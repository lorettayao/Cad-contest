module top(n0, n1, n6, n7, n2, n3, n8, n4, n5, n9, n10, n12, n13, n11, n14, n15, n16, n17, n18, n20, n19);
    input n0, n1, n2, n3, n4, n5;
    input [31:0] n6, n7, n8;
    output [31:0] n9, n10, n11;
    output n12, n13, n14, n15, n16, n17;
    output [7:0] n18, n19;
    output [15:0] n20;
    wire n0, n1, n2, n3, n4, n5;
    wire [31:0] n6, n7, n8;
    wire [31:0] n9, n10, n11;
    wire n12, n13, n14, n15, n16, n17;
    wire [7:0] n18, n19;
    wire [15:0] n20;
    wire [31:0] n21;
    wire [31:0] n22;
    wire [31:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [31:0] n26;
    wire [31:0] n27;
    wire [31:0] n28;
    wire [25:0] n29;
    wire [25:0] n30;
    wire [25:0] n31;
    wire [25:0] n32;
    wire [2:0] n33;
    wire [15:0] n34;
    wire [15:0] n35;
    wire [2:0] n36;
    wire [1:0] n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133;
    wire n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
    wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
    wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157;
    wire n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165;
    wire n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
    wire n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
    wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
    wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
    wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
    wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
    wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
    wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
    wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
    wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
    wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
    wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
    wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
    wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277;
    wire n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285;
    wire n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293;
    wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
    wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
    wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
    wire n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325;
    wire n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333;
    wire n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
    wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
    wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357;
    wire n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365;
    wire n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373;
    wire n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
    wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
    wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397;
    wire n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405;
    wire n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413;
    wire n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
    wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
    wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437;
    wire n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
    wire n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453;
    wire n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
    wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
    wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477;
    wire n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485;
    wire n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493;
    wire n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
    wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
    wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
    wire n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;
    wire n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533;
    wire n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541;
    wire n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549;
    wire n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557;
    wire n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565;
    wire n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573;
    wire n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581;
    wire n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589;
    wire n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597;
    wire n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605;
    wire n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613;
    wire n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
    wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629;
    wire n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637;
    wire n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645;
    wire n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653;
    wire n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661;
    wire n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669;
    wire n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677;
    wire n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685;
    wire n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693;
    wire n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701;
    wire n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709;
    wire n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717;
    wire n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725;
    wire n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733;
    wire n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741;
    wire n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749;
    wire n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757;
    wire n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765;
    wire n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773;
    wire n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781;
    wire n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789;
    wire n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797;
    wire n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805;
    wire n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813;
    wire n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821;
    wire n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829;
    wire n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837;
    wire n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845;
    wire n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853;
    wire n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861;
    wire n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869;
    wire n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877;
    wire n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885;
    wire n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893;
    wire n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
    wire n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909;
    wire n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917;
    wire n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925;
    wire n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;
    wire n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941;
    wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
    wire n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957;
    wire n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965;
    wire n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973;
    wire n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981;
    wire n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989;
    wire n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997;
    wire n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005;
    wire n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013;
    wire n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021;
    wire n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029;
    wire n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037;
    wire n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045;
    wire n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053;
    wire n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061;
    wire n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069;
    wire n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077;
    wire n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085;
    wire n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093;
    wire n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101;
    wire n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109;
    wire n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117;
    wire n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125;
    wire n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133;
    wire n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141;
    wire n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149;
    wire n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157;
    wire n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165;
    wire n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173;
    wire n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181;
    wire n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189;
    wire n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197;
    wire n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205;
    wire n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213;
    wire n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221;
    wire n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229;
    wire n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237;
    wire n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245;
    wire n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253;
    wire n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261;
    wire n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269;
    wire n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277;
    wire n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285;
    wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
    wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
    wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
    wire n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317;
    wire n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325;
    wire n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333;
    wire n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341;
    wire n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349;
    wire n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357;
    wire n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365;
    wire n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373;
    wire n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381;
    wire n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389;
    wire n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397;
    wire n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405;
    wire n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413;
    wire n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421;
    wire n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429;
    wire n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437;
    wire n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445;
    wire n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453;
    wire n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461;
    wire n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469;
    wire n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477;
    wire n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485;
    wire n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493;
    wire n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501;
    wire n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509;
    wire n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517;
    wire n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525;
    wire n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533;
    wire n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541;
    wire n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549;
    wire n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557;
    wire n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565;
    wire n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573;
    wire n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581;
    wire n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589;
    wire n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597;
    wire n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605;
    wire n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613;
    wire n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621;
    wire n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629;
    wire n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637;
    wire n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645;
    wire n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653;
    wire n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661;
    wire n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669;
    wire n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677;
    wire n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685;
    wire n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693;
    wire n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701;
    wire n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709;
    wire n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717;
    wire n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725;
    wire n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733;
    wire n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741;
    wire n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749;
    wire n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757;
    wire n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765;
    wire n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773;
    wire n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781;
    wire n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789;
    wire n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797;
    wire n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805;
    wire n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813;
    wire n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821;
    wire n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829;
    wire n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837;
    wire n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845;
    wire n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853;
    wire n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861;
    wire n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869;
    wire n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877;
    wire n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885;
    wire n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893;
    wire n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901;
    wire n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909;
    wire n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917;
    wire n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925;
    wire n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933;
    wire n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941;
    wire n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949;
    wire n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957;
    wire n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965;
    wire n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973;
    wire n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981;
    wire n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989;
    wire n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997;
    wire n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005;
    wire n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013;
    wire n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021;
    wire n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029;
    wire n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037;
    wire n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045;
    wire n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053;
    wire n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061;
    wire n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069;
    wire n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077;
    wire n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085;
    wire n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093;
    wire n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101;
    wire n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109;
    wire n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117;
    wire n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125;
    wire n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133;
    wire n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141;
    wire n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149;
    wire n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157;
    wire n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165;
    wire n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173;
    wire n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181;
    wire n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189;
    wire n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197;
    wire n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205;
    wire n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213;
    wire n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221;
    wire n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229;
    wire n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237;
    wire n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245;
    wire n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253;
    wire n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261;
    wire n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269;
    wire n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277;
    wire n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285;
    wire n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293;
    wire n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301;
    wire n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309;
    wire n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317;
    wire n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325;
    wire n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333;
    wire n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341;
    wire n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349;
    wire n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357;
    wire n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365;
    wire n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373;
    wire n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381;
    wire n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389;
    wire n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397;
    wire n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405;
    wire n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413;
    wire n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421;
    wire n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429;
    wire n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437;
    wire n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445;
    wire n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453;
    wire n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461;
    wire n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469;
    wire n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477;
    wire n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485;
    wire n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493;
    wire n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501;
    wire n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509;
    wire n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517;
    wire n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525;
    wire n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533;
    wire n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541;
    wire n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549;
    wire n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557;
    wire n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565;
    wire n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573;
    wire n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581;
    wire n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589;
    wire n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597;
    wire n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605;
    wire n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613;
    wire n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621;
    wire n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629;
    wire n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637;
    wire n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645;
    wire n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653;
    wire n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661;
    wire n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669;
    wire n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677;
    wire n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685;
    wire n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693;
    buf g0(n19[0], 1'b0);
    buf g1(n19[1], 1'b0);
    buf g2(n19[2], 1'b0);
    buf g3(n19[3], 1'b0);
    buf g4(n18[0], 1'b0);
    buf g5(n18[1], 1'b0);
    buf g6(n18[2], 1'b0);
    buf g7(n18[3], 1'b0);
    buf g8(n18[4], 1'b0);
    buf g9(n18[5], 1'b0);
    buf g10(n18[6], 1'b0);
    buf g11(n18[7], 1'b0);
    not g12(n4465 ,n1);
    not g13(n4464 ,n5);
    or g14(n4526 ,n4443 ,n4381);
    or g15(n4552 ,n4446 ,n4371);
    or g16(n4549 ,n4457 ,n4391);
    or g17(n4542 ,n4454 ,n4386);
    or g18(n4529 ,n4458 ,n4392);
    or g19(n4504 ,n4462 ,n4397);
    or g20(n4503 ,n4461 ,n4395);
    or g21(n4502 ,n4456 ,n4343);
    or g22(n4528 ,n4452 ,n4388);
    or g23(n4501 ,n4453 ,n4390);
    or g24(n4500 ,n4451 ,n4389);
    or g25(n4527 ,n4449 ,n4385);
    or g26(n4499 ,n4450 ,n4387);
    or g27(n4498 ,n4447 ,n4384);
    or g28(n4548 ,n4440 ,n4373);
    or g29(n4541 ,n4444 ,n4383);
    or g30(n4555 ,n4460 ,n4362);
    or g31(n4497 ,n4445 ,n4368);
    or g32(n4496 ,n4442 ,n4382);
    or g33(n4495 ,n4441 ,n4380);
    or g34(n4540 ,n4438 ,n4375);
    or g35(n4525 ,n4448 ,n4378);
    or g36(n4494 ,n4439 ,n4377);
    or g37(n4524 ,n4437 ,n4374);
    or g38(n4493 ,n4455 ,n4376);
    or g39(n4492 ,n4436 ,n4393);
    or g40(n4551 ,n4427 ,n4359);
    or g41(n4547 ,n4432 ,n4366);
    or g42(n4539 ,n4434 ,n4370);
    or g43(n4523 ,n4435 ,n4372);
    or g44(n4522 ,n4433 ,n4369);
    or g45(n4538 ,n4430 ,n4364);
    or g46(n4534 ,n4414 ,n4350);
    or g47(n4546 ,n4424 ,n4354);
    or g48(n4520 ,n4429 ,n4365);
    or g49(n4519 ,n4428 ,n4363);
    or g50(n4537 ,n4426 ,n4361);
    or g51(n4518 ,n4425 ,n4394);
    or g52(n4554 ,n4459 ,n4399);
    or g53(n4553 ,n4415 ,n4347);
    or g54(n4536 ,n4422 ,n4356);
    or g55(n4517 ,n4423 ,n4358);
    or g56(n4516 ,n4421 ,n4357);
    or g57(n4535 ,n4419 ,n4353);
    or g58(n4515 ,n4420 ,n4355);
    or g59(n4514 ,n4418 ,n4352);
    or g60(n4550 ,n4411 ,n4336);
    or g61(n4545 ,n4416 ,n4349);
    or g62(n4521 ,n4463 ,n4379);
    or g63(n4513 ,n4417 ,n4351);
    or g64(n4512 ,n4413 ,n4360);
    or g65(n4511 ,n4412 ,n4348);
    or g66(n4544 ,n4408 ,n4339);
    or g67(n4533 ,n4410 ,n4346);
    or g68(n4510 ,n4409 ,n4345);
    or g69(n4532 ,n4406 ,n4341);
    or g70(n4509 ,n4407 ,n4344);
    or g71(n4508 ,n4405 ,n4342);
    or g72(n4543 ,n4401 ,n4398);
    or g73(n4531 ,n4403 ,n4338);
    or g74(n4507 ,n4404 ,n4340);
    or g75(n4506 ,n4402 ,n4337);
    or g76(n4530 ,n4431 ,n4396);
    or g77(n4505 ,n4400 ,n4367);
    nor g78(n4463 ,n4206 ,n4215);
    nor g79(n4462 ,n4206 ,n4209);
    nor g80(n4461 ,n4206 ,n4267);
    nor g81(n4460 ,n4206 ,n4301);
    nor g82(n4459 ,n4206 ,n4212);
    nor g83(n4458 ,n4207 ,n4317);
    nor g84(n4457 ,n4206 ,n4313);
    nor g85(n4456 ,n4206 ,n4321);
    nor g86(n4455 ,n4206 ,n4328);
    nor g87(n4454 ,n4207 ,n4309);
    nor g88(n4453 ,n4207 ,n4310);
    nor g89(n4452 ,n4207 ,n4311);
    nor g90(n4451 ,n4207 ,n4260);
    nor g91(n4450 ,n4207 ,n4239);
    nor g92(n4449 ,n4207 ,n4293);
    nor g93(n4448 ,n4207 ,n4261);
    nor g94(n4447 ,n4206 ,n4298);
    nor g95(n4446 ,n4207 ,n4234);
    nor g96(n4445 ,n4206 ,n4289);
    nor g97(n4444 ,n4206 ,n4249);
    nor g98(n4443 ,n4207 ,n4228);
    nor g99(n4442 ,n4207 ,n4270);
    nor g100(n4441 ,n4207 ,n4256);
    nor g101(n4440 ,n4207 ,n4285);
    nor g102(n4439 ,n4206 ,n4211);
    nor g103(n4438 ,n4206 ,n4304);
    nor g104(n4437 ,n4207 ,n4236);
    nor g105(n4436 ,n4207 ,n4332);
    nor g106(n4435 ,n4206 ,n4251);
    nor g107(n4434 ,n4206 ,n4292);
    nor g108(n4433 ,n4207 ,n4248);
    nor g109(n4432 ,n4207 ,n4245);
    nor g110(n4431 ,n4207 ,n4221);
    nor g111(n4430 ,n4206 ,n4244);
    nor g112(n4429 ,n4206 ,n4282);
    nor g113(n4428 ,n4207 ,n4214);
    nor g114(n4427 ,n4206 ,n4208);
    nor g115(n4426 ,n4207 ,n4265);
    nor g116(n4425 ,n4206 ,n4275);
    nor g117(n4424 ,n4206 ,n4320);
    nor g118(n4423 ,n4206 ,n4277);
    nor g119(n4422 ,n4206 ,n4266);
    nor g120(n4421 ,n4207 ,n4329);
    nor g121(n4420 ,n4207 ,n4264);
    nor g122(n4419 ,n4206 ,n4318);
    nor g123(n4418 ,n4207 ,n4254);
    nor g124(n4417 ,n4207 ,n4314);
    nor g125(n4416 ,n4207 ,n4302);
    nor g126(n4415 ,n4207 ,n4290);
    nor g127(n4414 ,n4207 ,n4306);
    nor g128(n4413 ,n4207 ,n4307);
    nor g129(n4412 ,n4206 ,n4252);
    nor g130(n4411 ,n4206 ,n4308);
    nor g131(n4410 ,n4207 ,n4295);
    nor g132(n4409 ,n4206 ,n4286);
    nor g133(n4408 ,n4206 ,n4284);
    nor g134(n4407 ,n4206 ,n4242);
    nor g135(n4406 ,n4206 ,n4217);
    nor g136(n4405 ,n4206 ,n4281);
    nor g137(n4404 ,n4206 ,n4263);
    nor g138(n4403 ,n4206 ,n4273);
    nor g139(n4402 ,n4207 ,n4220);
    nor g140(n4401 ,n4207 ,n4237);
    nor g141(n4400 ,n4207 ,n4269);
    nor g142(n4399 ,n4224 ,n4204);
    nor g143(n4398 ,n4325 ,n4204);
    nor g144(n4397 ,n4319 ,n4204);
    nor g145(n4396 ,n4327 ,n4204);
    nor g146(n4395 ,n4303 ,n4205);
    nor g147(n4394 ,n4240 ,n4205);
    nor g148(n4393 ,n4333 ,n4204);
    nor g149(n4392 ,n4250 ,n4205);
    nor g150(n4391 ,n4276 ,n4205);
    nor g151(n4390 ,n4296 ,n4205);
    nor g152(n4389 ,n4305 ,n4205);
    nor g153(n4388 ,n4322 ,n4204);
    nor g154(n4387 ,n4233 ,n4204);
    nor g155(n4386 ,n4335 ,n4204);
    nor g156(n4385 ,n4259 ,n4204);
    nor g157(n4384 ,n4294 ,n4204);
    nor g158(n4383 ,n4218 ,n4204);
    nor g159(n4382 ,n4257 ,n4205);
    nor g160(n4381 ,n4272 ,n4204);
    nor g161(n4380 ,n4231 ,n4204);
    nor g162(n4379 ,n4225 ,n4204);
    nor g163(n4378 ,n4334 ,n4204);
    nor g164(n4377 ,n4287 ,n4204);
    nor g165(n4376 ,n4262 ,n4204);
    nor g166(n4375 ,n4300 ,n4204);
    nor g167(n4374 ,n4253 ,n4204);
    nor g168(n4373 ,n4216 ,n4204);
    nor g169(n4372 ,n4227 ,n4204);
    nor g170(n4371 ,n4226 ,n4205);
    nor g171(n4370 ,n4288 ,n4204);
    nor g172(n4369 ,n4247 ,n4204);
    nor g173(n4368 ,n4229 ,n4204);
    nor g174(n4367 ,n4213 ,n4204);
    nor g175(n4366 ,n4223 ,n4204);
    nor g176(n4365 ,n4243 ,n4205);
    nor g177(n4364 ,n4280 ,n4204);
    nor g178(n4363 ,n4241 ,n4204);
    nor g179(n4362 ,n4331 ,n4205);
    nor g180(n4361 ,n4222 ,n4205);
    nor g181(n4360 ,n4238 ,n4204);
    nor g182(n4359 ,n4258 ,n4204);
    nor g183(n4358 ,n4230 ,n4204);
    nor g184(n4357 ,n4330 ,n4204);
    nor g185(n4356 ,n4326 ,n4204);
    nor g186(n4355 ,n4324 ,n4204);
    nor g187(n4354 ,n4323 ,n4204);
    nor g188(n4353 ,n4315 ,n4205);
    nor g189(n4352 ,n4316 ,n4204);
    nor g190(n4351 ,n4312 ,n4204);
    nor g191(n4350 ,n4246 ,n4205);
    nor g192(n4349 ,n4299 ,n4204);
    nor g193(n4348 ,n4297 ,n4205);
    nor g194(n4347 ,n4255 ,n4204);
    nor g195(n4346 ,n4210 ,n4204);
    nor g196(n4345 ,n4291 ,n4204);
    nor g197(n4344 ,n4283 ,n4204);
    nor g198(n4343 ,n4271 ,n4204);
    nor g199(n4342 ,n4279 ,n4205);
    nor g200(n4341 ,n4232 ,n4204);
    nor g201(n4340 ,n4219 ,n4204);
    nor g202(n4339 ,n4278 ,n4204);
    nor g203(n4338 ,n4274 ,n4205);
    nor g204(n4337 ,n4268 ,n4204);
    nor g205(n4336 ,n4235 ,n4204);
    not g206(n4335 ,n21[18]);
    not g207(n4334 ,n21[1]);
    not g208(n4333 ,n22[0]);
    not g209(n4332 ,n23[0]);
    not g210(n4331 ,n21[31]);
    not g211(n4330 ,n22[24]);
    not g212(n4329 ,n23[24]);
    not g213(n4328 ,n23[1]);
    not g214(n4327 ,n21[6]);
    not g215(n4326 ,n21[12]);
    not g216(n4325 ,n21[19]);
    not g217(n4324 ,n22[23]);
    not g218(n4323 ,n21[22]);
    not g219(n4322 ,n21[4]);
    not g220(n4321 ,n23[10]);
    not g221(n4320 ,n24[22]);
    not g222(n4319 ,n22[12]);
    not g223(n4318 ,n24[11]);
    not g224(n4317 ,n24[5]);
    not g225(n4316 ,n22[22]);
    not g226(n4315 ,n21[11]);
    not g227(n4314 ,n23[21]);
    not g228(n4313 ,n24[25]);
    not g229(n4312 ,n22[21]);
    not g230(n4311 ,n24[4]);
    not g231(n4310 ,n23[9]);
    not g232(n4309 ,n24[18]);
    not g233(n4308 ,n24[26]);
    not g234(n4307 ,n23[20]);
    not g235(n4306 ,n24[10]);
    not g236(n4305 ,n22[8]);
    not g237(n4304 ,n24[16]);
    not g238(n4303 ,n22[11]);
    not g239(n4302 ,n24[21]);
    not g240(n4301 ,n24[31]);
    not g241(n4300 ,n21[16]);
    not g242(n4299 ,n21[21]);
    not g243(n4298 ,n23[6]);
    not g244(n4297 ,n22[19]);
    not g245(n4296 ,n22[9]);
    not g246(n4295 ,n24[9]);
    not g247(n4294 ,n22[6]);
    not g248(n4293 ,n24[3]);
    not g249(n4292 ,n24[15]);
    not g250(n4291 ,n22[18]);
    not g251(n4290 ,n24[29]);
    not g252(n4289 ,n23[5]);
    not g253(n4288 ,n21[15]);
    not g254(n4287 ,n22[2]);
    not g255(n4286 ,n23[18]);
    not g256(n4285 ,n24[24]);
    not g257(n4284 ,n24[20]);
    not g258(n4283 ,n22[17]);
    not g259(n4282 ,n23[28]);
    not g260(n4281 ,n23[16]);
    not g261(n4280 ,n21[14]);
    not g262(n4279 ,n22[16]);
    not g263(n4278 ,n21[20]);
    not g264(n4277 ,n23[25]);
    not g265(n4276 ,n21[25]);
    not g266(n4275 ,n23[26]);
    not g267(n4274 ,n21[7]);
    not g268(n4273 ,n24[7]);
    not g269(n4206 ,n4205);
    not g270(n4205 ,n4207);
    not g271(n4204 ,n4207);
    not g272(n4207 ,n6[5]);
    not g273(n4272 ,n21[2]);
    not g274(n4271 ,n22[10]);
    not g275(n4270 ,n23[4]);
    not g276(n4269 ,n23[13]);
    not g277(n4268 ,n22[14]);
    not g278(n4267 ,n23[11]);
    not g279(n4266 ,n24[12]);
    not g280(n4265 ,n24[13]);
    not g281(n4264 ,n23[23]);
    not g282(n4263 ,n23[15]);
    not g283(n4262 ,n22[1]);
    not g284(n4261 ,n24[1]);
    not g285(n4260 ,n23[8]);
    not g286(n4259 ,n21[3]);
    not g287(n4258 ,n21[27]);
    not g288(n4257 ,n22[4]);
    not g289(n4256 ,n23[3]);
    not g290(n4255 ,n21[29]);
    not g291(n4254 ,n23[22]);
    not g292(n4253 ,n21[0]);
    not g293(n4252 ,n23[19]);
    not g294(n4251 ,n23[31]);
    not g295(n4250 ,n21[5]);
    not g296(n4249 ,n24[17]);
    not g297(n4248 ,n23[30]);
    not g298(n4247 ,n22[30]);
    not g299(n4246 ,n21[10]);
    not g300(n4245 ,n24[23]);
    not g301(n4244 ,n24[14]);
    not g302(n4243 ,n22[28]);
    not g303(n4242 ,n23[17]);
    not g304(n4241 ,n22[27]);
    not g305(n4240 ,n22[26]);
    not g306(n4239 ,n23[7]);
    not g307(n4238 ,n22[20]);
    not g308(n4237 ,n24[19]);
    not g309(n4236 ,n24[0]);
    not g310(n4235 ,n21[26]);
    not g311(n4234 ,n24[28]);
    not g312(n4233 ,n22[7]);
    not g313(n4232 ,n21[8]);
    not g314(n4231 ,n22[3]);
    not g315(n4230 ,n22[25]);
    not g316(n4229 ,n22[5]);
    not g317(n4228 ,n24[2]);
    not g318(n4227 ,n22[31]);
    not g319(n4226 ,n21[28]);
    not g320(n4225 ,n22[29]);
    not g321(n4224 ,n21[30]);
    not g322(n4223 ,n21[23]);
    not g323(n4222 ,n21[13]);
    not g324(n4221 ,n24[6]);
    not g325(n4220 ,n23[14]);
    not g326(n4219 ,n22[15]);
    not g327(n4218 ,n21[17]);
    not g328(n4217 ,n24[8]);
    not g329(n4216 ,n21[24]);
    not g330(n4215 ,n23[29]);
    not g331(n4214 ,n23[27]);
    not g332(n4213 ,n22[13]);
    not g333(n4212 ,n24[30]);
    not g334(n4211 ,n23[2]);
    not g335(n4210 ,n21[9]);
    not g336(n4209 ,n23[12]);
    not g337(n4208 ,n24[27]);
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3266), .Q(n25[0]));
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3264), .Q(n25[1]));
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3280), .Q(n25[2]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3278), .Q(n25[3]));
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3273), .Q(n25[4]));
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3268), .Q(n25[5]));
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3263), .Q(n25[6]));
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3256), .Q(n25[7]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3253), .Q(n25[8]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3252), .Q(n25[9]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3247), .Q(n25[10]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3245), .Q(n25[11]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3242), .Q(n25[12]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3241), .Q(n25[13]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3240), .Q(n25[14]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3239), .Q(n25[15]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3238), .Q(n25[16]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3237), .Q(n25[17]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3236), .Q(n25[18]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3235), .Q(n25[19]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3234), .Q(n25[20]));
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3233), .Q(n25[21]));
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3232), .Q(n25[22]));
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3231), .Q(n25[23]));
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3229), .Q(n25[24]));
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3230), .Q(n25[25]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3228), .Q(n25[26]));
    dff g365(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3227), .Q(n25[27]));
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3226), .Q(n25[28]));
    dff g367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3225), .Q(n25[29]));
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3224), .Q(n25[30]));
    dff g369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3223), .Q(n25[31]));
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3222), .Q(n26[0]));
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3221), .Q(n26[1]));
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3220), .Q(n26[2]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3219), .Q(n26[3]));
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3218), .Q(n26[4]));
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3217), .Q(n26[5]));
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3216), .Q(n26[6]));
    dff g377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3215), .Q(n26[7]));
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3214), .Q(n26[8]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3213), .Q(n26[9]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3212), .Q(n26[10]));
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3211), .Q(n26[11]));
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3210), .Q(n26[12]));
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3207), .Q(n26[13]));
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3209), .Q(n26[14]));
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3208), .Q(n26[15]));
    dff g386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3206), .Q(n26[16]));
    dff g387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3204), .Q(n26[17]));
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3205), .Q(n26[18]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3203), .Q(n26[19]));
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3202), .Q(n26[20]));
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3200), .Q(n26[21]));
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3199), .Q(n26[22]));
    dff g393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3197), .Q(n26[23]));
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3195), .Q(n26[24]));
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3192), .Q(n26[25]));
    dff g396(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3190), .Q(n26[26]));
    dff g397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3191), .Q(n26[27]));
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3189), .Q(n26[28]));
    dff g399(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3188), .Q(n26[29]));
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3187), .Q(n26[30]));
    dff g401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3186), .Q(n26[31]));
    dff g402(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3178), .Q(n27[0]));
    dff g403(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3181), .Q(n27[1]));
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3174), .Q(n27[2]));
    dff g405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3172), .Q(n27[3]));
    dff g406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3169), .Q(n27[4]));
    dff g407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3165), .Q(n27[5]));
    dff g408(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3163), .Q(n27[6]));
    dff g409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3157), .Q(n27[7]));
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3155), .Q(n27[8]));
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3151), .Q(n27[9]));
    dff g412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3269), .Q(n27[10]));
    dff g413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3147), .Q(n27[11]));
    dff g414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3142), .Q(n27[12]));
    dff g415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3140), .Q(n27[13]));
    dff g416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3134), .Q(n27[14]));
    dff g417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3246), .Q(n27[15]));
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3128), .Q(n27[16]));
    dff g419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3126), .Q(n27[17]));
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3116), .Q(n27[18]));
    dff g421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3196), .Q(n27[19]));
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3118), .Q(n27[20]));
    dff g423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3113), .Q(n27[21]));
    dff g424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3110), .Q(n27[22]));
    dff g425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3243), .Q(n27[23]));
    dff g426(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3103), .Q(n27[24]));
    dff g427(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3100), .Q(n27[25]));
    dff g428(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3096), .Q(n27[26]));
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3272), .Q(n27[27]));
    dff g430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3094), .Q(n27[28]));
    dff g431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3154), .Q(n27[29]));
    dff g432(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3091), .Q(n27[30]));
    dff g433(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3309), .Q(n27[31]));
    dff g434(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3314), .Q(n28[0]));
    dff g435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3307), .Q(n28[1]));
    dff g436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3302), .Q(n28[2]));
    dff g437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3297), .Q(n28[3]));
    dff g438(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3296), .Q(n28[4]));
    dff g439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3292), .Q(n28[5]));
    dff g440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3290), .Q(n28[6]));
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3476), .Q(n28[7]));
    dff g442(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3089), .Q(n28[8]));
    dff g443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3285), .Q(n28[9]));
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3284), .Q(n28[10]));
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3283), .Q(n28[11]));
    dff g446(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3282), .Q(n28[12]));
    dff g447(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3281), .Q(n28[13]));
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3279), .Q(n28[14]));
    dff g449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3277), .Q(n28[15]));
    dff g450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3276), .Q(n28[16]));
    dff g451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3275), .Q(n28[17]));
    dff g452(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3274), .Q(n28[18]));
    dff g453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3271), .Q(n28[19]));
    dff g454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3270), .Q(n28[20]));
    dff g455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3267), .Q(n28[21]));
    dff g456(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3265), .Q(n28[22]));
    dff g457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3262), .Q(n28[23]));
    dff g458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3260), .Q(n28[24]));
    dff g459(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3258), .Q(n28[25]));
    dff g460(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3257), .Q(n28[26]));
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3255), .Q(n28[27]));
    dff g462(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3254), .Q(n28[28]));
    dff g463(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3251), .Q(n28[29]));
    dff g464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3250), .Q(n28[30]));
    dff g465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3248), .Q(n28[31]));
    dff g466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3559), .Q(n16));
    dff g467(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3558), .Q(n17));
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3185), .Q(n29[0]));
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3184), .Q(n29[1]));
    dff g470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3183), .Q(n29[2]));
    dff g471(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3180), .Q(n29[3]));
    dff g472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3179), .Q(n29[4]));
    dff g473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3177), .Q(n29[5]));
    dff g474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3176), .Q(n29[6]));
    dff g475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3175), .Q(n29[7]));
    dff g476(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3173), .Q(n29[8]));
    dff g477(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3171), .Q(n29[9]));
    dff g478(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3170), .Q(n29[10]));
    dff g479(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3168), .Q(n29[11]));
    dff g480(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3167), .Q(n29[12]));
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3166), .Q(n29[13]));
    dff g482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3164), .Q(n29[14]));
    dff g483(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3162), .Q(n29[15]));
    dff g484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3161), .Q(n29[16]));
    dff g485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3160), .Q(n29[17]));
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3159), .Q(n29[18]));
    dff g487(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3158), .Q(n29[19]));
    dff g488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3156), .Q(n29[20]));
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3244), .Q(n29[21]));
    dff g490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3153), .Q(n29[22]));
    dff g491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3249), .Q(n29[23]));
    dff g492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3152), .Q(n29[24]));
    dff g493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3150), .Q(n29[25]));
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3259), .Q(n30[0]));
    dff g495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3149), .Q(n30[1]));
    dff g496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3148), .Q(n30[2]));
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3145), .Q(n30[3]));
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3144), .Q(n30[4]));
    dff g499(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3143), .Q(n30[5]));
    dff g500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3141), .Q(n30[6]));
    dff g501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3139), .Q(n30[7]));
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3136), .Q(n30[8]));
    dff g503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3182), .Q(n30[9]));
    dff g504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3135), .Q(n30[10]));
    dff g505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3133), .Q(n30[11]));
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3132), .Q(n30[12]));
    dff g507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3131), .Q(n30[13]));
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3130), .Q(n30[14]));
    dff g509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3129), .Q(n30[15]));
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3127), .Q(n30[16]));
    dff g511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3125), .Q(n30[17]));
    dff g512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3124), .Q(n30[18]));
    dff g513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3123), .Q(n30[19]));
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3122), .Q(n30[20]));
    dff g515(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3121), .Q(n30[21]));
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3120), .Q(n30[22]));
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3119), .Q(n30[23]));
    dff g518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3201), .Q(n30[24]));
    dff g519(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3117), .Q(n30[25]));
    dff g520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3115), .Q(n31[0]));
    dff g521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3114), .Q(n31[1]));
    dff g522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3112), .Q(n31[2]));
    dff g523(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3111), .Q(n31[3]));
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3108), .Q(n31[4]));
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3107), .Q(n31[5]));
    dff g526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3106), .Q(n31[6]));
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3138), .Q(n31[7]));
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3105), .Q(n31[8]));
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3104), .Q(n31[9]));
    dff g530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3102), .Q(n31[10]));
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3101), .Q(n31[11]));
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3099), .Q(n31[12]));
    dff g533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3198), .Q(n31[13]));
    dff g534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3098), .Q(n31[14]));
    dff g535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3097), .Q(n31[15]));
    dff g536(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3261), .Q(n31[16]));
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3193), .Q(n31[17]));
    dff g538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3109), .Q(n31[18]));
    dff g539(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3095), .Q(n31[19]));
    dff g540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3137), .Q(n31[20]));
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3146), .Q(n31[21]));
    dff g542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3093), .Q(n31[22]));
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3092), .Q(n31[23]));
    dff g544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3194), .Q(n31[24]));
    dff g545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3090), .Q(n31[25]));
    dff g546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3286), .Q(n32[0]));
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3315), .Q(n32[1]));
    dff g548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3313), .Q(n32[2]));
    dff g549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3312), .Q(n32[3]));
    dff g550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3311), .Q(n32[4]));
    dff g551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3310), .Q(n32[5]));
    dff g552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3308), .Q(n32[6]));
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3306), .Q(n32[7]));
    dff g554(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3305), .Q(n32[8]));
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3304), .Q(n32[9]));
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3303), .Q(n32[10]));
    dff g557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3301), .Q(n32[11]));
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3300), .Q(n32[12]));
    dff g559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3299), .Q(n32[13]));
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3298), .Q(n32[14]));
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3295), .Q(n32[15]));
    dff g562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3294), .Q(n32[16]));
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3293), .Q(n32[17]));
    dff g564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3291), .Q(n32[18]));
    dff g565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3289), .Q(n32[19]));
    dff g566(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3288), .Q(n32[20]));
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3287), .Q(n32[21]));
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3316), .Q(n32[22]));
    dff g569(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3477), .Q(n32[23]));
    dff g570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3478), .Q(n32[24]));
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3479), .Q(n32[25]));
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2618), .Q(n128));
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2617), .Q(n129));
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2616), .Q(n130));
    dff g575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2615), .Q(n131));
    dff g576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4202), .Q(n11[0]));
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4198), .Q(n11[1]));
    dff g578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4201), .Q(n11[2]));
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4197), .Q(n11[3]));
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4200), .Q(n11[4]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4199), .Q(n11[5]));
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4203), .Q(n11[6]));
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4196), .Q(n11[7]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4195), .Q(n11[8]));
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4194), .Q(n11[9]));
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4193), .Q(n11[10]));
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4192), .Q(n11[11]));
    dff g588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4168), .Q(n11[12]));
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4190), .Q(n11[13]));
    dff g590(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4189), .Q(n11[14]));
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4188), .Q(n11[15]));
    dff g592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4187), .Q(n11[16]));
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4186), .Q(n11[17]));
    dff g594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4185), .Q(n11[18]));
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4184), .Q(n11[19]));
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4183), .Q(n11[20]));
    dff g597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4182), .Q(n11[21]));
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4181), .Q(n11[22]));
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4180), .Q(n11[23]));
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4179), .Q(n11[24]));
    dff g601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4178), .Q(n11[25]));
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4177), .Q(n11[26]));
    dff g603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4175), .Q(n11[27]));
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4176), .Q(n11[28]));
    dff g605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4174), .Q(n11[29]));
    dff g606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4173), .Q(n11[30]));
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4172), .Q(n11[31]));
    dff g608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3958), .Q(n14));
    dff g609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3957), .Q(n15));
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n33[0]));
    dff g611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1610), .Q(n33[1]));
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n33[2]));
    dff g613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1609), .Q(n19[4]));
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1608), .Q(n19[5]));
    dff g615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n19[6]));
    dff g616(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n19[7]));
    dff g617(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3581), .Q(n34[0]));
    dff g618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3580), .Q(n34[1]));
    dff g619(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3579), .Q(n34[2]));
    dff g620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3578), .Q(n34[3]));
    dff g621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3577), .Q(n34[4]));
    dff g622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3576), .Q(n34[5]));
    dff g623(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3575), .Q(n34[6]));
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3574), .Q(n34[7]));
    dff g625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3444), .Q(n21[0]));
    dff g626(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3443), .Q(n21[1]));
    dff g627(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3442), .Q(n21[2]));
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3441), .Q(n21[3]));
    dff g629(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3440), .Q(n21[4]));
    dff g630(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3439), .Q(n21[5]));
    dff g631(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3437), .Q(n21[6]));
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3438), .Q(n21[7]));
    dff g633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3436), .Q(n21[8]));
    dff g634(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3435), .Q(n21[9]));
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3434), .Q(n21[10]));
    dff g636(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3433), .Q(n21[11]));
    dff g637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3432), .Q(n21[12]));
    dff g638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3431), .Q(n21[13]));
    dff g639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3430), .Q(n21[14]));
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3429), .Q(n21[15]));
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3428), .Q(n21[16]));
    dff g642(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3427), .Q(n21[17]));
    dff g643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3426), .Q(n21[18]));
    dff g644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3425), .Q(n21[19]));
    dff g645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3424), .Q(n21[20]));
    dff g646(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3423), .Q(n21[21]));
    dff g647(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3422), .Q(n21[22]));
    dff g648(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3421), .Q(n21[23]));
    dff g649(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3420), .Q(n21[24]));
    dff g650(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3419), .Q(n21[25]));
    dff g651(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3418), .Q(n21[26]));
    dff g652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3417), .Q(n21[27]));
    dff g653(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3416), .Q(n21[28]));
    dff g654(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3415), .Q(n21[29]));
    dff g655(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3414), .Q(n21[30]));
    dff g656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3413), .Q(n21[31]));
    dff g657(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3412), .Q(n22[0]));
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3411), .Q(n22[1]));
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3410), .Q(n22[2]));
    dff g660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3409), .Q(n22[3]));
    dff g661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3408), .Q(n22[4]));
    dff g662(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3407), .Q(n22[5]));
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3406), .Q(n22[6]));
    dff g664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3405), .Q(n22[7]));
    dff g665(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3404), .Q(n22[8]));
    dff g666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3403), .Q(n22[9]));
    dff g667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3402), .Q(n22[10]));
    dff g668(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3401), .Q(n22[11]));
    dff g669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3400), .Q(n22[12]));
    dff g670(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3399), .Q(n22[13]));
    dff g671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3398), .Q(n22[14]));
    dff g672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3397), .Q(n22[15]));
    dff g673(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3396), .Q(n22[16]));
    dff g674(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3395), .Q(n22[17]));
    dff g675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3394), .Q(n22[18]));
    dff g676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3392), .Q(n22[19]));
    dff g677(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3393), .Q(n22[20]));
    dff g678(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3391), .Q(n22[21]));
    dff g679(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3390), .Q(n22[22]));
    dff g680(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3389), .Q(n22[23]));
    dff g681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3388), .Q(n22[24]));
    dff g682(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3387), .Q(n22[25]));
    dff g683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3386), .Q(n22[26]));
    dff g684(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3385), .Q(n22[27]));
    dff g685(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3384), .Q(n22[28]));
    dff g686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3383), .Q(n22[29]));
    dff g687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3382), .Q(n22[30]));
    dff g688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3381), .Q(n22[31]));
    dff g689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3380), .Q(n24[0]));
    dff g690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3379), .Q(n24[1]));
    dff g691(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3378), .Q(n24[2]));
    dff g692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3377), .Q(n24[3]));
    dff g693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3376), .Q(n24[4]));
    dff g694(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3375), .Q(n24[5]));
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3374), .Q(n24[6]));
    dff g696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3373), .Q(n24[7]));
    dff g697(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3372), .Q(n24[8]));
    dff g698(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3371), .Q(n24[9]));
    dff g699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3370), .Q(n24[10]));
    dff g700(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3369), .Q(n24[11]));
    dff g701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3368), .Q(n24[12]));
    dff g702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3367), .Q(n24[13]));
    dff g703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3366), .Q(n24[14]));
    dff g704(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3365), .Q(n24[15]));
    dff g705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3364), .Q(n24[16]));
    dff g706(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3363), .Q(n24[17]));
    dff g707(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3362), .Q(n24[18]));
    dff g708(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3361), .Q(n24[19]));
    dff g709(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3360), .Q(n24[20]));
    dff g710(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3359), .Q(n24[21]));
    dff g711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3358), .Q(n24[22]));
    dff g712(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3357), .Q(n24[23]));
    dff g713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3356), .Q(n24[24]));
    dff g714(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3355), .Q(n24[25]));
    dff g715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3354), .Q(n24[26]));
    dff g716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3353), .Q(n24[27]));
    dff g717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3352), .Q(n24[28]));
    dff g718(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3351), .Q(n24[29]));
    dff g719(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3350), .Q(n24[30]));
    dff g720(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3349), .Q(n24[31]));
    dff g721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3348), .Q(n23[0]));
    dff g722(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3347), .Q(n23[1]));
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3346), .Q(n23[2]));
    dff g724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3345), .Q(n23[3]));
    dff g725(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3344), .Q(n23[4]));
    dff g726(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3343), .Q(n23[5]));
    dff g727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3342), .Q(n23[6]));
    dff g728(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3341), .Q(n23[7]));
    dff g729(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3340), .Q(n23[8]));
    dff g730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3339), .Q(n23[9]));
    dff g731(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3338), .Q(n23[10]));
    dff g732(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3337), .Q(n23[11]));
    dff g733(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3336), .Q(n23[12]));
    dff g734(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3335), .Q(n23[13]));
    dff g735(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3334), .Q(n23[14]));
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3333), .Q(n23[15]));
    dff g737(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3332), .Q(n23[16]));
    dff g738(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3331), .Q(n23[17]));
    dff g739(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3328), .Q(n23[18]));
    dff g740(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3330), .Q(n23[19]));
    dff g741(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3329), .Q(n23[20]));
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3327), .Q(n23[21]));
    dff g743(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3326), .Q(n23[22]));
    dff g744(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3325), .Q(n23[23]));
    dff g745(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3324), .Q(n23[24]));
    dff g746(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3323), .Q(n23[25]));
    dff g747(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3322), .Q(n23[26]));
    dff g748(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3321), .Q(n23[27]));
    dff g749(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3320), .Q(n23[28]));
    dff g750(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3319), .Q(n23[29]));
    dff g751(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3318), .Q(n23[30]));
    dff g752(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3317), .Q(n23[31]));
    dff g753(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3951), .Q(n9[0]));
    dff g754(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3956), .Q(n9[1]));
    dff g755(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3955), .Q(n9[2]));
    dff g756(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3954), .Q(n9[3]));
    dff g757(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3953), .Q(n9[4]));
    dff g758(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4081), .Q(n9[5]));
    dff g759(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4169), .Q(n9[6]));
    dff g760(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4167), .Q(n9[7]));
    dff g761(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4171), .Q(n9[8]));
    dff g762(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4170), .Q(n9[9]));
    dff g763(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4191), .Q(n9[10]));
    dff g764(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4166), .Q(n9[11]));
    dff g765(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4163), .Q(n9[12]));
    dff g766(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4165), .Q(n9[13]));
    dff g767(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4164), .Q(n9[14]));
    dff g768(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4162), .Q(n9[15]));
    dff g769(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4161), .Q(n9[16]));
    dff g770(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4160), .Q(n9[17]));
    dff g771(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4159), .Q(n9[18]));
    dff g772(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4158), .Q(n9[19]));
    dff g773(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4157), .Q(n9[20]));
    dff g774(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4156), .Q(n9[21]));
    dff g775(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4155), .Q(n9[22]));
    dff g776(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4154), .Q(n9[23]));
    dff g777(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4153), .Q(n9[24]));
    dff g778(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4151), .Q(n9[25]));
    dff g779(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4152), .Q(n9[26]));
    dff g780(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4150), .Q(n9[27]));
    dff g781(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4149), .Q(n9[28]));
    dff g782(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4148), .Q(n9[29]));
    dff g783(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4147), .Q(n9[30]));
    dff g784(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4146), .Q(n9[31]));
    dff g785(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n12));
    dff g786(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4138), .Q(n10[0]));
    dff g787(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4137), .Q(n10[1]));
    dff g788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4135), .Q(n10[2]));
    dff g789(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4136), .Q(n10[3]));
    dff g790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4134), .Q(n10[4]));
    dff g791(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4133), .Q(n10[5]));
    dff g792(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4132), .Q(n10[6]));
    dff g793(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4130), .Q(n10[7]));
    dff g794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4131), .Q(n10[8]));
    dff g795(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4129), .Q(n10[9]));
    dff g796(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4128), .Q(n10[10]));
    dff g797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4127), .Q(n10[11]));
    dff g798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4126), .Q(n10[12]));
    dff g799(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4125), .Q(n10[13]));
    dff g800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4124), .Q(n10[14]));
    dff g801(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4123), .Q(n10[15]));
    dff g802(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4122), .Q(n10[16]));
    dff g803(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4121), .Q(n10[17]));
    dff g804(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4120), .Q(n10[18]));
    dff g805(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4119), .Q(n10[19]));
    dff g806(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4118), .Q(n10[20]));
    dff g807(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4117), .Q(n10[21]));
    dff g808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4116), .Q(n10[22]));
    dff g809(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4115), .Q(n10[23]));
    dff g810(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4114), .Q(n10[24]));
    dff g811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4113), .Q(n10[25]));
    dff g812(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4112), .Q(n10[26]));
    dff g813(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4111), .Q(n10[27]));
    dff g814(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4110), .Q(n10[28]));
    dff g815(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4109), .Q(n10[29]));
    dff g816(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4108), .Q(n10[30]));
    dff g817(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n4107), .Q(n10[31]));
    dff g818(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3657), .Q(n13));
    dff g819(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3571), .Q(n35[0]));
    dff g820(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3570), .Q(n35[1]));
    dff g821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3569), .Q(n35[2]));
    dff g822(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3568), .Q(n35[3]));
    dff g823(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3567), .Q(n35[4]));
    dff g824(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3566), .Q(n35[5]));
    dff g825(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3572), .Q(n35[6]));
    dff g826(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3573), .Q(n35[7]));
    dff g827(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3492), .Q(n36[0]));
    dff g828(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3583), .Q(n36[1]));
    dff g829(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3491), .Q(n36[2]));
    dff g830(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n20[0]));
    dff g831(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n20[1]));
    dff g832(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n20[2]));
    dff g833(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1612), .Q(n20[3]));
    dff g834(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1614), .Q(n20[4]));
    dff g835(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1613), .Q(n20[5]));
    dff g836(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n20[6]));
    dff g837(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n20[7]));
    dff g838(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1611), .Q(n20[8]));
    dff g839(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n20[9]));
    dff g840(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n20[10]));
    dff g841(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n20[11]));
    dff g842(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1591), .Q(n20[12]));
    dff g843(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n20[13]));
    dff g844(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1616), .Q(n20[14]));
    dff g845(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1615), .Q(n20[15]));
    or g846(n4203 ,n4010 ,n4142);
    or g847(n4202 ,n4019 ,n4106);
    or g848(n4201 ,n4018 ,n4104);
    or g849(n4200 ,n4014 ,n4140);
    or g850(n4199 ,n4012 ,n4141);
    or g851(n4198 ,n4021 ,n4105);
    or g852(n4197 ,n4016 ,n4139);
    or g853(n4196 ,n4008 ,n4143);
    or g854(n4195 ,n4006 ,n4144);
    or g855(n4194 ,n4004 ,n4145);
    or g856(n4193 ,n4002 ,n4055);
    or g857(n4192 ,n4000 ,n4102);
    or g858(n4191 ,n3467 ,n4076);
    or g859(n4190 ,n3996 ,n4098);
    or g860(n4189 ,n3994 ,n4100);
    or g861(n4188 ,n3992 ,n4099);
    or g862(n4187 ,n4054 ,n4097);
    or g863(n4186 ,n3988 ,n4096);
    or g864(n4185 ,n3986 ,n4095);
    or g865(n4184 ,n3984 ,n4094);
    or g866(n4183 ,n3983 ,n4093);
    or g867(n4182 ,n3980 ,n4092);
    or g868(n4181 ,n3978 ,n4091);
    or g869(n4180 ,n3976 ,n4090);
    or g870(n4179 ,n3974 ,n4089);
    or g871(n4178 ,n3972 ,n4088);
    or g872(n4177 ,n3968 ,n4087);
    or g873(n4176 ,n3966 ,n4085);
    or g874(n4175 ,n3969 ,n4086);
    or g875(n4174 ,n3964 ,n4084);
    or g876(n4173 ,n3962 ,n4083);
    or g877(n4172 ,n3960 ,n4082);
    or g878(n4171 ,n3469 ,n4078);
    or g879(n4170 ,n3468 ,n4077);
    or g880(n4169 ,n3471 ,n4080);
    or g881(n4168 ,n3998 ,n4101);
    or g882(n4167 ,n3470 ,n4079);
    or g883(n4166 ,n3466 ,n4075);
    or g884(n4165 ,n3464 ,n4073);
    or g885(n4164 ,n3463 ,n4072);
    or g886(n4163 ,n3465 ,n4074);
    or g887(n4162 ,n3462 ,n4071);
    or g888(n4161 ,n3461 ,n4070);
    or g889(n4160 ,n3460 ,n4069);
    or g890(n4159 ,n3459 ,n4068);
    or g891(n4158 ,n3458 ,n4067);
    or g892(n4157 ,n3457 ,n4066);
    or g893(n4156 ,n3456 ,n4065);
    or g894(n4155 ,n3455 ,n4064);
    or g895(n4154 ,n3454 ,n4063);
    or g896(n4153 ,n3453 ,n4062);
    or g897(n4152 ,n3451 ,n4060);
    or g898(n4151 ,n3452 ,n4061);
    or g899(n4150 ,n3450 ,n4059);
    or g900(n4149 ,n3449 ,n4058);
    or g901(n4148 ,n3448 ,n4057);
    or g902(n4147 ,n3447 ,n4056);
    or g903(n4146 ,n3446 ,n4103);
    or g904(n4145 ,n3611 ,n4003);
    or g905(n4144 ,n3612 ,n4005);
    or g906(n4143 ,n3613 ,n4007);
    or g907(n4142 ,n3614 ,n4009);
    or g908(n4141 ,n3615 ,n4011);
    or g909(n4140 ,n3616 ,n4013);
    or g910(n4139 ,n3617 ,n4015);
    or g911(n4138 ,n2589 ,n3990);
    or g912(n4137 ,n2592 ,n4053);
    or g913(n4136 ,n2403 ,n4051);
    or g914(n4135 ,n2596 ,n4052);
    or g915(n4134 ,n2603 ,n4050);
    or g916(n4133 ,n2606 ,n4049);
    or g917(n4132 ,n2608 ,n4048);
    or g918(n4131 ,n2613 ,n4046);
    or g919(n4130 ,n2400 ,n4047);
    or g920(n4129 ,n2424 ,n4045);
    or g921(n4128 ,n2441 ,n4044);
    or g922(n4127 ,n2444 ,n4043);
    or g923(n4126 ,n2585 ,n4042);
    or g924(n4125 ,n2395 ,n4041);
    or g925(n4124 ,n2604 ,n4040);
    or g926(n4123 ,n2393 ,n4039);
    or g927(n4122 ,n2609 ,n4038);
    or g928(n4121 ,n2407 ,n4037);
    or g929(n4120 ,n2387 ,n4035);
    or g930(n4119 ,n2388 ,n4036);
    or g931(n4118 ,n2583 ,n4034);
    or g932(n4117 ,n2422 ,n4033);
    or g933(n4116 ,n2601 ,n4032);
    or g934(n4115 ,n2383 ,n4031);
    or g935(n4114 ,n2607 ,n4030);
    or g936(n4113 ,n2396 ,n4029);
    or g937(n4112 ,n2595 ,n4028);
    or g938(n4111 ,n2401 ,n4027);
    or g939(n4110 ,n2456 ,n4025);
    or g940(n4109 ,n2380 ,n4026);
    or g941(n4108 ,n2588 ,n4024);
    or g942(n4107 ,n2378 ,n4023);
    or g943(n4106 ,n3620 ,n4022);
    or g944(n4105 ,n3619 ,n4020);
    or g945(n4104 ,n3618 ,n4017);
    or g946(n4103 ,n1848 ,n3989);
    or g947(n4102 ,n3631 ,n3999);
    or g948(n4101 ,n3653 ,n3997);
    or g949(n4100 ,n3602 ,n3993);
    or g950(n4099 ,n3601 ,n3991);
    or g951(n4098 ,n3582 ,n3995);
    or g952(n4097 ,n3600 ,n3925);
    or g953(n4096 ,n3599 ,n3987);
    or g954(n4095 ,n3598 ,n3985);
    or g955(n4094 ,n3597 ,n3981);
    or g956(n4093 ,n3596 ,n3982);
    or g957(n4092 ,n3595 ,n3979);
    or g958(n4091 ,n3594 ,n3977);
    or g959(n4090 ,n3593 ,n3975);
    or g960(n4089 ,n3592 ,n3973);
    or g961(n4088 ,n3591 ,n3971);
    or g962(n4087 ,n3590 ,n3970);
    or g963(n4086 ,n3589 ,n3967);
    or g964(n4085 ,n3588 ,n3965);
    or g965(n4084 ,n3587 ,n3963);
    or g966(n4083 ,n3586 ,n3961);
    or g967(n4082 ,n3585 ,n3959);
    or g968(n4081 ,n3706 ,n3952);
    or g969(n4080 ,n1852 ,n3950);
    or g970(n4079 ,n1842 ,n3949);
    or g971(n4078 ,n1841 ,n3948);
    or g972(n4077 ,n1840 ,n3947);
    or g973(n4076 ,n1827 ,n3946);
    or g974(n4075 ,n1851 ,n3944);
    or g975(n4074 ,n1845 ,n3945);
    or g976(n4073 ,n1838 ,n3943);
    or g977(n4072 ,n1850 ,n3942);
    or g978(n4071 ,n1836 ,n3941);
    or g979(n4070 ,n1849 ,n3940);
    or g980(n4069 ,n1847 ,n3939);
    or g981(n4068 ,n1835 ,n3938);
    or g982(n4067 ,n1834 ,n3937);
    or g983(n4066 ,n1829 ,n3936);
    or g984(n4065 ,n1833 ,n3935);
    or g985(n4064 ,n1832 ,n3934);
    or g986(n4063 ,n1837 ,n3933);
    or g987(n4062 ,n1843 ,n3932);
    or g988(n4061 ,n1844 ,n3931);
    or g989(n4060 ,n1828 ,n3930);
    or g990(n4059 ,n1830 ,n3929);
    or g991(n4058 ,n1831 ,n3928);
    or g992(n4057 ,n1839 ,n3927);
    or g993(n4056 ,n1846 ,n3926);
    or g994(n4055 ,n3610 ,n4001);
    or g995(n4054 ,n3855 ,n3854);
    or g996(n4053 ,n2593 ,n3761);
    or g997(n4052 ,n2404 ,n3760);
    or g998(n4051 ,n2602 ,n3759);
    or g999(n4050 ,n2402 ,n3758);
    or g1000(n4049 ,n2610 ,n3757);
    or g1001(n4048 ,n2614 ,n3756);
    or g1002(n4047 ,n2612 ,n3755);
    or g1003(n4046 ,n2399 ,n3754);
    or g1004(n4045 ,n2462 ,n3753);
    or g1005(n4044 ,n2429 ,n3752);
    or g1006(n4043 ,n2459 ,n3751);
    or g1007(n4042 ,n2397 ,n3750);
    or g1008(n4041 ,n2591 ,n3749);
    or g1009(n4040 ,n2598 ,n3748);
    or g1010(n4039 ,n2605 ,n3747);
    or g1011(n4038 ,n2392 ,n3746);
    or g1012(n4037 ,n2377 ,n3744);
    or g1013(n4036 ,n2594 ,n3743);
    or g1014(n4035 ,n2390 ,n3745);
    or g1015(n4034 ,n2386 ,n3742);
    or g1016(n4033 ,n2434 ,n3741);
    or g1017(n4032 ,n2586 ,n3740);
    or g1018(n4031 ,n2597 ,n3739);
    or g1019(n4030 ,n2611 ,n3738);
    or g1020(n4029 ,n2382 ,n3737);
    or g1021(n4028 ,n2394 ,n3736);
    or g1022(n4027 ,n2461 ,n3735);
    or g1023(n4026 ,n2428 ,n3733);
    or g1024(n4025 ,n2381 ,n3734);
    or g1025(n4024 ,n2587 ,n3732);
    or g1026(n4023 ,n2600 ,n3828);
    or g1027(n4022 ,n3917 ,n3913);
    or g1028(n4021 ,n3916 ,n3915);
    or g1029(n4020 ,n3914 ,n3912);
    or g1030(n4019 ,n3919 ,n3918);
    or g1031(n4018 ,n3911 ,n3910);
    or g1032(n4017 ,n3909 ,n3908);
    or g1033(n4016 ,n3906 ,n3907);
    or g1034(n4015 ,n3904 ,n3905);
    or g1035(n4014 ,n3903 ,n3902);
    or g1036(n4013 ,n3901 ,n3900);
    or g1037(n4012 ,n3897 ,n3899);
    or g1038(n4011 ,n3898 ,n3896);
    or g1039(n4010 ,n3895 ,n3894);
    or g1040(n4009 ,n3893 ,n3892);
    or g1041(n4008 ,n3890 ,n3891);
    or g1042(n4007 ,n3889 ,n3888);
    or g1043(n4006 ,n3887 ,n3886);
    or g1044(n4005 ,n3885 ,n3884);
    or g1045(n4004 ,n3883 ,n3882);
    or g1046(n4003 ,n3881 ,n3880);
    or g1047(n4002 ,n3878 ,n3879);
    or g1048(n4001 ,n3877 ,n3924);
    or g1049(n4000 ,n3874 ,n3875);
    or g1050(n3999 ,n3873 ,n3872);
    or g1051(n3998 ,n3871 ,n3870);
    or g1052(n3997 ,n3869 ,n3868);
    or g1053(n3996 ,n3862 ,n3865);
    or g1054(n3995 ,n3867 ,n3866);
    or g1055(n3994 ,n3864 ,n3863);
    or g1056(n3993 ,n3861 ,n3860);
    or g1057(n3992 ,n3858 ,n3859);
    or g1058(n3991 ,n3857 ,n3856);
    or g1059(n3990 ,n2590 ,n3762);
    or g1060(n3989 ,n3765 ,n3691);
    or g1061(n3988 ,n3851 ,n3850);
    or g1062(n3987 ,n3849 ,n3848);
    or g1063(n3986 ,n3847 ,n3846);
    or g1064(n3985 ,n3845 ,n3844);
    or g1065(n3984 ,n3842 ,n3843);
    or g1066(n3983 ,n3839 ,n3838);
    or g1067(n3982 ,n3837 ,n3836);
    or g1068(n3981 ,n3841 ,n3840);
    or g1069(n3980 ,n3833 ,n3835);
    or g1070(n3979 ,n3834 ,n3832);
    or g1071(n3978 ,n3831 ,n3830);
    or g1072(n3977 ,n3829 ,n3731);
    or g1073(n3976 ,n3826 ,n3827);
    or g1074(n3975 ,n3825 ,n3824);
    or g1075(n3974 ,n3823 ,n3822);
    or g1076(n3973 ,n3821 ,n3820);
    or g1077(n3972 ,n3819 ,n3818);
    or g1078(n3971 ,n3817 ,n3816);
    or g1079(n3970 ,n3813 ,n3812);
    or g1080(n3969 ,n3810 ,n3811);
    or g1081(n3968 ,n3815 ,n3814);
    or g1082(n3967 ,n3809 ,n3808);
    or g1083(n3966 ,n3807 ,n3806);
    or g1084(n3965 ,n3805 ,n3804);
    or g1085(n3964 ,n3803 ,n3801);
    or g1086(n3963 ,n3802 ,n3800);
    or g1087(n3962 ,n3799 ,n3798);
    or g1088(n3961 ,n3797 ,n3796);
    or g1089(n3960 ,n3794 ,n3795);
    or g1090(n3959 ,n3793 ,n3792);
    or g1091(n3958 ,n3713 ,n3764);
    or g1092(n3957 ,n3712 ,n3763);
    or g1093(n3956 ,n3710 ,n3876);
    or g1094(n3955 ,n3709 ,n3923);
    or g1095(n3954 ,n3708 ,n3922);
    or g1096(n3953 ,n3730 ,n3920);
    or g1097(n3952 ,n1800 ,n3791);
    or g1098(n3951 ,n3711 ,n3921);
    or g1099(n3950 ,n3790 ,n3705);
    or g1100(n3949 ,n3789 ,n3704);
    or g1101(n3948 ,n3788 ,n3703);
    or g1102(n3947 ,n3787 ,n3702);
    or g1103(n3946 ,n3786 ,n3707);
    or g1104(n3945 ,n3784 ,n3715);
    or g1105(n3944 ,n3785 ,n3714);
    or g1106(n3943 ,n3783 ,n3716);
    or g1107(n3942 ,n3782 ,n3717);
    or g1108(n3941 ,n3781 ,n3718);
    or g1109(n3940 ,n3780 ,n3719);
    or g1110(n3939 ,n3779 ,n3720);
    or g1111(n3938 ,n3778 ,n3721);
    or g1112(n3937 ,n3777 ,n3722);
    or g1113(n3936 ,n3776 ,n3723);
    or g1114(n3935 ,n3775 ,n3724);
    or g1115(n3934 ,n3774 ,n3725);
    or g1116(n3933 ,n3773 ,n3726);
    or g1117(n3932 ,n3772 ,n3727);
    or g1118(n3931 ,n3771 ,n3728);
    or g1119(n3930 ,n3770 ,n3729);
    or g1120(n3929 ,n3769 ,n3672);
    or g1121(n3928 ,n3768 ,n3694);
    or g1122(n3927 ,n3767 ,n3693);
    or g1123(n3926 ,n3766 ,n3692);
    or g1124(n3925 ,n3852 ,n3853);
    nor g1125(n3924 ,n1387 ,n3699);
    nor g1126(n3923 ,n1123 ,n3701);
    nor g1127(n3922 ,n1076 ,n3701);
    nor g1128(n3921 ,n1171 ,n3701);
    nor g1129(n3920 ,n1021 ,n3701);
    nor g1130(n3919 ,n1333 ,n3696);
    nor g1131(n3918 ,n1366 ,n3697);
    nor g1132(n3917 ,n1324 ,n3698);
    nor g1133(n3916 ,n946 ,n3696);
    nor g1134(n3915 ,n1393 ,n3697);
    nor g1135(n3914 ,n955 ,n3698);
    nor g1136(n3913 ,n958 ,n3699);
    nor g1137(n3912 ,n1392 ,n3699);
    nor g1138(n3911 ,n963 ,n3696);
    nor g1139(n3910 ,n1340 ,n3697);
    nor g1140(n3909 ,n947 ,n3698);
    nor g1141(n3908 ,n1326 ,n3699);
    nor g1142(n3907 ,n1354 ,n3697);
    nor g1143(n3906 ,n1329 ,n3696);
    nor g1144(n3905 ,n1388 ,n3699);
    nor g1145(n3904 ,n1391 ,n3698);
    nor g1146(n3903 ,n1394 ,n3696);
    nor g1147(n3902 ,n1309 ,n3697);
    nor g1148(n3901 ,n1318 ,n3698);
    nor g1149(n3900 ,n944 ,n3699);
    nor g1150(n3899 ,n1389 ,n3697);
    nor g1151(n3898 ,n1363 ,n3698);
    nor g1152(n3897 ,n1368 ,n3696);
    nor g1153(n3896 ,n937 ,n3699);
    nor g1154(n3895 ,n1314 ,n3696);
    nor g1155(n3894 ,n1315 ,n3697);
    nor g1156(n3893 ,n1379 ,n3698);
    nor g1157(n3892 ,n1383 ,n3699);
    nor g1158(n3891 ,n1370 ,n3697);
    nor g1159(n3890 ,n1325 ,n3696);
    nor g1160(n3889 ,n1362 ,n3698);
    nor g1161(n3888 ,n1390 ,n3699);
    nor g1162(n3887 ,n1372 ,n3696);
    nor g1163(n3886 ,n960 ,n3697);
    nor g1164(n3885 ,n1381 ,n3698);
    nor g1165(n3884 ,n1355 ,n3699);
    nor g1166(n3883 ,n1360 ,n3696);
    nor g1167(n3882 ,n1319 ,n3697);
    nor g1168(n3881 ,n1395 ,n3698);
    nor g1169(n3880 ,n1384 ,n3699);
    nor g1170(n3879 ,n1346 ,n3697);
    nor g1171(n3878 ,n1403 ,n3696);
    nor g1172(n3877 ,n1300 ,n3698);
    nor g1173(n3876 ,n1052 ,n3701);
    nor g1174(n3875 ,n1308 ,n3697);
    nor g1175(n3874 ,n1358 ,n3696);
    nor g1176(n3873 ,n1356 ,n3698);
    nor g1177(n3872 ,n1353 ,n3699);
    nor g1178(n3871 ,n948 ,n3696);
    nor g1179(n3870 ,n1334 ,n3697);
    nor g1180(n3869 ,n1331 ,n3698);
    nor g1181(n3868 ,n950 ,n3699);
    nor g1182(n3867 ,n959 ,n3698);
    nor g1183(n3866 ,n1357 ,n3699);
    nor g1184(n3865 ,n1316 ,n3697);
    nor g1185(n3864 ,n957 ,n3696);
    nor g1186(n3863 ,n1382 ,n3697);
    nor g1187(n3862 ,n1408 ,n3696);
    nor g1188(n3861 ,n1361 ,n3698);
    nor g1189(n3860 ,n1307 ,n3699);
    nor g1190(n3859 ,n962 ,n3697);
    nor g1191(n3858 ,n1407 ,n3696);
    nor g1192(n3857 ,n1349 ,n3698);
    nor g1193(n3856 ,n961 ,n3699);
    nor g1194(n3855 ,n1298 ,n3696);
    nor g1195(n3854 ,n1375 ,n3697);
    nor g1196(n3853 ,n941 ,n3699);
    nor g1197(n3852 ,n1398 ,n3698);
    nor g1198(n3851 ,n1320 ,n3696);
    nor g1199(n3850 ,n1378 ,n3697);
    nor g1200(n3849 ,n1376 ,n3698);
    nor g1201(n3848 ,n1338 ,n3699);
    nor g1202(n3847 ,n1385 ,n3696);
    nor g1203(n3846 ,n952 ,n3697);
    nor g1204(n3845 ,n945 ,n3698);
    nor g1205(n3844 ,n1351 ,n3699);
    nor g1206(n3843 ,n1406 ,n3697);
    nor g1207(n3842 ,n1374 ,n3696);
    nor g1208(n3841 ,n1310 ,n3698);
    nor g1209(n3840 ,n1303 ,n3699);
    nor g1210(n3839 ,n1328 ,n3696);
    nor g1211(n3838 ,n1339 ,n3697);
    nor g1212(n3837 ,n1321 ,n3698);
    nor g1213(n3836 ,n1342 ,n3699);
    nor g1214(n3835 ,n954 ,n3697);
    nor g1215(n3834 ,n1317 ,n3698);
    nor g1216(n3833 ,n939 ,n3696);
    nor g1217(n3832 ,n1359 ,n3699);
    nor g1218(n3831 ,n1337 ,n3696);
    nor g1219(n3830 ,n1347 ,n3697);
    nor g1220(n3829 ,n1344 ,n3698);
    or g1221(n3828 ,n3621 ,n3659);
    nor g1222(n3827 ,n1386 ,n3697);
    nor g1223(n3826 ,n1373 ,n3696);
    nor g1224(n3825 ,n1302 ,n3698);
    nor g1225(n3824 ,n1330 ,n3699);
    nor g1226(n3823 ,n1404 ,n3696);
    nor g1227(n3822 ,n1350 ,n3697);
    nor g1228(n3821 ,n1367 ,n3698);
    nor g1229(n3820 ,n965 ,n3699);
    nor g1230(n3819 ,n1364 ,n3696);
    nor g1231(n3818 ,n964 ,n3697);
    nor g1232(n3817 ,n956 ,n3698);
    nor g1233(n3816 ,n1313 ,n3699);
    nor g1234(n3815 ,n1371 ,n3696);
    nor g1235(n3814 ,n1365 ,n3697);
    nor g1236(n3813 ,n940 ,n3698);
    nor g1237(n3812 ,n1409 ,n3699);
    nor g1238(n3811 ,n1352 ,n3697);
    nor g1239(n3810 ,n1402 ,n3696);
    nor g1240(n3809 ,n1336 ,n3698);
    nor g1241(n3808 ,n1322 ,n3699);
    nor g1242(n3807 ,n1399 ,n3696);
    nor g1243(n3806 ,n1312 ,n3697);
    nor g1244(n3805 ,n1400 ,n3698);
    nor g1245(n3804 ,n1332 ,n3699);
    nor g1246(n3803 ,n1323 ,n3696);
    nor g1247(n3802 ,n1405 ,n3698);
    nor g1248(n3801 ,n938 ,n3697);
    nor g1249(n3800 ,n936 ,n3699);
    nor g1250(n3799 ,n942 ,n3696);
    nor g1251(n3798 ,n1306 ,n3697);
    nor g1252(n3797 ,n1345 ,n3698);
    nor g1253(n3796 ,n1369 ,n3699);
    nor g1254(n3795 ,n966 ,n3697);
    nor g1255(n3794 ,n1397 ,n3696);
    nor g1256(n3793 ,n1305 ,n3698);
    nor g1257(n3792 ,n1327 ,n3699);
    nor g1258(n3791 ,n844 ,n3658);
    nor g1259(n3790 ,n861 ,n3700);
    nor g1260(n3789 ,n847 ,n3700);
    nor g1261(n3788 ,n862 ,n3700);
    nor g1262(n3787 ,n854 ,n3700);
    nor g1263(n3786 ,n851 ,n3700);
    nor g1264(n3785 ,n846 ,n3700);
    nor g1265(n3784 ,n849 ,n3700);
    nor g1266(n3783 ,n859 ,n3700);
    nor g1267(n3782 ,n860 ,n3700);
    nor g1268(n3781 ,n853 ,n3700);
    nor g1269(n3780 ,n867 ,n3700);
    nor g1270(n3779 ,n845 ,n3700);
    nor g1271(n3778 ,n863 ,n3700);
    nor g1272(n3777 ,n858 ,n3700);
    nor g1273(n3776 ,n848 ,n3700);
    nor g1274(n3775 ,n850 ,n3700);
    nor g1275(n3774 ,n865 ,n3700);
    nor g1276(n3773 ,n855 ,n3700);
    nor g1277(n3772 ,n864 ,n3700);
    nor g1278(n3771 ,n869 ,n3700);
    nor g1279(n3770 ,n868 ,n3700);
    nor g1280(n3769 ,n852 ,n3700);
    nor g1281(n3768 ,n866 ,n3700);
    nor g1282(n3767 ,n857 ,n3700);
    nor g1283(n3766 ,n870 ,n3700);
    nor g1284(n3765 ,n856 ,n3700);
    nor g1285(n3764 ,n799 ,n3655);
    nor g1286(n3763 ,n814 ,n3656);
    or g1287(n3762 ,n3651 ,n3690);
    or g1288(n3761 ,n3650 ,n3689);
    or g1289(n3760 ,n3649 ,n3688);
    or g1290(n3759 ,n3648 ,n3687);
    or g1291(n3758 ,n3647 ,n3686);
    or g1292(n3757 ,n3646 ,n3685);
    or g1293(n3756 ,n3645 ,n3684);
    or g1294(n3755 ,n3644 ,n3683);
    or g1295(n3754 ,n3643 ,n3682);
    or g1296(n3753 ,n3642 ,n3681);
    or g1297(n3752 ,n3641 ,n3680);
    or g1298(n3751 ,n3640 ,n3679);
    or g1299(n3750 ,n3639 ,n3678);
    or g1300(n3749 ,n3638 ,n3677);
    or g1301(n3748 ,n3637 ,n3676);
    or g1302(n3747 ,n3636 ,n3675);
    or g1303(n3746 ,n3635 ,n3674);
    or g1304(n3745 ,n3633 ,n3695);
    or g1305(n3744 ,n3634 ,n3673);
    or g1306(n3743 ,n3632 ,n3671);
    or g1307(n3742 ,n3654 ,n3670);
    or g1308(n3741 ,n3630 ,n3669);
    or g1309(n3740 ,n3629 ,n3668);
    or g1310(n3739 ,n3628 ,n3667);
    or g1311(n3738 ,n3627 ,n3666);
    or g1312(n3737 ,n3626 ,n3665);
    or g1313(n3736 ,n3625 ,n3664);
    or g1314(n3735 ,n3624 ,n3663);
    or g1315(n3734 ,n3623 ,n3662);
    or g1316(n3733 ,n3622 ,n3661);
    or g1317(n3732 ,n3652 ,n3660);
    nor g1318(n3731 ,n1311 ,n3699);
    nor g1319(n3730 ,n1573 ,n3604);
    nor g1320(n3729 ,n1557 ,n3604);
    nor g1321(n3728 ,n1511 ,n3604);
    nor g1322(n3727 ,n1568 ,n3604);
    nor g1323(n3726 ,n1537 ,n3604);
    nor g1324(n3725 ,n1522 ,n3604);
    nor g1325(n3724 ,n980 ,n3604);
    nor g1326(n3723 ,n1473 ,n3604);
    nor g1327(n3722 ,n990 ,n3604);
    nor g1328(n3721 ,n1575 ,n3604);
    nor g1329(n3720 ,n1452 ,n3604);
    nor g1330(n3719 ,n1534 ,n3604);
    nor g1331(n3718 ,n993 ,n3604);
    nor g1332(n3717 ,n1416 ,n3604);
    nor g1333(n3716 ,n1561 ,n3604);
    nor g1334(n3715 ,n1445 ,n3604);
    nor g1335(n3714 ,n1483 ,n3604);
    nor g1336(n3713 ,n1524 ,n3607);
    nor g1337(n3712 ,n1474 ,n3609);
    nor g1338(n3711 ,n1493 ,n3604);
    nor g1339(n3710 ,n1472 ,n3604);
    nor g1340(n3709 ,n1476 ,n3604);
    nor g1341(n3708 ,n1533 ,n3604);
    nor g1342(n3707 ,n1442 ,n3604);
    nor g1343(n3706 ,n1540 ,n3604);
    nor g1344(n3705 ,n1531 ,n3604);
    nor g1345(n3704 ,n1579 ,n3604);
    nor g1346(n3703 ,n1585 ,n3604);
    nor g1347(n3702 ,n979 ,n3604);
    nor g1348(n3695 ,n1512 ,n3605);
    nor g1349(n3694 ,n1574 ,n3604);
    nor g1350(n3693 ,n1008 ,n3604);
    nor g1351(n3692 ,n1432 ,n3604);
    nor g1352(n3691 ,n1469 ,n3604);
    nor g1353(n3690 ,n1502 ,n3605);
    nor g1354(n3689 ,n1470 ,n3605);
    nor g1355(n3688 ,n1419 ,n3605);
    nor g1356(n3687 ,n1551 ,n3605);
    nor g1357(n3686 ,n988 ,n3605);
    nor g1358(n3685 ,n1517 ,n3605);
    nor g1359(n3684 ,n1556 ,n3605);
    nor g1360(n3683 ,n1446 ,n3605);
    nor g1361(n3682 ,n1589 ,n3605);
    nor g1362(n3681 ,n1436 ,n3605);
    nor g1363(n3680 ,n1499 ,n3605);
    nor g1364(n3679 ,n1459 ,n3605);
    nor g1365(n3678 ,n1480 ,n3605);
    nor g1366(n3677 ,n1015 ,n3605);
    nor g1367(n3676 ,n1563 ,n3605);
    nor g1368(n3675 ,n1447 ,n3605);
    nor g1369(n3674 ,n1503 ,n3605);
    nor g1370(n3673 ,n996 ,n3605);
    nor g1371(n3672 ,n1560 ,n3604);
    nor g1372(n3671 ,n1542 ,n3605);
    nor g1373(n3670 ,n1451 ,n3605);
    nor g1374(n3669 ,n1494 ,n3605);
    nor g1375(n3668 ,n1462 ,n3605);
    nor g1376(n3667 ,n1544 ,n3605);
    nor g1377(n3666 ,n976 ,n3605);
    nor g1378(n3665 ,n1433 ,n3605);
    nor g1379(n3664 ,n1013 ,n3605);
    nor g1380(n3663 ,n1586 ,n3605);
    nor g1381(n3662 ,n1007 ,n3605);
    nor g1382(n3661 ,n1420 ,n3605);
    nor g1383(n3660 ,n1530 ,n3605);
    nor g1384(n3659 ,n1508 ,n3605);
    or g1385(n3658 ,n1764 ,n3603);
    nor g1386(n3657 ,n811 ,n3584);
    or g1387(n3656 ,n1729 ,n3608);
    or g1388(n3655 ,n1729 ,n3606);
    or g1389(n3701 ,n1738 ,n802);
    or g1390(n3700 ,n1716 ,n802);
    or g1391(n3699 ,n6[5] ,n800);
    or g1392(n3698 ,n6[5] ,n801);
    or g1393(n3697 ,n844 ,n800);
    or g1394(n3696 ,n844 ,n801);
    nor g1395(n3654 ,n1043 ,n3564);
    nor g1396(n3653 ,n1564 ,n3563);
    nor g1397(n3652 ,n1163 ,n3564);
    nor g1398(n3651 ,n1151 ,n3564);
    nor g1399(n3650 ,n1116 ,n3564);
    nor g1400(n3649 ,n1173 ,n3564);
    nor g1401(n3648 ,n1203 ,n3564);
    nor g1402(n3647 ,n1090 ,n3564);
    nor g1403(n3646 ,n1053 ,n3564);
    nor g1404(n3645 ,n1162 ,n3564);
    nor g1405(n3644 ,n1048 ,n3564);
    nor g1406(n3643 ,n1078 ,n3564);
    nor g1407(n3642 ,n1178 ,n3564);
    nor g1408(n3641 ,n1136 ,n3564);
    nor g1409(n3640 ,n1217 ,n3564);
    nor g1410(n3639 ,n1143 ,n3564);
    nor g1411(n3638 ,n1071 ,n3564);
    nor g1412(n3637 ,n1182 ,n3564);
    nor g1413(n3636 ,n1131 ,n3564);
    nor g1414(n3635 ,n1181 ,n3564);
    nor g1415(n3634 ,n1029 ,n3564);
    nor g1416(n3633 ,n1210 ,n3564);
    nor g1417(n3632 ,n1033 ,n3564);
    nor g1418(n3631 ,n1465 ,n3563);
    nor g1419(n3630 ,n1194 ,n3564);
    nor g1420(n3629 ,n1170 ,n3564);
    nor g1421(n3628 ,n1216 ,n3564);
    nor g1422(n3627 ,n1062 ,n3564);
    nor g1423(n3626 ,n1110 ,n3564);
    nor g1424(n3625 ,n1220 ,n3564);
    nor g1425(n3624 ,n1036 ,n3564);
    nor g1426(n3623 ,n1167 ,n3564);
    nor g1427(n3622 ,n1112 ,n3564);
    nor g1428(n3621 ,n1041 ,n3564);
    nor g1429(n3620 ,n1541 ,n3563);
    nor g1430(n3619 ,n989 ,n3563);
    nor g1431(n3618 ,n1566 ,n3563);
    nor g1432(n3617 ,n974 ,n3563);
    nor g1433(n3616 ,n1514 ,n3563);
    nor g1434(n3615 ,n1491 ,n3563);
    nor g1435(n3614 ,n1492 ,n3563);
    nor g1436(n3613 ,n999 ,n3563);
    nor g1437(n3612 ,n1454 ,n3563);
    nor g1438(n3611 ,n1518 ,n3563);
    nor g1439(n3610 ,n1484 ,n3563);
    not g1440(n3609 ,n3608);
    not g1441(n3607 ,n3606);
    not g1442(n3603 ,n3604);
    nor g1443(n3602 ,n1578 ,n3563);
    nor g1444(n3601 ,n1550 ,n3563);
    nor g1445(n3600 ,n969 ,n3563);
    nor g1446(n3599 ,n1440 ,n3563);
    nor g1447(n3598 ,n1536 ,n3563);
    nor g1448(n3597 ,n1457 ,n3563);
    nor g1449(n3596 ,n1538 ,n3563);
    nor g1450(n3595 ,n1455 ,n3563);
    nor g1451(n3594 ,n1545 ,n3563);
    nor g1452(n3593 ,n1562 ,n3563);
    nor g1453(n3592 ,n1581 ,n3563);
    nor g1454(n3591 ,n971 ,n3563);
    nor g1455(n3590 ,n1453 ,n3563);
    nor g1456(n3589 ,n1489 ,n3563);
    nor g1457(n3588 ,n1411 ,n3563);
    nor g1458(n3587 ,n1429 ,n3563);
    nor g1459(n3586 ,n1001 ,n3563);
    nor g1460(n3585 ,n1584 ,n3563);
    nor g1461(n3584 ,n13 ,n3551);
    or g1462(n3583 ,n3482 ,n3539);
    nor g1463(n3582 ,n1571 ,n3563);
    nor g1464(n3581 ,n839 ,n3547);
    nor g1465(n3580 ,n811 ,n3555);
    nor g1466(n3579 ,n811 ,n3554);
    nor g1467(n3578 ,n812 ,n3553);
    nor g1468(n3577 ,n813 ,n3552);
    nor g1469(n3576 ,n841 ,n3560);
    nor g1470(n3575 ,n839 ,n3561);
    nor g1471(n3574 ,n811 ,n3549);
    nor g1472(n3573 ,n839 ,n3540);
    nor g1473(n3572 ,n841 ,n3546);
    nor g1474(n3571 ,n813 ,n3538);
    nor g1475(n3570 ,n811 ,n3545);
    nor g1476(n3569 ,n839 ,n3544);
    nor g1477(n3568 ,n811 ,n3542);
    nor g1478(n3567 ,n810 ,n3543);
    nor g1479(n3566 ,n799 ,n3541);
    nor g1480(n3608 ,n810 ,n3556);
    nor g1481(n3606 ,n839 ,n3557);
    nor g1482(n3605 ,n810 ,n3550);
    nor g1483(n3604 ,n839 ,n3548);
    not g1484(n3562 ,n3563);
    nor g1485(n3561 ,n3514 ,n3525);
    nor g1486(n3560 ,n3515 ,n3520);
    nor g1487(n3559 ,n839 ,n3504);
    nor g1488(n3558 ,n841 ,n3503);
    or g1489(n3557 ,n1730 ,n3536);
    or g1490(n3556 ,n1730 ,n3535);
    nor g1491(n3555 ,n3519 ,n3524);
    nor g1492(n3554 ,n3518 ,n3523);
    nor g1493(n3553 ,n3517 ,n3522);
    nor g1494(n3552 ,n3516 ,n3521);
    nor g1495(n3565 ,n1221 ,n3535);
    or g1496(n3564 ,n814 ,n3534);
    nor g1497(n3563 ,n812 ,n3537);
    not g1498(n3551 ,n3550);
    nor g1499(n3549 ,n3513 ,n3533);
    nor g1500(n3548 ,n1736 ,n3535);
    xnor g1501(n3547 ,n3500 ,n34[0]);
    nor g1502(n3546 ,n3507 ,n3527);
    nor g1503(n3545 ,n3510 ,n3526);
    nor g1504(n3544 ,n3509 ,n3531);
    nor g1505(n3543 ,n3512 ,n3529);
    nor g1506(n3542 ,n3508 ,n3530);
    nor g1507(n3541 ,n3511 ,n3528);
    nor g1508(n3540 ,n3506 ,n3532);
    or g1509(n3539 ,n3445 ,n3505);
    xnor g1510(n3538 ,n3502 ,n35[0]);
    nor g1511(n3550 ,n1733 ,n3535);
    not g1512(n3537 ,n3536);
    not g1513(n3534 ,n3535);
    nor g1514(n3533 ,n1083 ,n3499);
    nor g1515(n3532 ,n1060 ,n3501);
    nor g1516(n3531 ,n1042 ,n3501);
    nor g1517(n3530 ,n1028 ,n3501);
    nor g1518(n3529 ,n1200 ,n3501);
    nor g1519(n3528 ,n1126 ,n3501);
    nor g1520(n3527 ,n1191 ,n3501);
    nor g1521(n3526 ,n1119 ,n3501);
    nor g1522(n3525 ,n1097 ,n3499);
    nor g1523(n3524 ,n1172 ,n3499);
    nor g1524(n3523 ,n1105 ,n3499);
    nor g1525(n3522 ,n1199 ,n3499);
    nor g1526(n3521 ,n1211 ,n3499);
    nor g1527(n3520 ,n1183 ,n3499);
    nor g1528(n3536 ,n978 ,n3499);
    nor g1529(n3535 ,n975 ,n3499);
    nor g1530(n3519 ,n949 ,n3500);
    nor g1531(n3518 ,n1348 ,n3500);
    nor g1532(n3517 ,n1341 ,n3500);
    nor g1533(n3516 ,n1401 ,n3500);
    nor g1534(n3515 ,n953 ,n3500);
    nor g1535(n3514 ,n1396 ,n3500);
    nor g1536(n3513 ,n1380 ,n3500);
    nor g1537(n3512 ,n1304 ,n3502);
    nor g1538(n3511 ,n943 ,n3502);
    nor g1539(n3510 ,n1410 ,n3502);
    nor g1540(n3509 ,n1299 ,n3502);
    nor g1541(n3508 ,n1335 ,n3502);
    nor g1542(n3507 ,n951 ,n3502);
    nor g1543(n3506 ,n1343 ,n3502);
    nor g1544(n3505 ,n3480 ,n3501);
    nor g1545(n3504 ,n16 ,n3500);
    nor g1546(n3503 ,n17 ,n3502);
    not g1547(n3501 ,n3502);
    nor g1548(n3502 ,n1729 ,n3498);
    not g1549(n3499 ,n3500);
    nor g1550(n3500 ,n1729 ,n3497);
    not g1551(n3498 ,n3497);
    nor g1552(n3497 ,n3485 ,n3496);
    or g1553(n3496 ,n3488 ,n3494);
    not g1554(n3495 ,n3494);
    nor g1555(n3494 ,n3493 ,n3490);
    nor g1556(n3493 ,n844 ,n3486);
    or g1557(n3492 ,n3483 ,n3489);
    or g1558(n3491 ,n3484 ,n3487);
    nor g1559(n3490 ,n6[5] ,n3472);
    nor g1560(n3489 ,n1731 ,n3480);
    nor g1561(n3488 ,n6[5] ,n3474);
    nor g1562(n3487 ,n1735 ,n3480);
    nor g1563(n3486 ,n1756 ,n3473);
    nor g1564(n3485 ,n844 ,n3475);
    nor g1565(n3484 ,n1528 ,n3481);
    nor g1566(n3483 ,n1546 ,n3481);
    nor g1567(n3482 ,n1003 ,n3481);
    not g1568(n3480 ,n3481);
    or g1569(n3479 ,n2925 ,n2696);
    or g1570(n3478 ,n2927 ,n2697);
    or g1571(n3477 ,n2928 ,n2698);
    or g1572(n3476 ,n2929 ,n3079);
    or g1573(n3475 ,n1887 ,n2726);
    or g1574(n3474 ,n1886 ,n2725);
    or g1575(n3473 ,n1859 ,n2909);
    nor g1576(n3472 ,n1883 ,n2724);
    or g1577(n3471 ,n2458 ,n2457);
    or g1578(n3470 ,n2454 ,n2453);
    or g1579(n3469 ,n2452 ,n2451);
    or g1580(n3468 ,n2450 ,n2449);
    or g1581(n3467 ,n2446 ,n2445);
    or g1582(n3466 ,n2443 ,n2442);
    or g1583(n3465 ,n2440 ,n2439);
    or g1584(n3464 ,n2437 ,n2436);
    or g1585(n3463 ,n2433 ,n2432);
    or g1586(n3462 ,n2431 ,n2430);
    or g1587(n3461 ,n2599 ,n2427);
    or g1588(n3460 ,n2426 ,n2425);
    or g1589(n3459 ,n2385 ,n2423);
    or g1590(n3458 ,n2421 ,n2420);
    or g1591(n3457 ,n2419 ,n2418);
    or g1592(n3456 ,n2384 ,n2417);
    or g1593(n3455 ,n2416 ,n2405);
    or g1594(n3454 ,n2411 ,n2415);
    or g1595(n3453 ,n2435 ,n2455);
    or g1596(n3452 ,n2391 ,n2413);
    or g1597(n3451 ,n2375 ,n2376);
    or g1598(n3450 ,n2389 ,n2412);
    or g1599(n3449 ,n2398 ,n2410);
    or g1600(n3448 ,n2414 ,n2408);
    or g1601(n3447 ,n2438 ,n2460);
    or g1602(n3446 ,n2584 ,n2406);
    nor g1603(n3445 ,n1766 ,n2730);
    nor g1604(n3444 ,n810 ,n2374);
    nor g1605(n3443 ,n799 ,n2582);
    nor g1606(n3442 ,n810 ,n2581);
    nor g1607(n3441 ,n811 ,n2580);
    nor g1608(n3440 ,n811 ,n2578);
    nor g1609(n3439 ,n810 ,n2577);
    nor g1610(n3438 ,n810 ,n2575);
    nor g1611(n3437 ,n813 ,n2576);
    nor g1612(n3436 ,n810 ,n2574);
    nor g1613(n3435 ,n810 ,n2573);
    nor g1614(n3434 ,n810 ,n2572);
    nor g1615(n3433 ,n812 ,n2571);
    nor g1616(n3432 ,n812 ,n2569);
    nor g1617(n3431 ,n811 ,n2568);
    nor g1618(n3430 ,n812 ,n2567);
    nor g1619(n3429 ,n812 ,n2566);
    nor g1620(n3428 ,n841 ,n2565);
    nor g1621(n3427 ,n841 ,n2564);
    nor g1622(n3426 ,n812 ,n2562);
    nor g1623(n3425 ,n812 ,n2561);
    nor g1624(n3424 ,n810 ,n2560);
    nor g1625(n3423 ,n810 ,n2558);
    nor g1626(n3422 ,n811 ,n2557);
    nor g1627(n3421 ,n810 ,n2556);
    nor g1628(n3420 ,n812 ,n2555);
    nor g1629(n3419 ,n799 ,n2554);
    nor g1630(n3418 ,n839 ,n2553);
    nor g1631(n3417 ,n839 ,n2552);
    nor g1632(n3416 ,n799 ,n2551);
    nor g1633(n3415 ,n810 ,n2550);
    nor g1634(n3414 ,n839 ,n2549);
    nor g1635(n3413 ,n811 ,n2548);
    nor g1636(n3412 ,n814 ,n2373);
    nor g1637(n3411 ,n839 ,n2547);
    nor g1638(n3410 ,n841 ,n2546);
    nor g1639(n3409 ,n813 ,n2545);
    nor g1640(n3408 ,n812 ,n2544);
    nor g1641(n3407 ,n813 ,n2543);
    nor g1642(n3406 ,n814 ,n2542);
    nor g1643(n3405 ,n813 ,n2541);
    nor g1644(n3404 ,n811 ,n2540);
    nor g1645(n3403 ,n812 ,n2539);
    nor g1646(n3402 ,n811 ,n2538);
    nor g1647(n3401 ,n811 ,n2537);
    nor g1648(n3400 ,n812 ,n2536);
    nor g1649(n3399 ,n810 ,n2535);
    nor g1650(n3398 ,n811 ,n2534);
    nor g1651(n3397 ,n810 ,n2532);
    nor g1652(n3396 ,n810 ,n2531);
    nor g1653(n3395 ,n814 ,n2530);
    nor g1654(n3394 ,n813 ,n2529);
    nor g1655(n3393 ,n813 ,n2527);
    nor g1656(n3392 ,n813 ,n2528);
    nor g1657(n3391 ,n799 ,n2526);
    nor g1658(n3390 ,n813 ,n2525);
    nor g1659(n3389 ,n799 ,n2524);
    nor g1660(n3388 ,n813 ,n2523);
    nor g1661(n3387 ,n799 ,n2522);
    nor g1662(n3386 ,n812 ,n2521);
    nor g1663(n3385 ,n812 ,n2520);
    nor g1664(n3384 ,n799 ,n2570);
    nor g1665(n3383 ,n813 ,n2519);
    nor g1666(n3382 ,n813 ,n2518);
    nor g1667(n3381 ,n814 ,n2517);
    nor g1668(n3380 ,n811 ,n2372);
    nor g1669(n3379 ,n810 ,n2516);
    nor g1670(n3378 ,n811 ,n2515);
    nor g1671(n3377 ,n811 ,n2514);
    nor g1672(n3376 ,n812 ,n2513);
    nor g1673(n3375 ,n811 ,n2512);
    nor g1674(n3374 ,n812 ,n2511);
    nor g1675(n3373 ,n812 ,n2510);
    nor g1676(n3372 ,n811 ,n2509);
    nor g1677(n3371 ,n811 ,n2508);
    nor g1678(n3370 ,n813 ,n2507);
    nor g1679(n3369 ,n811 ,n2506);
    nor g1680(n3368 ,n841 ,n2505);
    nor g1681(n3367 ,n841 ,n2504);
    nor g1682(n3366 ,n814 ,n2503);
    nor g1683(n3365 ,n812 ,n2502);
    nor g1684(n3364 ,n799 ,n2501);
    nor g1685(n3363 ,n841 ,n2500);
    nor g1686(n3362 ,n810 ,n2499);
    nor g1687(n3361 ,n810 ,n2498);
    nor g1688(n3360 ,n814 ,n2448);
    nor g1689(n3359 ,n814 ,n2497);
    nor g1690(n3358 ,n841 ,n2496);
    nor g1691(n3357 ,n812 ,n2495);
    nor g1692(n3356 ,n813 ,n2533);
    nor g1693(n3355 ,n841 ,n2494);
    nor g1694(n3354 ,n811 ,n2493);
    nor g1695(n3353 ,n810 ,n2492);
    nor g1696(n3352 ,n811 ,n2563);
    nor g1697(n3351 ,n799 ,n2491);
    nor g1698(n3350 ,n841 ,n2490);
    nor g1699(n3349 ,n810 ,n2489);
    nor g1700(n3348 ,n811 ,n2729);
    nor g1701(n3347 ,n813 ,n2488);
    nor g1702(n3346 ,n811 ,n2487);
    nor g1703(n3345 ,n812 ,n2486);
    nor g1704(n3344 ,n811 ,n2379);
    nor g1705(n3343 ,n811 ,n2485);
    nor g1706(n3342 ,n813 ,n2484);
    nor g1707(n3341 ,n839 ,n2483);
    nor g1708(n3340 ,n799 ,n2482);
    nor g1709(n3339 ,n813 ,n2481);
    nor g1710(n3338 ,n814 ,n2480);
    nor g1711(n3337 ,n814 ,n2479);
    nor g1712(n3336 ,n814 ,n2478);
    nor g1713(n3335 ,n810 ,n2477);
    nor g1714(n3334 ,n799 ,n2476);
    nor g1715(n3333 ,n813 ,n2475);
    nor g1716(n3332 ,n813 ,n2409);
    nor g1717(n3331 ,n810 ,n2474);
    nor g1718(n3330 ,n812 ,n2472);
    nor g1719(n3329 ,n812 ,n2471);
    nor g1720(n3328 ,n811 ,n2473);
    nor g1721(n3327 ,n813 ,n2470);
    nor g1722(n3326 ,n813 ,n2469);
    nor g1723(n3325 ,n811 ,n2468);
    nor g1724(n3324 ,n814 ,n2447);
    nor g1725(n3323 ,n812 ,n2467);
    nor g1726(n3322 ,n841 ,n2466);
    nor g1727(n3321 ,n814 ,n2465);
    nor g1728(n3320 ,n841 ,n2579);
    nor g1729(n3319 ,n812 ,n2464);
    nor g1730(n3318 ,n841 ,n2559);
    nor g1731(n3317 ,n810 ,n2463);
    or g1732(n3316 ,n2930 ,n2699);
    or g1733(n3315 ,n2959 ,n2721);
    or g1734(n3314 ,n2955 ,n3086);
    or g1735(n3313 ,n2958 ,n2720);
    or g1736(n3312 ,n2957 ,n2719);
    or g1737(n3311 ,n2954 ,n2718);
    or g1738(n3310 ,n2953 ,n2717);
    or g1739(n3309 ,n2956 ,n3087);
    or g1740(n3308 ,n2952 ,n2716);
    or g1741(n3307 ,n2950 ,n3085);
    or g1742(n3306 ,n2951 ,n2715);
    or g1743(n3305 ,n2949 ,n2714);
    or g1744(n3304 ,n2948 ,n2713);
    or g1745(n3303 ,n2947 ,n2712);
    or g1746(n3302 ,n2945 ,n3084);
    or g1747(n3301 ,n2946 ,n2711);
    or g1748(n3300 ,n2944 ,n2710);
    or g1749(n3299 ,n2943 ,n2709);
    or g1750(n3298 ,n2941 ,n2708);
    or g1751(n3297 ,n2942 ,n3083);
    or g1752(n3296 ,n2939 ,n3082);
    or g1753(n3295 ,n2940 ,n2707);
    or g1754(n3294 ,n2938 ,n2706);
    or g1755(n3293 ,n2936 ,n2704);
    or g1756(n3292 ,n2937 ,n3081);
    or g1757(n3291 ,n2935 ,n2703);
    or g1758(n3290 ,n2931 ,n3080);
    or g1759(n3289 ,n2934 ,n2702);
    or g1760(n3288 ,n2933 ,n2701);
    or g1761(n3287 ,n2932 ,n2700);
    nor g1762(n3481 ,n810 ,n2730);
    or g1763(n3286 ,n2727 ,n2722);
    or g1764(n3285 ,n2924 ,n3077);
    or g1765(n3284 ,n2923 ,n3076);
    or g1766(n3283 ,n2922 ,n3075);
    or g1767(n3282 ,n2921 ,n3073);
    or g1768(n3281 ,n2920 ,n3072);
    or g1769(n3280 ,n2914 ,n3066);
    or g1770(n3279 ,n2918 ,n3071);
    or g1771(n3278 ,n2910 ,n3063);
    or g1772(n3277 ,n2916 ,n3070);
    or g1773(n3276 ,n2913 ,n3067);
    or g1774(n3275 ,n2911 ,n3065);
    or g1775(n3274 ,n3088 ,n3064);
    or g1776(n3273 ,n2908 ,n3061);
    or g1777(n3272 ,n2893 ,n3074);
    or g1778(n3271 ,n2907 ,n3062);
    or g1779(n3270 ,n2905 ,n3060);
    or g1780(n3269 ,n2779 ,n2976);
    or g1781(n3268 ,n2903 ,n3058);
    or g1782(n3267 ,n2904 ,n3059);
    or g1783(n3266 ,n2919 ,n3069);
    or g1784(n3265 ,n2901 ,n3057);
    or g1785(n3264 ,n2917 ,n3068);
    or g1786(n3263 ,n2898 ,n3055);
    or g1787(n3262 ,n2900 ,n3056);
    or g1788(n3261 ,n2899 ,n2691);
    or g1789(n3260 ,n2896 ,n3053);
    or g1790(n3259 ,n2780 ,n2654);
    or g1791(n3258 ,n2894 ,n3050);
    or g1792(n3257 ,n2891 ,n3049);
    or g1793(n3256 ,n2890 ,n3052);
    or g1794(n3255 ,n2889 ,n3047);
    or g1795(n3254 ,n2887 ,n3046);
    or g1796(n3253 ,n2888 ,n3048);
    or g1797(n3252 ,n2885 ,n3044);
    or g1798(n3251 ,n2886 ,n3045);
    or g1799(n3250 ,n2884 ,n3043);
    or g1800(n3249 ,n2784 ,n2655);
    or g1801(n3248 ,n2882 ,n3042);
    or g1802(n3247 ,n2883 ,n3041);
    or g1803(n3246 ,n2763 ,n2972);
    or g1804(n3245 ,n2879 ,n3040);
    or g1805(n3244 ,n2878 ,n2657);
    or g1806(n3243 ,n2739 ,n3051);
    or g1807(n3242 ,n2877 ,n3038);
    or g1808(n3241 ,n2876 ,n3036);
    or g1809(n3240 ,n2873 ,n3035);
    or g1810(n3239 ,n2872 ,n3034);
    or g1811(n3238 ,n2871 ,n3032);
    or g1812(n3237 ,n2870 ,n3031);
    or g1813(n3236 ,n2869 ,n3030);
    or g1814(n3235 ,n2868 ,n3027);
    or g1815(n3234 ,n2867 ,n3029);
    or g1816(n3233 ,n2866 ,n3028);
    or g1817(n3232 ,n2865 ,n3026);
    or g1818(n3231 ,n2864 ,n3025);
    or g1819(n3230 ,n2862 ,n3023);
    or g1820(n3229 ,n2863 ,n3024);
    or g1821(n3228 ,n2861 ,n3022);
    or g1822(n3227 ,n2860 ,n3021);
    or g1823(n3226 ,n2859 ,n3020);
    or g1824(n3225 ,n2858 ,n3019);
    or g1825(n3224 ,n2857 ,n3018);
    or g1826(n3223 ,n2856 ,n3017);
    or g1827(n3222 ,n2855 ,n3015);
    or g1828(n3221 ,n2854 ,n3016);
    or g1829(n3220 ,n2853 ,n3014);
    or g1830(n3219 ,n2852 ,n3013);
    or g1831(n3218 ,n2851 ,n3012);
    or g1832(n3217 ,n2850 ,n3011);
    or g1833(n3216 ,n2849 ,n3010);
    or g1834(n3215 ,n2848 ,n3009);
    or g1835(n3214 ,n2847 ,n3008);
    or g1836(n3213 ,n2846 ,n3007);
    or g1837(n3212 ,n2845 ,n3006);
    or g1838(n3211 ,n2844 ,n2966);
    or g1839(n3210 ,n2842 ,n3005);
    or g1840(n3209 ,n2841 ,n3004);
    or g1841(n3208 ,n2840 ,n3002);
    or g1842(n3207 ,n2843 ,n3003);
    or g1843(n3206 ,n2839 ,n3001);
    or g1844(n3205 ,n2837 ,n2999);
    or g1845(n3204 ,n2838 ,n3000);
    or g1846(n3203 ,n2836 ,n2998);
    or g1847(n3202 ,n2833 ,n2997);
    or g1848(n3201 ,n2751 ,n2634);
    or g1849(n3200 ,n2832 ,n2996);
    or g1850(n3199 ,n2831 ,n2995);
    or g1851(n3198 ,n2734 ,n2623);
    or g1852(n3197 ,n2829 ,n2994);
    or g1853(n3196 ,n2752 ,n2969);
    or g1854(n3195 ,n2827 ,n2993);
    or g1855(n3194 ,n2830 ,n2620);
    or g1856(n3193 ,n2789 ,n2622);
    or g1857(n3192 ,n2824 ,n2992);
    or g1858(n3191 ,n2822 ,n2989);
    or g1859(n3190 ,n2823 ,n2991);
    or g1860(n3189 ,n2821 ,n2988);
    or g1861(n3188 ,n2820 ,n2987);
    or g1862(n3187 ,n2818 ,n2986);
    or g1863(n3186 ,n2816 ,n2985);
    or g1864(n3185 ,n2815 ,n2673);
    or g1865(n3184 ,n2813 ,n2672);
    or g1866(n3183 ,n2812 ,n2671);
    or g1867(n3182 ,n2769 ,n2647);
    or g1868(n3181 ,n2808 ,n2982);
    or g1869(n3180 ,n2811 ,n2670);
    or g1870(n3179 ,n2810 ,n2669);
    or g1871(n3178 ,n2814 ,n2983);
    or g1872(n3177 ,n2825 ,n2668);
    or g1873(n3176 ,n2807 ,n2693);
    or g1874(n3175 ,n2805 ,n2667);
    or g1875(n3174 ,n2806 ,n3033);
    or g1876(n3173 ,n2804 ,n2666);
    or g1877(n3172 ,n2802 ,n2981);
    or g1878(n3171 ,n2803 ,n2665);
    or g1879(n3170 ,n2801 ,n2664);
    or g1880(n3169 ,n2771 ,n2984);
    or g1881(n3168 ,n2800 ,n2663);
    or g1882(n3167 ,n2799 ,n2662);
    or g1883(n3166 ,n2798 ,n2661);
    or g1884(n3165 ,n2796 ,n2979);
    or g1885(n3164 ,n2797 ,n2674);
    or g1886(n3163 ,n2793 ,n2980);
    or g1887(n3162 ,n2795 ,n2676);
    or g1888(n3161 ,n2794 ,n2660);
    or g1889(n3160 ,n2792 ,n2659);
    or g1890(n3159 ,n2791 ,n2658);
    or g1891(n3158 ,n2790 ,n2680);
    or g1892(n3157 ,n2788 ,n3037);
    or g1893(n3156 ,n2787 ,n2681);
    or g1894(n3155 ,n2880 ,n2978);
    or g1895(n3154 ,n2817 ,n2990);
    or g1896(n3153 ,n2785 ,n2656);
    or g1897(n3152 ,n2783 ,n2686);
    or g1898(n3151 ,n2897 ,n2977);
    or g1899(n3150 ,n2781 ,n2687);
    or g1900(n3149 ,n2902 ,n2653);
    or g1901(n3148 ,n2778 ,n2689);
    or g1902(n3147 ,n2776 ,n3039);
    or g1903(n3146 ,n2826 ,n2705);
    or g1904(n3145 ,n2777 ,n2652);
    or g1905(n3144 ,n2912 ,n2690);
    or g1906(n3143 ,n2774 ,n2651);
    or g1907(n3142 ,n2775 ,n2975);
    or g1908(n3141 ,n2772 ,n2650);
    or g1909(n3140 ,n2768 ,n2974);
    or g1910(n3139 ,n2834 ,n2649);
    or g1911(n3138 ,n2740 ,n2626);
    or g1912(n3137 ,n2835 ,n2694);
    or g1913(n3136 ,n2770 ,n2648);
    or g1914(n3135 ,n2767 ,n2646);
    or g1915(n3134 ,n2828 ,n2973);
    or g1916(n3133 ,n2766 ,n2679);
    or g1917(n3132 ,n2764 ,n2645);
    or g1918(n3131 ,n2874 ,n2643);
    or g1919(n3130 ,n2762 ,n2684);
    or g1920(n3129 ,n2761 ,n2642);
    or g1921(n3128 ,n2895 ,n2971);
    or g1922(n3127 ,n2760 ,n2641);
    or g1923(n3126 ,n2756 ,n2970);
    or g1924(n3125 ,n2759 ,n2640);
    or g1925(n3124 ,n2758 ,n2639);
    or g1926(n3123 ,n2915 ,n2638);
    or g1927(n3122 ,n2755 ,n2637);
    or g1928(n3121 ,n2742 ,n2636);
    or g1929(n3120 ,n2757 ,n2635);
    or g1930(n3119 ,n2753 ,n2685);
    or g1931(n3118 ,n2749 ,n3054);
    or g1932(n3117 ,n2809 ,n2633);
    or g1933(n3116 ,n2754 ,n2965);
    or g1934(n3115 ,n2748 ,n2632);
    or g1935(n3114 ,n2747 ,n2631);
    or g1936(n3113 ,n2746 ,n2968);
    or g1937(n3112 ,n2881 ,n2682);
    or g1938(n3111 ,n2745 ,n2630);
    or g1939(n3110 ,n2743 ,n2967);
    or g1940(n3109 ,n2773 ,n2688);
    or g1941(n3108 ,n2744 ,n2629);
    or g1942(n3107 ,n2750 ,n2628);
    or g1943(n3106 ,n2741 ,n2627);
    or g1944(n3105 ,n2765 ,n2625);
    or g1945(n3104 ,n2738 ,n2695);
    or g1946(n3103 ,n2782 ,n2964);
    or g1947(n3102 ,n2737 ,n2644);
    or g1948(n3101 ,n2736 ,n2677);
    or g1949(n3100 ,n2875 ,n2963);
    or g1950(n3099 ,n2735 ,n2624);
    or g1951(n3098 ,n2892 ,n2683);
    or g1952(n3097 ,n2733 ,n2692);
    or g1953(n3096 ,n2732 ,n2962);
    or g1954(n3095 ,n2786 ,n2678);
    or g1955(n3094 ,n2906 ,n2961);
    or g1956(n3093 ,n2731 ,n2621);
    or g1957(n3092 ,n2819 ,n2675);
    or g1958(n3091 ,n2723 ,n2960);
    or g1959(n3090 ,n2728 ,n2619);
    or g1960(n3089 ,n2926 ,n3078);
    nor g1961(n3088 ,n1385 ,n827);
    nor g1962(n3087 ,n927 ,n832);
    nor g1963(n3086 ,n885 ,n829);
    nor g1964(n3085 ,n911 ,n829);
    nor g1965(n3084 ,n914 ,n829);
    nor g1966(n3083 ,n933 ,n829);
    nor g1967(n3082 ,n891 ,n2121);
    nor g1968(n3081 ,n930 ,n829);
    nor g1969(n3080 ,n906 ,n829);
    nor g1970(n3079 ,n878 ,n2121);
    nor g1971(n3078 ,n873 ,n829);
    nor g1972(n3077 ,n912 ,n829);
    nor g1973(n3076 ,n922 ,n829);
    nor g1974(n3075 ,n877 ,n829);
    nor g1975(n3074 ,n931 ,n832);
    nor g1976(n3073 ,n889 ,n829);
    nor g1977(n3072 ,n893 ,n2121);
    nor g1978(n3071 ,n932 ,n829);
    nor g1979(n3070 ,n905 ,n829);
    nor g1980(n3069 ,n885 ,n838);
    nor g1981(n3068 ,n911 ,n838);
    nor g1982(n3067 ,n876 ,n829);
    nor g1983(n3066 ,n914 ,n838);
    nor g1984(n3065 ,n915 ,n829);
    nor g1985(n3064 ,n919 ,n829);
    nor g1986(n3063 ,n933 ,n838);
    nor g1987(n3062 ,n904 ,n829);
    nor g1988(n3061 ,n891 ,n2124);
    nor g1989(n3060 ,n896 ,n829);
    nor g1990(n3059 ,n923 ,n829);
    nor g1991(n3058 ,n930 ,n838);
    nor g1992(n3057 ,n910 ,n829);
    nor g1993(n3056 ,n875 ,n829);
    nor g1994(n3055 ,n906 ,n838);
    nor g1995(n3054 ,n896 ,n832);
    nor g1996(n3053 ,n898 ,n2121);
    nor g1997(n3052 ,n878 ,n2124);
    nor g1998(n3051 ,n875 ,n832);
    nor g1999(n3050 ,n879 ,n829);
    nor g2000(n3049 ,n895 ,n829);
    nor g2001(n3048 ,n873 ,n838);
    nor g2002(n3047 ,n931 ,n2121);
    nor g2003(n3046 ,n907 ,n2121);
    nor g2004(n3045 ,n881 ,n829);
    nor g2005(n3044 ,n912 ,n838);
    nor g2006(n3043 ,n883 ,n829);
    nor g2007(n3042 ,n927 ,n829);
    nor g2008(n3041 ,n922 ,n838);
    nor g2009(n3040 ,n877 ,n838);
    nor g2010(n3039 ,n877 ,n2122);
    nor g2011(n3038 ,n889 ,n838);
    nor g2012(n3037 ,n878 ,n832);
    nor g2013(n3036 ,n893 ,n2124);
    nor g2014(n3035 ,n932 ,n838);
    nor g2015(n3034 ,n905 ,n838);
    nor g2016(n3033 ,n914 ,n832);
    nor g2017(n3032 ,n876 ,n838);
    nor g2018(n3031 ,n915 ,n838);
    nor g2019(n3030 ,n919 ,n838);
    nor g2020(n3029 ,n896 ,n838);
    nor g2021(n3028 ,n923 ,n838);
    nor g2022(n3027 ,n904 ,n838);
    nor g2023(n3026 ,n910 ,n838);
    nor g2024(n3025 ,n875 ,n838);
    nor g2025(n3024 ,n898 ,n2124);
    nor g2026(n3023 ,n879 ,n838);
    nor g2027(n3022 ,n895 ,n838);
    nor g2028(n3021 ,n931 ,n2124);
    nor g2029(n3020 ,n907 ,n2124);
    nor g2030(n3019 ,n881 ,n838);
    nor g2031(n3018 ,n883 ,n838);
    nor g2032(n3017 ,n927 ,n838);
    nor g2033(n3016 ,n911 ,n835);
    nor g2034(n3015 ,n885 ,n835);
    nor g2035(n3014 ,n914 ,n835);
    nor g2036(n3013 ,n933 ,n835);
    nor g2037(n3012 ,n891 ,n2123);
    nor g2038(n3011 ,n930 ,n835);
    nor g2039(n3010 ,n906 ,n835);
    nor g2040(n3009 ,n878 ,n2123);
    nor g2041(n3008 ,n873 ,n835);
    nor g2042(n3007 ,n912 ,n835);
    nor g2043(n3006 ,n922 ,n835);
    nor g2044(n3005 ,n889 ,n835);
    nor g2045(n3004 ,n932 ,n835);
    nor g2046(n3003 ,n893 ,n2123);
    nor g2047(n3002 ,n905 ,n835);
    nor g2048(n3001 ,n876 ,n835);
    nor g2049(n3000 ,n915 ,n835);
    nor g2050(n2999 ,n919 ,n835);
    nor g2051(n2998 ,n904 ,n835);
    nor g2052(n2997 ,n896 ,n835);
    nor g2053(n2996 ,n923 ,n835);
    nor g2054(n2995 ,n910 ,n835);
    nor g2055(n2994 ,n875 ,n835);
    nor g2056(n2993 ,n898 ,n835);
    nor g2057(n2992 ,n879 ,n2123);
    nor g2058(n2991 ,n895 ,n835);
    nor g2059(n2990 ,n881 ,n2122);
    nor g2060(n2989 ,n931 ,n835);
    nor g2061(n2988 ,n907 ,n2123);
    nor g2062(n2987 ,n881 ,n2123);
    nor g2063(n2986 ,n883 ,n835);
    nor g2064(n2985 ,n927 ,n835);
    nor g2065(n2984 ,n891 ,n832);
    nor g2066(n2983 ,n885 ,n832);
    nor g2067(n2982 ,n911 ,n832);
    nor g2068(n2981 ,n933 ,n832);
    nor g2069(n2980 ,n906 ,n832);
    nor g2070(n2979 ,n930 ,n2122);
    nor g2071(n2978 ,n873 ,n832);
    nor g2072(n2977 ,n912 ,n832);
    nor g2073(n2976 ,n922 ,n832);
    nor g2074(n2975 ,n889 ,n832);
    nor g2075(n2974 ,n893 ,n832);
    nor g2076(n2973 ,n932 ,n832);
    nor g2077(n2972 ,n905 ,n832);
    nor g2078(n2971 ,n876 ,n832);
    nor g2079(n2970 ,n915 ,n832);
    nor g2080(n2969 ,n904 ,n832);
    nor g2081(n2968 ,n923 ,n2122);
    nor g2082(n2967 ,n910 ,n832);
    nor g2083(n2966 ,n877 ,n835);
    nor g2084(n2965 ,n919 ,n832);
    nor g2085(n2964 ,n898 ,n2122);
    nor g2086(n2963 ,n879 ,n2122);
    nor g2087(n2962 ,n895 ,n832);
    nor g2088(n2961 ,n907 ,n832);
    nor g2089(n2960 ,n883 ,n832);
    nor g2090(n2959 ,n1241 ,n827);
    nor g2091(n2958 ,n897 ,n827);
    nor g2092(n2957 ,n903 ,n827);
    nor g2093(n2956 ,n966 ,n830);
    nor g2094(n2955 ,n1333 ,n827);
    nor g2095(n2954 ,n1229 ,n827);
    nor g2096(n2953 ,n1248 ,n827);
    nor g2097(n2952 ,n1257 ,n827);
    nor g2098(n2951 ,n1247 ,n827);
    nor g2099(n2950 ,n946 ,n827);
    nor g2100(n2949 ,n1255 ,n827);
    nor g2101(n2948 ,n892 ,n827);
    nor g2102(n2947 ,n1224 ,n828);
    nor g2103(n2946 ,n1233 ,n828);
    nor g2104(n2945 ,n963 ,n828);
    nor g2105(n2944 ,n1223 ,n827);
    nor g2106(n2943 ,n1261 ,n827);
    nor g2107(n2942 ,n1329 ,n828);
    nor g2108(n2941 ,n926 ,n828);
    nor g2109(n2940 ,n1288 ,n828);
    nor g2110(n2939 ,n1394 ,n828);
    nor g2111(n2938 ,n1293 ,n827);
    nor g2112(n2937 ,n1368 ,n827);
    nor g2113(n2936 ,n1279 ,n827);
    nor g2114(n2935 ,n1264 ,n827);
    nor g2115(n2934 ,n1252 ,n827);
    nor g2116(n2933 ,n1235 ,n828);
    nor g2117(n2932 ,n1275 ,n828);
    nor g2118(n2931 ,n1314 ,n827);
    nor g2119(n2930 ,n1273 ,n827);
    nor g2120(n2929 ,n1325 ,n828);
    nor g2121(n2928 ,n1262 ,n827);
    nor g2122(n2927 ,n902 ,n827);
    nor g2123(n2926 ,n1372 ,n828);
    nor g2124(n2925 ,n908 ,n828);
    nor g2125(n2924 ,n1360 ,n827);
    nor g2126(n2923 ,n1403 ,n827);
    nor g2127(n2922 ,n1358 ,n827);
    nor g2128(n2921 ,n948 ,n828);
    nor g2129(n2920 ,n1408 ,n828);
    nor g2130(n2919 ,n958 ,n836);
    nor g2131(n2918 ,n957 ,n828);
    nor g2132(n2917 ,n1392 ,n836);
    nor g2133(n2916 ,n1407 ,n828);
    nor g2134(n2915 ,n1251 ,n833);
    nor g2135(n2914 ,n1326 ,n836);
    nor g2136(n2913 ,n1298 ,n828);
    nor g2137(n2912 ,n1290 ,n833);
    nor g2138(n2911 ,n1320 ,n828);
    nor g2139(n2910 ,n1388 ,n836);
    or g2140(n2909 ,n1580 ,n1884);
    nor g2141(n2908 ,n944 ,n836);
    nor g2142(n2907 ,n1374 ,n827);
    nor g2143(n2906 ,n1312 ,n830);
    nor g2144(n2905 ,n1328 ,n828);
    nor g2145(n2904 ,n939 ,n828);
    nor g2146(n2903 ,n937 ,n836);
    nor g2147(n2902 ,n1272 ,n833);
    nor g2148(n2901 ,n1337 ,n828);
    nor g2149(n2900 ,n1373 ,n828);
    nor g2150(n2899 ,n1232 ,n830);
    nor g2151(n2898 ,n1383 ,n836);
    nor g2152(n2897 ,n1319 ,n830);
    nor g2153(n2896 ,n1404 ,n828);
    nor g2154(n2895 ,n1375 ,n830);
    nor g2155(n2894 ,n1364 ,n828);
    nor g2156(n2893 ,n1352 ,n830);
    nor g2157(n2892 ,n1289 ,n830);
    nor g2158(n2891 ,n1371 ,n827);
    nor g2159(n2890 ,n1390 ,n836);
    nor g2160(n2889 ,n1402 ,n828);
    nor g2161(n2888 ,n1355 ,n836);
    nor g2162(n2887 ,n1399 ,n827);
    nor g2163(n2886 ,n1323 ,n827);
    nor g2164(n2885 ,n1384 ,n836);
    nor g2165(n2884 ,n942 ,n827);
    nor g2166(n2883 ,n1387 ,n836);
    nor g2167(n2882 ,n1397 ,n827);
    nor g2168(n2881 ,n909 ,n830);
    nor g2169(n2880 ,n960 ,n830);
    nor g2170(n2879 ,n1353 ,n836);
    nor g2171(n2878 ,n1291 ,n837);
    nor g2172(n2877 ,n950 ,n837);
    nor g2173(n2876 ,n1357 ,n837);
    nor g2174(n2875 ,n964 ,n830);
    nor g2175(n2874 ,n1260 ,n833);
    nor g2176(n2873 ,n1307 ,n836);
    nor g2177(n2872 ,n961 ,n836);
    nor g2178(n2871 ,n941 ,n837);
    nor g2179(n2870 ,n1338 ,n837);
    nor g2180(n2869 ,n1351 ,n837);
    nor g2181(n2868 ,n1303 ,n837);
    nor g2182(n2867 ,n1342 ,n836);
    nor g2183(n2866 ,n1359 ,n836);
    nor g2184(n2865 ,n1311 ,n836);
    nor g2185(n2864 ,n1330 ,n836);
    nor g2186(n2863 ,n965 ,n836);
    nor g2187(n2862 ,n1313 ,n837);
    nor g2188(n2861 ,n1409 ,n837);
    nor g2189(n2860 ,n1322 ,n836);
    nor g2190(n2859 ,n1332 ,n836);
    nor g2191(n2858 ,n936 ,n837);
    nor g2192(n2857 ,n1369 ,n836);
    nor g2193(n2856 ,n1327 ,n836);
    nor g2194(n2855 ,n1324 ,n833);
    nor g2195(n2854 ,n955 ,n833);
    nor g2196(n2853 ,n947 ,n833);
    nor g2197(n2852 ,n1391 ,n833);
    nor g2198(n2851 ,n1318 ,n833);
    nor g2199(n2850 ,n1363 ,n833);
    nor g2200(n2849 ,n1379 ,n833);
    nor g2201(n2848 ,n1362 ,n833);
    nor g2202(n2847 ,n1381 ,n834);
    nor g2203(n2846 ,n1395 ,n834);
    nor g2204(n2845 ,n1300 ,n834);
    nor g2205(n2844 ,n1356 ,n833);
    nor g2206(n2843 ,n959 ,n833);
    nor g2207(n2842 ,n1331 ,n834);
    nor g2208(n2841 ,n1361 ,n834);
    nor g2209(n2840 ,n1349 ,n834);
    nor g2210(n2839 ,n1398 ,n834);
    nor g2211(n2838 ,n1376 ,n833);
    nor g2212(n2837 ,n945 ,n833);
    nor g2213(n2836 ,n1310 ,n833);
    nor g2214(n2835 ,n894 ,n830);
    nor g2215(n2834 ,n1256 ,n833);
    nor g2216(n2833 ,n1321 ,n833);
    nor g2217(n2832 ,n1317 ,n834);
    nor g2218(n2831 ,n1344 ,n834);
    nor g2219(n2830 ,n1239 ,n830);
    nor g2220(n2829 ,n1302 ,n833);
    nor g2221(n2828 ,n1382 ,n831);
    nor g2222(n2827 ,n1367 ,n833);
    nor g2223(n2826 ,n1271 ,n831);
    nor g2224(n2825 ,n1244 ,n837);
    nor g2225(n2824 ,n956 ,n834);
    nor g2226(n2823 ,n940 ,n833);
    nor g2227(n2822 ,n1336 ,n833);
    nor g2228(n2821 ,n1400 ,n834);
    nor g2229(n2820 ,n1405 ,n834);
    nor g2230(n2819 ,n882 ,n831);
    nor g2231(n2818 ,n1345 ,n833);
    nor g2232(n2817 ,n938 ,n830);
    nor g2233(n2816 ,n1305 ,n833);
    nor g2234(n2815 ,n1240 ,n837);
    nor g2235(n2814 ,n1366 ,n830);
    nor g2236(n2813 ,n1292 ,n836);
    nor g2237(n2812 ,n1226 ,n836);
    nor g2238(n2811 ,n1276 ,n836);
    nor g2239(n2810 ,n916 ,n837);
    nor g2240(n2809 ,n1245 ,n833);
    nor g2241(n2808 ,n1393 ,n831);
    nor g2242(n2807 ,n1234 ,n837);
    nor g2243(n2806 ,n1340 ,n831);
    nor g2244(n2805 ,n1269 ,n837);
    nor g2245(n2804 ,n1284 ,n837);
    nor g2246(n2803 ,n935 ,n837);
    nor g2247(n2802 ,n1354 ,n831);
    nor g2248(n2801 ,n1246 ,n837);
    nor g2249(n2800 ,n924 ,n836);
    nor g2250(n2799 ,n884 ,n837);
    nor g2251(n2798 ,n1265 ,n837);
    nor g2252(n2797 ,n901 ,n837);
    nor g2253(n2796 ,n1389 ,n831);
    nor g2254(n2795 ,n1227 ,n837);
    nor g2255(n2794 ,n928 ,n837);
    nor g2256(n2793 ,n1315 ,n830);
    nor g2257(n2792 ,n1231 ,n837);
    nor g2258(n2791 ,n1278 ,n836);
    nor g2259(n2790 ,n1268 ,n837);
    nor g2260(n2789 ,n1285 ,n830);
    nor g2261(n2788 ,n1370 ,n830);
    nor g2262(n2787 ,n890 ,n836);
    nor g2263(n2786 ,n929 ,n830);
    nor g2264(n2785 ,n1286 ,n836);
    nor g2265(n2784 ,n1243 ,n836);
    nor g2266(n2783 ,n917 ,n836);
    nor g2267(n2782 ,n1350 ,n830);
    nor g2268(n2781 ,n1253 ,n837);
    nor g2269(n2780 ,n1295 ,n834);
    nor g2270(n2779 ,n1346 ,n831);
    nor g2271(n2778 ,n921 ,n834);
    nor g2272(n2777 ,n1282 ,n834);
    nor g2273(n2776 ,n1308 ,n831);
    nor g2274(n2775 ,n1334 ,n830);
    nor g2275(n2774 ,n1236 ,n834);
    nor g2276(n2773 ,n1294 ,n830);
    nor g2277(n2772 ,n880 ,n834);
    nor g2278(n2771 ,n1309 ,n831);
    nor g2279(n2770 ,n1280 ,n834);
    nor g2280(n2769 ,n1250 ,n833);
    nor g2281(n2768 ,n1316 ,n830);
    nor g2282(n2767 ,n886 ,n834);
    nor g2283(n2766 ,n900 ,n834);
    nor g2284(n2765 ,n925 ,n830);
    nor g2285(n2764 ,n1281 ,n834);
    nor g2286(n2763 ,n962 ,n831);
    nor g2287(n2762 ,n913 ,n834);
    nor g2288(n2761 ,n1249 ,n834);
    nor g2289(n2760 ,n1266 ,n834);
    nor g2290(n2759 ,n1225 ,n833);
    nor g2291(n2758 ,n1242 ,n834);
    nor g2292(n2757 ,n1237 ,n833);
    nor g2293(n2756 ,n1378 ,n831);
    nor g2294(n2755 ,n1230 ,n833);
    nor g2295(n2754 ,n952 ,n830);
    nor g2296(n2753 ,n1263 ,n833);
    nor g2297(n2752 ,n1406 ,n830);
    nor g2298(n2751 ,n918 ,n833);
    nor g2299(n2750 ,n1274 ,n830);
    nor g2300(n2749 ,n1339 ,n831);
    nor g2301(n2748 ,n1254 ,n831);
    nor g2302(n2747 ,n887 ,n831);
    nor g2303(n2746 ,n954 ,n831);
    nor g2304(n2745 ,n920 ,n831);
    nor g2305(n2744 ,n1267 ,n831);
    nor g2306(n2743 ,n1347 ,n830);
    nor g2307(n2742 ,n899 ,n834);
    nor g2308(n2741 ,n1297 ,n831);
    nor g2309(n2740 ,n1287 ,n831);
    nor g2310(n2739 ,n1386 ,n831);
    nor g2311(n2738 ,n1283 ,n831);
    nor g2312(n2737 ,n1238 ,n831);
    nor g2313(n2736 ,n934 ,n831);
    nor g2314(n2735 ,n1277 ,n830);
    nor g2315(n2734 ,n1228 ,n831);
    nor g2316(n2733 ,n1296 ,n830);
    nor g2317(n2732 ,n1365 ,n830);
    nor g2318(n2731 ,n874 ,n830);
    xnor g2319(n2729 ,n1862 ,n23[0]);
    nor g2320(n2728 ,n1258 ,n830);
    nor g2321(n2727 ,n1270 ,n828);
    or g2322(n2726 ,n1821 ,n1885);
    or g2323(n2725 ,n1814 ,n1882);
    or g2324(n2724 ,n1806 ,n1881);
    nor g2325(n2723 ,n1306 ,n831);
    nor g2326(n2722 ,n861 ,n829);
    nor g2327(n2721 ,n847 ,n2121);
    nor g2328(n2720 ,n862 ,n829);
    nor g2329(n2719 ,n854 ,n829);
    nor g2330(n2718 ,n851 ,n2121);
    nor g2331(n2717 ,n846 ,n829);
    nor g2332(n2716 ,n849 ,n829);
    nor g2333(n2715 ,n859 ,n829);
    nor g2334(n2714 ,n860 ,n829);
    nor g2335(n2713 ,n853 ,n2121);
    nor g2336(n2712 ,n867 ,n829);
    nor g2337(n2711 ,n845 ,n829);
    nor g2338(n2710 ,n863 ,n829);
    nor g2339(n2709 ,n858 ,n829);
    nor g2340(n2708 ,n848 ,n829);
    nor g2341(n2707 ,n850 ,n829);
    nor g2342(n2706 ,n865 ,n829);
    nor g2343(n2705 ,n852 ,n832);
    nor g2344(n2704 ,n855 ,n2121);
    nor g2345(n2703 ,n864 ,n829);
    nor g2346(n2702 ,n869 ,n829);
    nor g2347(n2701 ,n868 ,n829);
    nor g2348(n2700 ,n852 ,n829);
    nor g2349(n2699 ,n866 ,n829);
    nor g2350(n2698 ,n857 ,n829);
    nor g2351(n2697 ,n870 ,n829);
    nor g2352(n2696 ,n856 ,n829);
    nor g2353(n2695 ,n853 ,n2122);
    nor g2354(n2694 ,n868 ,n832);
    nor g2355(n2693 ,n849 ,n838);
    nor g2356(n2692 ,n850 ,n832);
    nor g2357(n2691 ,n865 ,n2122);
    nor g2358(n2690 ,n851 ,n835);
    nor g2359(n2689 ,n862 ,n2123);
    nor g2360(n2688 ,n864 ,n832);
    nor g2361(n2687 ,n856 ,n2124);
    nor g2362(n2686 ,n870 ,n838);
    nor g2363(n2685 ,n857 ,n835);
    nor g2364(n2684 ,n848 ,n835);
    nor g2365(n2683 ,n848 ,n832);
    nor g2366(n2682 ,n862 ,n832);
    nor g2367(n2681 ,n868 ,n838);
    nor g2368(n2680 ,n869 ,n2124);
    nor g2369(n2679 ,n845 ,n2123);
    nor g2370(n2678 ,n869 ,n832);
    nor g2371(n2677 ,n845 ,n2122);
    nor g2372(n2676 ,n850 ,n838);
    nor g2373(n2675 ,n857 ,n832);
    nor g2374(n2674 ,n848 ,n838);
    nor g2375(n2673 ,n861 ,n838);
    nor g2376(n2672 ,n847 ,n838);
    nor g2377(n2671 ,n862 ,n2124);
    nor g2378(n2670 ,n854 ,n838);
    nor g2379(n2669 ,n851 ,n838);
    nor g2380(n2668 ,n846 ,n838);
    nor g2381(n2667 ,n859 ,n838);
    nor g2382(n2666 ,n860 ,n838);
    nor g2383(n2665 ,n853 ,n838);
    nor g2384(n2664 ,n867 ,n838);
    nor g2385(n2663 ,n845 ,n2124);
    nor g2386(n2662 ,n863 ,n838);
    nor g2387(n2661 ,n858 ,n838);
    nor g2388(n2660 ,n865 ,n838);
    nor g2389(n2659 ,n855 ,n838);
    nor g2390(n2658 ,n864 ,n838);
    nor g2391(n2657 ,n852 ,n838);
    nor g2392(n2656 ,n866 ,n838);
    nor g2393(n2655 ,n857 ,n838);
    nor g2394(n2654 ,n861 ,n835);
    nor g2395(n2653 ,n847 ,n835);
    nor g2396(n2652 ,n854 ,n835);
    nor g2397(n2651 ,n846 ,n835);
    nor g2398(n2650 ,n849 ,n2123);
    nor g2399(n2649 ,n859 ,n835);
    nor g2400(n2648 ,n860 ,n835);
    nor g2401(n2647 ,n853 ,n835);
    nor g2402(n2646 ,n867 ,n835);
    nor g2403(n2645 ,n863 ,n835);
    nor g2404(n2644 ,n867 ,n832);
    nor g2405(n2643 ,n858 ,n835);
    nor g2406(n2642 ,n850 ,n835);
    nor g2407(n2641 ,n865 ,n2123);
    nor g2408(n2640 ,n855 ,n835);
    nor g2409(n2639 ,n864 ,n835);
    nor g2410(n2638 ,n869 ,n835);
    nor g2411(n2637 ,n868 ,n835);
    nor g2412(n2636 ,n852 ,n835);
    nor g2413(n2635 ,n866 ,n835);
    nor g2414(n2634 ,n870 ,n835);
    nor g2415(n2633 ,n856 ,n835);
    nor g2416(n2632 ,n861 ,n832);
    nor g2417(n2631 ,n847 ,n832);
    nor g2418(n2630 ,n854 ,n832);
    nor g2419(n2629 ,n851 ,n832);
    nor g2420(n2628 ,n846 ,n832);
    nor g2421(n2627 ,n849 ,n2122);
    nor g2422(n2626 ,n859 ,n832);
    nor g2423(n2625 ,n860 ,n832);
    nor g2424(n2624 ,n863 ,n832);
    nor g2425(n2623 ,n858 ,n832);
    nor g2426(n2622 ,n855 ,n832);
    nor g2427(n2621 ,n866 ,n832);
    nor g2428(n2620 ,n870 ,n832);
    nor g2429(n2619 ,n856 ,n832);
    nor g2430(n2618 ,n839 ,n1876);
    nor g2431(n2617 ,n841 ,n1877);
    nor g2432(n2616 ,n811 ,n1878);
    nor g2433(n2615 ,n813 ,n1879);
    or g2434(n2614 ,n2356 ,n2347);
    or g2435(n2613 ,n2364 ,n2238);
    or g2436(n2612 ,n2355 ,n2360);
    or g2437(n2611 ,n2351 ,n2298);
    or g2438(n2610 ,n2341 ,n2338);
    or g2439(n2609 ,n2361 ,n2350);
    or g2440(n2608 ,n2343 ,n2345);
    or g2441(n2607 ,n2342 ,n2363);
    or g2442(n2606 ,n2332 ,n2177);
    or g2443(n2605 ,n2331 ,n2333);
    or g2444(n2604 ,n2318 ,n2310);
    or g2445(n2603 ,n2367 ,n2339);
    or g2446(n2602 ,n2319 ,n2321);
    or g2447(n2601 ,n2290 ,n2280);
    or g2448(n2600 ,n2311 ,n2358);
    or g2449(n2599 ,n2221 ,n2220);
    or g2450(n2598 ,n2317 ,n2314);
    or g2451(n2597 ,n2309 ,n2359);
    or g2452(n2596 ,n2326 ,n2313);
    or g2453(n2595 ,n2340 ,n2362);
    or g2454(n2594 ,n2330 ,n2336);
    or g2455(n2593 ,n2300 ,n2302);
    or g2456(n2592 ,n2304 ,n2299);
    or g2457(n2591 ,n2297 ,n2301);
    or g2458(n2590 ,n2183 ,n2293);
    or g2459(n2589 ,n2184 ,n2306);
    or g2460(n2588 ,n2273 ,n2289);
    or g2461(n2587 ,n2279 ,n2288);
    or g2462(n2586 ,n2284 ,n2287);
    or g2463(n2585 ,n2277 ,n2283);
    or g2464(n2584 ,n2186 ,n2278);
    or g2465(n2583 ,n2202 ,n2168);
    nor g2466(n2582 ,n2004 ,n2138);
    nor g2467(n2581 ,n2002 ,n2137);
    nor g2468(n2580 ,n2001 ,n2136);
    nor g2469(n2579 ,n1912 ,n2084);
    nor g2470(n2578 ,n2000 ,n2134);
    nor g2471(n2577 ,n1999 ,n2133);
    nor g2472(n2576 ,n1998 ,n2132);
    nor g2473(n2575 ,n1997 ,n2131);
    nor g2474(n2574 ,n2120 ,n2130);
    nor g2475(n2573 ,n1994 ,n2129);
    nor g2476(n2572 ,n1993 ,n2128);
    nor g2477(n2571 ,n1992 ,n2126);
    nor g2478(n2570 ,n1943 ,n2070);
    nor g2479(n2569 ,n1991 ,n2371);
    nor g2480(n2568 ,n1990 ,n1996);
    nor g2481(n2567 ,n1931 ,n2119);
    nor g2482(n2566 ,n1989 ,n2118);
    nor g2483(n2565 ,n1987 ,n2117);
    nor g2484(n2564 ,n1986 ,n2116);
    nor g2485(n2563 ,n1927 ,n2110);
    nor g2486(n2562 ,n1985 ,n2115);
    nor g2487(n2561 ,n1984 ,n2114);
    nor g2488(n2560 ,n1982 ,n2113);
    nor g2489(n2559 ,n2006 ,n2020);
    nor g2490(n2558 ,n1981 ,n2112);
    nor g2491(n2557 ,n1892 ,n2111);
    nor g2492(n2556 ,n1980 ,n2109);
    nor g2493(n2555 ,n1977 ,n2108);
    nor g2494(n2554 ,n1976 ,n2107);
    nor g2495(n2553 ,n2007 ,n2105);
    nor g2496(n2552 ,n2008 ,n2104);
    nor g2497(n2551 ,n1972 ,n2103);
    nor g2498(n2550 ,n1971 ,n2102);
    nor g2499(n2549 ,n2009 ,n2101);
    nor g2500(n2548 ,n1970 ,n2100);
    nor g2501(n2547 ,n1969 ,n2099);
    nor g2502(n2546 ,n2010 ,n2098);
    nor g2503(n2545 ,n1968 ,n2097);
    nor g2504(n2544 ,n1966 ,n2096);
    nor g2505(n2543 ,n1964 ,n2095);
    nor g2506(n2542 ,n1913 ,n2094);
    nor g2507(n2541 ,n1963 ,n2093);
    nor g2508(n2540 ,n1962 ,n2092);
    nor g2509(n2539 ,n1960 ,n2091);
    nor g2510(n2538 ,n1926 ,n2090);
    nor g2511(n2537 ,n1958 ,n2089);
    nor g2512(n2536 ,n1956 ,n2088);
    nor g2513(n2535 ,n1955 ,n2087);
    nor g2514(n2534 ,n1936 ,n2086);
    nor g2515(n2533 ,n1961 ,n2045);
    nor g2516(n2532 ,n1954 ,n2085);
    nor g2517(n2531 ,n1953 ,n2082);
    nor g2518(n2530 ,n1952 ,n2081);
    nor g2519(n2529 ,n1951 ,n2080);
    nor g2520(n2528 ,n1950 ,n2079);
    nor g2521(n2527 ,n1948 ,n2078);
    nor g2522(n2526 ,n1947 ,n2077);
    nor g2523(n2525 ,n1959 ,n2076);
    nor g2524(n2524 ,n1967 ,n2075);
    nor g2525(n2523 ,n1973 ,n2074);
    nor g2526(n2522 ,n1945 ,n2073);
    nor g2527(n2521 ,n1979 ,n2072);
    nor g2528(n2520 ,n1944 ,n2071);
    nor g2529(n2519 ,n1942 ,n2139);
    nor g2530(n2518 ,n1901 ,n2069);
    nor g2531(n2517 ,n1941 ,n2068);
    nor g2532(n2516 ,n1940 ,n2067);
    nor g2533(n2515 ,n2003 ,n2066);
    nor g2534(n2514 ,n1908 ,n2065);
    nor g2535(n2513 ,n2011 ,n2064);
    nor g2536(n2512 ,n1924 ,n2063);
    nor g2537(n2511 ,n1889 ,n2062);
    nor g2538(n2510 ,n1910 ,n2061);
    nor g2539(n2509 ,n1911 ,n2060);
    nor g2540(n2508 ,n1937 ,n2059);
    nor g2541(n2507 ,n1920 ,n2058);
    nor g2542(n2506 ,n1917 ,n2057);
    nor g2543(n2505 ,n1935 ,n2056);
    nor g2544(n2504 ,n1978 ,n2055);
    nor g2545(n2503 ,n1928 ,n2054);
    nor g2546(n2502 ,n1929 ,n2053);
    nor g2547(n2501 ,n1933 ,n2051);
    nor g2548(n2500 ,n1934 ,n2052);
    nor g2549(n2499 ,n1938 ,n2050);
    nor g2550(n2498 ,n1939 ,n2049);
    nor g2551(n2497 ,n1907 ,n2047);
    nor g2552(n2496 ,n1946 ,n2046);
    nor g2553(n2495 ,n1957 ,n2083);
    nor g2554(n2494 ,n1930 ,n2106);
    nor g2555(n2493 ,n1965 ,n2044);
    nor g2556(n2492 ,n1974 ,n2043);
    nor g2557(n2491 ,n1983 ,n2127);
    nor g2558(n2490 ,n1988 ,n2042);
    nor g2559(n2489 ,n1995 ,n2041);
    nor g2560(n2488 ,n1888 ,n2012);
    nor g2561(n2487 ,n1890 ,n2040);
    nor g2562(n2486 ,n1891 ,n2039);
    nor g2563(n2485 ,n1923 ,n2037);
    nor g2564(n2484 ,n1894 ,n2036);
    nor g2565(n2483 ,n1895 ,n2035);
    nor g2566(n2482 ,n1922 ,n2034);
    nor g2567(n2481 ,n1921 ,n2033);
    nor g2568(n2480 ,n1898 ,n2032);
    nor g2569(n2479 ,n1897 ,n2013);
    nor g2570(n2478 ,n1919 ,n2015);
    nor g2571(n2477 ,n1918 ,n2014);
    nor g2572(n2476 ,n1899 ,n2030);
    nor g2573(n2475 ,n1900 ,n2029);
    nor g2574(n2474 ,n1905 ,n2016);
    nor g2575(n2473 ,n1902 ,n2028);
    nor g2576(n2472 ,n1903 ,n2027);
    nor g2577(n2471 ,n1915 ,n2017);
    nor g2578(n2470 ,n1904 ,n2026);
    nor g2579(n2469 ,n1906 ,n2025);
    nor g2580(n2468 ,n1896 ,n2018);
    nor g2581(n2467 ,n1914 ,n2023);
    nor g2582(n2466 ,n1925 ,n2022);
    nor g2583(n2465 ,n1949 ,n2021);
    nor g2584(n2464 ,n1975 ,n2135);
    nor g2585(n2463 ,n2005 ,n2019);
    or g2586(n2462 ,n2169 ,n2195);
    or g2587(n2461 ,n2259 ,n2348);
    or g2588(n2460 ,n2247 ,n2270);
    or g2589(n2459 ,n2366 ,n2324);
    or g2590(n2458 ,n2257 ,n2256);
    or g2591(n2457 ,n2255 ,n2254);
    or g2592(n2456 ,n2222 ,n2153);
    or g2593(n2455 ,n2244 ,n2272);
    or g2594(n2454 ,n2251 ,n2370);
    or g2595(n2453 ,n2249 ,n2248);
    or g2596(n2452 ,n2245 ,n2246);
    or g2597(n2451 ,n2325 ,n2234);
    or g2598(n2450 ,n2243 ,n2125);
    or g2599(n2449 ,n2242 ,n2241);
    nor g2600(n2448 ,n1932 ,n2048);
    nor g2601(n2447 ,n1909 ,n2024);
    or g2602(n2446 ,n2239 ,n2240);
    or g2603(n2445 ,n2269 ,n2172);
    or g2604(n2444 ,n2252 ,n2334);
    or g2605(n2443 ,n2237 ,n2236);
    or g2606(n2442 ,n2235 ,n2144);
    or g2607(n2441 ,n2215 ,n2207);
    or g2608(n2440 ,n2233 ,n2232);
    or g2609(n2439 ,n2268 ,n2231);
    or g2610(n2438 ,n2187 ,n2337);
    or g2611(n2437 ,n2229 ,n2142);
    or g2612(n2436 ,n2228 ,n2145);
    or g2613(n2435 ,n2198 ,n2260);
    or g2614(n2434 ,n2224 ,n2262);
    or g2615(n2433 ,n2227 ,n2271);
    or g2616(n2432 ,n2267 ,n2225);
    or g2617(n2431 ,n2223 ,n2276);
    or g2618(n2430 ,n2292 ,n2307);
    or g2619(n2429 ,n2357 ,n2368);
    or g2620(n2428 ,n2250 ,n2261);
    or g2621(n2427 ,n2365 ,n2219);
    or g2622(n2426 ,n2217 ,n2143);
    or g2623(n2425 ,n2216 ,n2157);
    or g2624(n2424 ,n2263 ,n2226);
    or g2625(n2423 ,n2166 ,n2212);
    or g2626(n2422 ,n2323 ,n2218);
    or g2627(n2421 ,n2210 ,n2176);
    or g2628(n2420 ,n2209 ,n2208);
    or g2629(n2419 ,n2205 ,n2206);
    or g2630(n2418 ,n2152 ,n2204);
    or g2631(n2417 ,n2158 ,n2201);
    or g2632(n2416 ,n2200 ,n2182);
    or g2633(n2415 ,n2203 ,n2199);
    or g2634(n2414 ,n2167 ,n2189);
    or g2635(n2413 ,n2141 ,n2196);
    or g2636(n2412 ,n2181 ,n2173);
    or g2637(n2411 ,n2190 ,n2197);
    or g2638(n2410 ,n2175 ,n2266);
    nor g2639(n2409 ,n1916 ,n2031);
    or g2640(n2408 ,n2188 ,n2230);
    or g2641(n2407 ,n2148 ,n2147);
    or g2642(n2406 ,n2282 ,n2281);
    or g2643(n2405 ,n2178 ,n2174);
    or g2644(n2404 ,n2308 ,n2312);
    or g2645(n2403 ,n2315 ,n2179);
    or g2646(n2402 ,n2329 ,n2327);
    or g2647(n2401 ,n2349 ,n2369);
    or g2648(n2400 ,n2354 ,n2352);
    or g2649(n2399 ,n2253 ,n2258);
    or g2650(n2398 ,n2191 ,n2180);
    or g2651(n2397 ,n2291 ,n2285);
    or g2652(n2396 ,n2156 ,n2155);
    or g2653(n2395 ,n2294 ,n2295);
    or g2654(n2394 ,n2154 ,n2171);
    or g2655(n2393 ,n2335 ,n2328);
    or g2656(n2392 ,n2346 ,n2353);
    or g2657(n2391 ,n2149 ,n2140);
    or g2658(n2390 ,n2322 ,n2170);
    or g2659(n2389 ,n2192 ,n2159);
    or g2660(n2388 ,n2275 ,n2163);
    or g2661(n2387 ,n2160 ,n2286);
    or g2662(n2386 ,n2274 ,n2265);
    or g2663(n2385 ,n2213 ,n2214);
    or g2664(n2384 ,n2164 ,n2161);
    or g2665(n2383 ,n2303 ,n2316);
    or g2666(n2382 ,n2344 ,n2185);
    or g2667(n2381 ,n2264 ,n2162);
    or g2668(n2380 ,n2211 ,n2150);
    nor g2669(n2379 ,n1893 ,n2038);
    or g2670(n2378 ,n2305 ,n2320);
    or g2671(n2377 ,n2151 ,n2165);
    or g2672(n2376 ,n2296 ,n2193);
    or g2673(n2375 ,n2194 ,n2146);
    xnor g2674(n2374 ,n1872 ,n21[0]);
    xnor g2675(n2373 ,n1861 ,n22[0]);
    xnor g2676(n2372 ,n1873 ,n24[0]);
    nor g2677(n2730 ,n1739 ,n1880);
    nor g2678(n2371 ,n1050 ,n821);
    nor g2679(n2370 ,n1241 ,n818);
    nor g2680(n2369 ,n1402 ,n818);
    nor g2681(n2368 ,n1300 ,n820);
    nor g2682(n2367 ,n1309 ,n826);
    nor g2683(n2366 ,n1353 ,n824);
    nor g2684(n2365 ,n1246 ,n824);
    nor g2685(n2364 ,n960 ,n826);
    nor g2686(n2363 ,n1404 ,n817);
    nor g2687(n2362 ,n1371 ,n818);
    nor g2688(n2361 ,n1375 ,n825);
    nor g2689(n2360 ,n1362 ,n820);
    nor g2690(n2359 ,n1302 ,n819);
    nor g2691(n2358 ,n1305 ,n820);
    nor g2692(n2357 ,n1387 ,n823);
    nor g2693(n2356 ,n1383 ,n824);
    nor g2694(n2355 ,n1390 ,n824);
    nor g2695(n2354 ,n1370 ,n826);
    nor g2696(n2353 ,n1398 ,n820);
    nor g2697(n2352 ,n1325 ,n818);
    nor g2698(n2351 ,n965 ,n823);
    nor g2699(n2350 ,n1298 ,n817);
    nor g2700(n2349 ,n1352 ,n826);
    nor g2701(n2348 ,n1336 ,n819);
    nor g2702(n2347 ,n1379 ,n820);
    nor g2703(n2346 ,n941 ,n824);
    nor g2704(n2345 ,n1314 ,n818);
    nor g2705(n2344 ,n1313 ,n823);
    nor g2706(n2343 ,n1315 ,n825);
    nor g2707(n2342 ,n1350 ,n826);
    nor g2708(n2341 ,n937 ,n824);
    nor g2709(n2340 ,n1365 ,n825);
    nor g2710(n2339 ,n1394 ,n817);
    nor g2711(n2338 ,n1363 ,n819);
    nor g2712(n2337 ,n902 ,n818);
    nor g2713(n2336 ,n1310 ,n820);
    nor g2714(n2335 ,n962 ,n826);
    nor g2715(n2334 ,n1358 ,n817);
    nor g2716(n2333 ,n1349 ,n819);
    nor g2717(n2332 ,n1389 ,n825);
    nor g2718(n2331 ,n961 ,n823);
    nor g2719(n2330 ,n1303 ,n823);
    nor g2720(n2329 ,n944 ,n823);
    nor g2721(n2328 ,n1407 ,n817);
    nor g2722(n2327 ,n1318 ,n819);
    nor g2723(n2326 ,n1340 ,n825);
    nor g2724(n2325 ,n1226 ,n823);
    nor g2725(n2324 ,n1356 ,n819);
    nor g2726(n2323 ,n954 ,n825);
    nor g2727(n2322 ,n1351 ,n823);
    nor g2728(n2321 ,n1391 ,n819);
    nor g2729(n2320 ,n1397 ,n817);
    nor g2730(n2319 ,n1388 ,n824);
    nor g2731(n2318 ,n1382 ,n825);
    nor g2732(n2317 ,n1307 ,n823);
    nor g2733(n2316 ,n1373 ,n817);
    nor g2734(n2315 ,n1354 ,n825);
    nor g2735(n2314 ,n1361 ,n819);
    nor g2736(n2313 ,n963 ,n817);
    nor g2737(n2312 ,n947 ,n820);
    nor g2738(n2311 ,n1327 ,n823);
    nor g2739(n2310 ,n957 ,n818);
    nor g2740(n2309 ,n1330 ,n823);
    nor g2741(n2308 ,n1326 ,n823);
    nor g2742(n2307 ,n1250 ,n819);
    nor g2743(n2306 ,n1333 ,n817);
    nor g2744(n2305 ,n966 ,n826);
    nor g2745(n2304 ,n1393 ,n825);
    nor g2746(n2303 ,n1386 ,n825);
    nor g2747(n2302 ,n955 ,n819);
    nor g2748(n2301 ,n959 ,n819);
    nor g2749(n2300 ,n1392 ,n823);
    nor g2750(n2299 ,n946 ,n817);
    nor g2751(n2298 ,n1367 ,n819);
    nor g2752(n2297 ,n1357 ,n823);
    nor g2753(n2296 ,n890 ,n823);
    nor g2754(n2295 ,n1408 ,n817);
    nor g2755(n2294 ,n1316 ,n825);
    nor g2756(n2293 ,n1324 ,n819);
    nor g2757(n2292 ,n935 ,n823);
    nor g2758(n2291 ,n950 ,n823);
    nor g2759(n2290 ,n1347 ,n825);
    nor g2760(n2289 ,n942 ,n817);
    nor g2761(n2288 ,n1345 ,n819);
    nor g2762(n2287 ,n1344 ,n819);
    nor g2763(n2286 ,n1385 ,n817);
    nor g2764(n2285 ,n1331 ,n819);
    nor g2765(n2284 ,n1311 ,n824);
    nor g2766(n2283 ,n948 ,n817);
    nor g2767(n2282 ,n1253 ,n824);
    nor g2768(n2281 ,n1245 ,n819);
    nor g2769(n2280 ,n1337 ,n817);
    nor g2770(n2279 ,n1369 ,n823);
    nor g2771(n2278 ,n908 ,n817);
    nor g2772(n2277 ,n1334 ,n825);
    nor g2773(n2276 ,n892 ,n817);
    nor g2774(n2275 ,n1406 ,n825);
    nor g2775(n2274 ,n1342 ,n823);
    nor g2776(n2273 ,n1306 ,n825);
    nor g2777(n2272 ,n1242 ,n820);
    nor g2778(n2271 ,n1255 ,n818);
    nor g2779(n2270 ,n918 ,n820);
    nor g2780(n2269 ,n916 ,n824);
    nor g2781(n2268 ,n1234 ,n823);
    nor g2782(n2267 ,n1284 ,n824);
    nor g2783(n2266 ,n1237 ,n819);
    nor g2784(n2265 ,n1321 ,n819);
    nor g2785(n2264 ,n1332 ,n824);
    nor g2786(n2263 ,n1319 ,n825);
    nor g2787(n2262 ,n1317 ,n820);
    nor g2788(n2261 ,n1405 ,n819);
    nor g2789(n2260 ,n1264 ,n818);
    nor g2790(n2259 ,n1322 ,n824);
    nor g2791(n2258 ,n1381 ,n820);
    nor g2792(n2257 ,n1254 ,n825);
    nor g2793(n2256 ,n1270 ,n817);
    nor g2794(n2255 ,n1240 ,n823);
    nor g2795(n2254 ,n1295 ,n820);
    nor g2796(n2253 ,n1355 ,n823);
    nor g2797(n2252 ,n1308 ,n826);
    nor g2798(n2251 ,n887 ,n826);
    nor g2799(n2250 ,n936 ,n824);
    nor g2800(n2249 ,n1292 ,n823);
    nor g2801(n2248 ,n1272 ,n820);
    nor g2802(n2247 ,n917 ,n823);
    nor g2803(n2246 ,n897 ,n817);
    nor g2804(n2245 ,n909 ,n825);
    nor g2805(n2244 ,n1278 ,n823);
    nor g2806(n2243 ,n920 ,n825);
    nor g2807(n2242 ,n1276 ,n824);
    nor g2808(n2241 ,n1282 ,n819);
    nor g2809(n2240 ,n1229 ,n818);
    nor g2810(n2239 ,n1267 ,n826);
    nor g2811(n2238 ,n1372 ,n817);
    nor g2812(n2237 ,n1274 ,n825);
    nor g2813(n2236 ,n1248 ,n818);
    nor g2814(n2235 ,n1244 ,n823);
    nor g2815(n2234 ,n921 ,n819);
    nor g2816(n2233 ,n1297 ,n826);
    nor g2817(n2232 ,n1257 ,n818);
    nor g2818(n2231 ,n880 ,n820);
    nor g2819(n2230 ,n1263 ,n819);
    nor g2820(n2229 ,n1287 ,n826);
    nor g2821(n2228 ,n1269 ,n823);
    nor g2822(n2227 ,n925 ,n826);
    nor g2823(n2226 ,n1360 ,n818);
    nor g2824(n2225 ,n1280 ,n819);
    nor g2825(n2224 ,n1359 ,n824);
    nor g2826(n2223 ,n1283 ,n825);
    nor g2827(n2222 ,n1312 ,n825);
    nor g2828(n2221 ,n1238 ,n826);
    nor g2829(n2220 ,n1224 ,n817);
    nor g2830(n2219 ,n886 ,n819);
    nor g2831(n2218 ,n939 ,n817);
    nor g2832(n2217 ,n934 ,n825);
    nor g2833(n2216 ,n924 ,n824);
    nor g2834(n2215 ,n1346 ,n825);
    nor g2835(n2214 ,n1223 ,n818);
    nor g2836(n2213 ,n1277 ,n825);
    nor g2837(n2212 ,n1281 ,n820);
    nor g2838(n2211 ,n938 ,n826);
    nor g2839(n2210 ,n1228 ,n825);
    nor g2840(n2209 ,n1265 ,n824);
    nor g2841(n2208 ,n1260 ,n819);
    nor g2842(n2207 ,n1403 ,n817);
    nor g2843(n2206 ,n926 ,n817);
    nor g2844(n2205 ,n1289 ,n825);
    nor g2845(n2204 ,n913 ,n819);
    nor g2846(n2203 ,n1231 ,n824);
    nor g2847(n2202 ,n1339 ,n826);
    nor g2848(n2201 ,n1249 ,n820);
    nor g2849(n2200 ,n1232 ,n826);
    nor g2850(n2199 ,n1225 ,n820);
    nor g2851(n2198 ,n1294 ,n826);
    nor g2852(n2197 ,n1279 ,n817);
    nor g2853(n2196 ,n1251 ,n820);
    nor g2854(n2195 ,n1395 ,n820);
    nor g2855(n2194 ,n894 ,n826);
    nor g2856(n2193 ,n1230 ,n820);
    nor g2857(n2192 ,n1271 ,n826);
    nor g2858(n2191 ,n874 ,n825);
    nor g2859(n2190 ,n1285 ,n825);
    nor g2860(n2189 ,n1262 ,n818);
    nor g2861(n2188 ,n1243 ,n824);
    nor g2862(n2187 ,n1239 ,n825);
    nor g2863(n2186 ,n1258 ,n826);
    nor g2864(n2185 ,n956 ,n819);
    nor g2865(n2184 ,n1366 ,n826);
    nor g2866(n2183 ,n958 ,n823);
    nor g2867(n2182 ,n1293 ,n817);
    nor g2868(n2181 ,n1291 ,n823);
    nor g2869(n2180 ,n1273 ,n817);
    nor g2870(n2179 ,n1329 ,n818);
    nor g2871(n2178 ,n928 ,n823);
    nor g2872(n2177 ,n1368 ,n818);
    nor g2873(n2176 ,n1261 ,n818);
    nor g2874(n2175 ,n1286 ,n824);
    nor g2875(n2174 ,n1266 ,n819);
    nor g2876(n2173 ,n899 ,n819);
    nor g2877(n2172 ,n1290 ,n820);
    nor g2878(n2171 ,n940 ,n820);
    nor g2879(n2170 ,n945 ,n820);
    nor g2880(n2169 ,n1384 ,n824);
    nor g2881(n2168 ,n1328 ,n818);
    nor g2882(n2167 ,n882 ,n826);
    nor g2883(n2166 ,n884 ,n824);
    nor g2884(n2165 ,n1376 ,n819);
    nor g2885(n2164 ,n1296 ,n825);
    nor g2886(n2163 ,n1374 ,n818);
    nor g2887(n2162 ,n1400 ,n819);
    nor g2888(n2161 ,n1288 ,n817);
    nor g2889(n2160 ,n952 ,n825);
    nor g2890(n2159 ,n1275 ,n817);
    nor g2891(n2158 ,n1227 ,n823);
    nor g2892(n2157 ,n900 ,n820);
    nor g2893(n2156 ,n964 ,n826);
    nor g2894(n2155 ,n1364 ,n817);
    nor g2895(n2154 ,n1409 ,n823);
    nor g2896(n2153 ,n1399 ,n818);
    nor g2897(n2152 ,n901 ,n824);
    nor g2898(n2151 ,n1338 ,n824);
    nor g2899(n2150 ,n1323 ,n818);
    nor g2900(n2149 ,n929 ,n826);
    nor g2901(n2148 ,n1378 ,n826);
    nor g2902(n2147 ,n1320 ,n818);
    nor g2903(n2146 ,n1235 ,n817);
    nor g2904(n2145 ,n1256 ,n820);
    nor g2905(n2144 ,n1236 ,n820);
    nor g2906(n2143 ,n1233 ,n817);
    nor g2907(n2142 ,n1247 ,n818);
    nor g2908(n2141 ,n1268 ,n824);
    nor g2909(n2140 ,n1252 ,n818);
    nor g2910(n2139 ,n1201 ,n815);
    nor g2911(n2138 ,n1139 ,n821);
    nor g2912(n2137 ,n1185 ,n821);
    nor g2913(n2136 ,n1189 ,n821);
    nor g2914(n2135 ,n1064 ,n816);
    nor g2915(n2134 ,n1134 ,n821);
    nor g2916(n2133 ,n1030 ,n821);
    nor g2917(n2132 ,n1215 ,n821);
    nor g2918(n2131 ,n1176 ,n821);
    nor g2919(n2130 ,n1137 ,n821);
    nor g2920(n2129 ,n1169 ,n821);
    nor g2921(n2128 ,n1103 ,n821);
    nor g2922(n2127 ,n1056 ,n822);
    nor g2923(n2126 ,n1051 ,n821);
    nor g2924(n2125 ,n903 ,n818);
    not g2925(n2124 ,n837);
    not g2926(n838 ,n837);
    not g2927(n836 ,n2124);
    not g2928(n2123 ,n834);
    not g2929(n835 ,n834);
    not g2930(n833 ,n2123);
    not g2931(n2122 ,n831);
    not g2932(n832 ,n831);
    not g2933(n830 ,n2122);
    not g2934(n2121 ,n828);
    not g2935(n829 ,n828);
    not g2936(n827 ,n2121);
    nor g2937(n2120 ,n1444 ,n806);
    nor g2938(n2119 ,n1206 ,n821);
    nor g2939(n2118 ,n1069 ,n821);
    nor g2940(n2117 ,n1065 ,n821);
    nor g2941(n2116 ,n1114 ,n821);
    nor g2942(n2115 ,n1208 ,n821);
    nor g2943(n2114 ,n1121 ,n821);
    nor g2944(n2113 ,n1155 ,n821);
    nor g2945(n2112 ,n1077 ,n821);
    nor g2946(n2111 ,n1102 ,n821);
    nor g2947(n2110 ,n1045 ,n822);
    nor g2948(n2109 ,n1195 ,n821);
    nor g2949(n2108 ,n1128 ,n821);
    nor g2950(n2107 ,n1205 ,n821);
    nor g2951(n2106 ,n1132 ,n822);
    nor g2952(n2105 ,n1127 ,n821);
    nor g2953(n2104 ,n1213 ,n821);
    nor g2954(n2103 ,n1038 ,n821);
    nor g2955(n2102 ,n1080 ,n821);
    nor g2956(n2101 ,n1113 ,n821);
    nor g2957(n2100 ,n1072 ,n821);
    nor g2958(n2099 ,n1196 ,n815);
    nor g2959(n2098 ,n1098 ,n815);
    nor g2960(n2097 ,n1212 ,n815);
    nor g2961(n2096 ,n1070 ,n815);
    nor g2962(n2095 ,n1081 ,n815);
    nor g2963(n2094 ,n1088 ,n815);
    nor g2964(n2093 ,n1122 ,n815);
    nor g2965(n2092 ,n1047 ,n815);
    nor g2966(n2091 ,n1104 ,n815);
    nor g2967(n2090 ,n1109 ,n815);
    nor g2968(n2089 ,n1160 ,n815);
    nor g2969(n2088 ,n1067 ,n815);
    nor g2970(n2087 ,n1100 ,n815);
    nor g2971(n2086 ,n1124 ,n815);
    nor g2972(n2085 ,n1193 ,n815);
    nor g2973(n2084 ,n1148 ,n816);
    nor g2974(n2083 ,n1085 ,n822);
    nor g2975(n2082 ,n1026 ,n815);
    nor g2976(n2081 ,n1204 ,n815);
    nor g2977(n2080 ,n1147 ,n815);
    nor g2978(n2079 ,n1120 ,n815);
    nor g2979(n2078 ,n1099 ,n815);
    nor g2980(n2077 ,n1068 ,n815);
    nor g2981(n2076 ,n1096 ,n815);
    nor g2982(n2075 ,n1129 ,n815);
    nor g2983(n2074 ,n1108 ,n815);
    nor g2984(n2073 ,n1158 ,n815);
    nor g2985(n2072 ,n1063 ,n815);
    nor g2986(n2071 ,n1058 ,n815);
    nor g2987(n2070 ,n1039 ,n815);
    nor g2988(n2069 ,n1165 ,n815);
    nor g2989(n2068 ,n1091 ,n815);
    nor g2990(n2067 ,n1177 ,n822);
    nor g2991(n2066 ,n1187 ,n822);
    nor g2992(n2065 ,n1020 ,n822);
    nor g2993(n2064 ,n1179 ,n822);
    nor g2994(n2063 ,n1034 ,n822);
    nor g2995(n2062 ,n1192 ,n822);
    nor g2996(n2061 ,n1022 ,n822);
    nor g2997(n2060 ,n1135 ,n822);
    nor g2998(n2059 ,n1168 ,n822);
    nor g2999(n2058 ,n1180 ,n822);
    nor g3000(n2057 ,n1117 ,n822);
    nor g3001(n2056 ,n1152 ,n822);
    nor g3002(n2055 ,n1130 ,n822);
    nor g3003(n2054 ,n1040 ,n822);
    nor g3004(n2053 ,n1057 ,n822);
    nor g3005(n2052 ,n1111 ,n822);
    nor g3006(n2051 ,n1140 ,n822);
    nor g3007(n2050 ,n1061 ,n822);
    nor g3008(n2049 ,n1159 ,n822);
    nor g3009(n2048 ,n1095 ,n822);
    nor g3010(n2047 ,n1149 ,n822);
    nor g3011(n2046 ,n1202 ,n822);
    nor g3012(n2045 ,n1046 ,n822);
    nor g3013(n2044 ,n1094 ,n822);
    nor g3014(n2043 ,n1186 ,n822);
    nor g3015(n2042 ,n1073 ,n822);
    nor g3016(n2041 ,n1037 ,n822);
    nor g3017(n2040 ,n1218 ,n816);
    nor g3018(n2039 ,n1092 ,n816);
    nor g3019(n2038 ,n1035 ,n816);
    nor g3020(n2037 ,n1175 ,n816);
    nor g3021(n2036 ,n1075 ,n816);
    nor g3022(n2035 ,n1166 ,n816);
    nor g3023(n2034 ,n1174 ,n816);
    nor g3024(n2033 ,n1141 ,n816);
    nor g3025(n2032 ,n1145 ,n816);
    nor g3026(n2031 ,n1133 ,n816);
    nor g3027(n2030 ,n1101 ,n816);
    nor g3028(n2029 ,n1184 ,n816);
    nor g3029(n2028 ,n1079 ,n816);
    nor g3030(n2027 ,n1142 ,n816);
    nor g3031(n2026 ,n1138 ,n816);
    nor g3032(n2025 ,n1055 ,n816);
    nor g3033(n2024 ,n1198 ,n816);
    nor g3034(n2023 ,n1214 ,n816);
    nor g3035(n2022 ,n1118 ,n816);
    nor g3036(n2021 ,n1164 ,n816);
    nor g3037(n2020 ,n1025 ,n816);
    nor g3038(n2019 ,n1107 ,n816);
    nor g3039(n2018 ,n1146 ,n816);
    nor g3040(n2017 ,n1054 ,n816);
    nor g3041(n2016 ,n1153 ,n816);
    nor g3042(n2015 ,n1023 ,n816);
    nor g3043(n2014 ,n1059 ,n816);
    nor g3044(n2013 ,n1024 ,n816);
    nor g3045(n2012 ,n1027 ,n816);
    nor g3046(n2011 ,n1438 ,n809);
    nor g3047(n2010 ,n1485 ,n808);
    nor g3048(n2009 ,n1488 ,n806);
    nor g3049(n2008 ,n1448 ,n1872);
    nor g3050(n2007 ,n1463 ,n806);
    nor g3051(n2006 ,n1441 ,n807);
    nor g3052(n2005 ,n1588 ,n807);
    nor g3053(n2004 ,n1587 ,n1872);
    nor g3054(n2003 ,n994 ,n809);
    nor g3055(n2002 ,n1002 ,n806);
    nor g3056(n2001 ,n1443 ,n1872);
    nor g3057(n2000 ,n1418 ,n806);
    nor g3058(n1999 ,n1486 ,n1872);
    nor g3059(n1998 ,n1434 ,n806);
    nor g3060(n1997 ,n1526 ,n1872);
    nor g3061(n1996 ,n1209 ,n821);
    nor g3062(n1995 ,n1543 ,n1873);
    nor g3063(n1994 ,n1516 ,n806);
    nor g3064(n1993 ,n1467 ,n1872);
    nor g3065(n1992 ,n992 ,n806);
    nor g3066(n1991 ,n1468 ,n1872);
    nor g3067(n1990 ,n1012 ,n806);
    nor g3068(n1989 ,n1504 ,n1872);
    nor g3069(n1988 ,n1422 ,n809);
    nor g3070(n1987 ,n1567 ,n806);
    nor g3071(n1986 ,n1017 ,n1872);
    nor g3072(n1985 ,n1558 ,n806);
    nor g3073(n1984 ,n1016 ,n1872);
    nor g3074(n1983 ,n1437 ,n1873);
    nor g3075(n1982 ,n1487 ,n806);
    nor g3076(n1981 ,n1577 ,n1872);
    nor g3077(n1980 ,n1427 ,n806);
    nor g3078(n1979 ,n991 ,n808);
    nor g3079(n1978 ,n1481 ,n809);
    nor g3080(n1977 ,n985 ,n1872);
    nor g3081(n1976 ,n968 ,n806);
    nor g3082(n1975 ,n1009 ,n1862);
    nor g3083(n1974 ,n983 ,n1873);
    nor g3084(n1973 ,n1559 ,n1861);
    nor g3085(n1972 ,n1477 ,n1872);
    nor g3086(n1971 ,n1570 ,n806);
    nor g3087(n1970 ,n984 ,n1872);
    nor g3088(n1969 ,n1471 ,n808);
    nor g3089(n1968 ,n1482 ,n1861);
    nor g3090(n1967 ,n998 ,n808);
    nor g3091(n1966 ,n1014 ,n1861);
    nor g3092(n1965 ,n1430 ,n809);
    nor g3093(n1964 ,n1415 ,n808);
    nor g3094(n1963 ,n1554 ,n1861);
    nor g3095(n1962 ,n997 ,n808);
    nor g3096(n1961 ,n1414 ,n1873);
    nor g3097(n1960 ,n1515 ,n1861);
    nor g3098(n1959 ,n981 ,n808);
    nor g3099(n1958 ,n1509 ,n1861);
    nor g3100(n1957 ,n1583 ,n809);
    nor g3101(n1956 ,n982 ,n808);
    nor g3102(n1955 ,n972 ,n1861);
    nor g3103(n1954 ,n1548 ,n808);
    nor g3104(n1953 ,n1547 ,n1861);
    nor g3105(n1952 ,n1576 ,n808);
    nor g3106(n1951 ,n1413 ,n1861);
    nor g3107(n1950 ,n1527 ,n808);
    nor g3108(n1949 ,n1010 ,n807);
    nor g3109(n1948 ,n1495 ,n1861);
    nor g3110(n1947 ,n1426 ,n808);
    nor g3111(n1946 ,n1500 ,n1873);
    nor g3112(n1945 ,n1549 ,n1861);
    nor g3113(n1944 ,n1450 ,n808);
    nor g3114(n1943 ,n1458 ,n1861);
    nor g3115(n1942 ,n1479 ,n808);
    nor g3116(n1941 ,n1435 ,n1861);
    nor g3117(n1940 ,n1464 ,n809);
    nor g3118(n1939 ,n1553 ,n1873);
    nor g3119(n1938 ,n1535 ,n809);
    nor g3120(n1937 ,n1011 ,n1873);
    nor g3121(n1936 ,n1510 ,n808);
    nor g3122(n1935 ,n1529 ,n809);
    nor g3123(n1934 ,n1431 ,n1873);
    nor g3124(n1933 ,n1539 ,n809);
    nor g3125(n1932 ,n1424 ,n1873);
    nor g3126(n1931 ,n1572 ,n806);
    nor g3127(n1930 ,n1439 ,n809);
    nor g3128(n1929 ,n1421 ,n1873);
    nor g3129(n1928 ,n995 ,n809);
    nor g3130(n1927 ,n986 ,n1873);
    nor g3131(n1926 ,n1569 ,n1861);
    nor g3132(n1925 ,n1006 ,n1862);
    nor g3133(n1924 ,n1449 ,n809);
    nor g3134(n1923 ,n1428 ,n807);
    nor g3135(n1922 ,n1525 ,n1862);
    nor g3136(n1921 ,n1425 ,n807);
    nor g3137(n1920 ,n967 ,n1873);
    nor g3138(n1919 ,n1456 ,n1862);
    nor g3139(n1918 ,n1466 ,n807);
    nor g3140(n1917 ,n1555 ,n809);
    nor g3141(n1916 ,n1552 ,n1862);
    nor g3142(n1915 ,n1506 ,n807);
    nor g3143(n1914 ,n970 ,n1862);
    nor g3144(n1913 ,n1461 ,n808);
    nor g3145(n1912 ,n987 ,n807);
    nor g3146(n1911 ,n1004 ,n1873);
    nor g3147(n1910 ,n1519 ,n809);
    nor g3148(n1909 ,n1521 ,n1862);
    nor g3149(n1908 ,n1490 ,n1873);
    nor g3150(n1907 ,n1478 ,n809);
    nor g3151(n1906 ,n1523 ,n807);
    nor g3152(n1905 ,n1423 ,n1862);
    nor g3153(n1904 ,n1501 ,n807);
    nor g3154(n1903 ,n1513 ,n1862);
    nor g3155(n1902 ,n1005 ,n807);
    nor g3156(n1901 ,n1582 ,n808);
    nor g3157(n1900 ,n1412 ,n1862);
    nor g3158(n1899 ,n1565 ,n807);
    nor g3159(n1898 ,n1475 ,n1862);
    nor g3160(n1897 ,n1498 ,n807);
    nor g3161(n1896 ,n973 ,n1862);
    nor g3162(n1895 ,n1019 ,n807);
    nor g3163(n1894 ,n1505 ,n1862);
    nor g3164(n1893 ,n977 ,n807);
    nor g3165(n1892 ,n1507 ,n806);
    nor g3166(n1891 ,n1417 ,n1862);
    nor g3167(n1890 ,n1532 ,n807);
    nor g3168(n1889 ,n1000 ,n809);
    nor g3169(n1888 ,n1496 ,n807);
    or g3170(n1887 ,n1868 ,n1867);
    or g3171(n1886 ,n1865 ,n1866);
    or g3172(n1885 ,n1782 ,n1869);
    or g3173(n1884 ,n1856 ,n1857);
    or g3174(n1883 ,n1870 ,n1871);
    or g3175(n1882 ,n1772 ,n1855);
    or g3176(n1881 ,n1740 ,n1858);
    or g3177(n1880 ,n1796 ,n1860);
    nor g3178(n1879 ,n131 ,n1862);
    nor g3179(n1878 ,n130 ,n1873);
    nor g3180(n1877 ,n129 ,n1861);
    nor g3181(n1876 ,n128 ,n1872);
    nor g3182(n837 ,n839 ,n821);
    nor g3183(n834 ,n813 ,n815);
    nor g3184(n831 ,n839 ,n822);
    nor g3185(n828 ,n810 ,n816);
    not g3186(n825 ,n1875);
    not g3187(n826 ,n1875);
    not g3188(n823 ,n1874);
    not g3189(n824 ,n1874);
    or g3190(n1871 ,n1803 ,n1809);
    or g3191(n1870 ,n1497 ,n1823);
    or g3192(n1869 ,n1808 ,n1819);
    or g3193(n1868 ,n1520 ,n1811);
    or g3194(n1867 ,n1824 ,n1822);
    or g3195(n1866 ,n1818 ,n1817);
    or g3196(n1865 ,n1460 ,n1825);
    nor g3197(n1875 ,n871 ,n803);
    nor g3198(n1874 ,n871 ,n1802);
    nor g3199(n1873 ,n871 ,n804);
    nor g3200(n1872 ,n871 ,n805);
    not g3201(n819 ,n1864);
    not g3202(n820 ,n1864);
    not g3203(n817 ,n1863);
    not g3204(n818 ,n1863);
    or g3205(n1860 ,n1737 ,n1826);
    or g3206(n1859 ,n1816 ,n1815);
    or g3207(n1858 ,n1820 ,n1804);
    or g3208(n1857 ,n1807 ,n1812);
    or g3209(n1856 ,n1813 ,n1805);
    or g3210(n1855 ,n1853 ,n1810);
    nor g3211(n1854 ,n799 ,n1799);
    nor g3212(n1864 ,n6[5] ,n1801);
    nor g3213(n1863 ,n37[0] ,n803);
    nor g3214(n1862 ,n37[0] ,n804);
    nor g3215(n1861 ,n37[0] ,n805);
    or g3216(n1853 ,n1779 ,n1780);
    nor g3217(n1852 ,n1087 ,n1765);
    nor g3218(n1851 ,n1106 ,n1765);
    nor g3219(n1850 ,n1044 ,n1765);
    nor g3220(n1849 ,n1049 ,n1765);
    nor g3221(n1848 ,n1125 ,n1765);
    nor g3222(n1847 ,n1157 ,n1765);
    nor g3223(n1846 ,n1197 ,n1765);
    nor g3224(n1845 ,n1084 ,n1765);
    nor g3225(n1844 ,n1156 ,n1765);
    nor g3226(n1843 ,n1093 ,n1765);
    nor g3227(n1842 ,n1086 ,n1765);
    nor g3228(n1841 ,n1031 ,n1765);
    nor g3229(n1840 ,n1032 ,n1765);
    nor g3230(n1839 ,n1144 ,n1765);
    nor g3231(n1838 ,n1074 ,n1765);
    nor g3232(n1837 ,n1219 ,n1765);
    nor g3233(n1836 ,n1161 ,n1765);
    nor g3234(n1835 ,n1150 ,n1765);
    nor g3235(n1834 ,n1207 ,n1765);
    nor g3236(n1833 ,n1115 ,n1765);
    nor g3237(n1832 ,n1066 ,n1765);
    nor g3238(n1831 ,n1089 ,n1765);
    nor g3239(n1830 ,n1188 ,n1765);
    nor g3240(n1829 ,n1190 ,n1765);
    nor g3241(n1828 ,n1082 ,n1765);
    nor g3242(n1827 ,n1154 ,n1765);
    nor g3243(n1826 ,n1018 ,n1768);
    or g3244(n1825 ,n1777 ,n1776);
    or g3245(n1824 ,n1775 ,n1789);
    or g3246(n1823 ,n1788 ,n1792);
    or g3247(n1822 ,n1786 ,n1785);
    or g3248(n1821 ,n1784 ,n1783);
    or g3249(n1820 ,n1787 ,n1750);
    or g3250(n1819 ,n1751 ,n1778);
    or g3251(n1818 ,n1774 ,n1794);
    or g3252(n1817 ,n1755 ,n1760);
    or g3253(n1816 ,n1762 ,n1770);
    or g3254(n1815 ,n1769 ,n1797);
    or g3255(n1814 ,n1773 ,n1771);
    or g3256(n1813 ,n1781 ,n1761);
    or g3257(n1812 ,n1749 ,n1763);
    or g3258(n1811 ,n1791 ,n1758);
    or g3259(n1810 ,n1790 ,n1795);
    or g3260(n1809 ,n1753 ,n1752);
    or g3261(n1808 ,n1747 ,n1748);
    or g3262(n1807 ,n1745 ,n1757);
    or g3263(n1806 ,n1741 ,n1742);
    or g3264(n1805 ,n1759 ,n1744);
    or g3265(n1804 ,n1743 ,n1746);
    or g3266(n1803 ,n1793 ,n1754);
    or g3267(n1802 ,n6[5] ,n1766);
    or g3268(n1801 ,n37[0] ,n1766);
    nor g3269(n1800 ,n6[5] ,n1765);
    nor g3270(n1799 ,n12 ,n1767);
    or g3271(n1797 ,n1663 ,n1686);
    nor g3272(n1796 ,n4464 ,n1734);
    or g3273(n1795 ,n1666 ,n1644);
    or g3274(n1794 ,n1681 ,n1715);
    or g3275(n1793 ,n1709 ,n1712);
    or g3276(n1792 ,n1710 ,n1651);
    or g3277(n1791 ,n1701 ,n1700);
    or g3278(n1790 ,n1638 ,n1670);
    or g3279(n1789 ,n1699 ,n1713);
    or g3280(n1788 ,n1630 ,n1652);
    or g3281(n1787 ,n1706 ,n1689);
    or g3282(n1786 ,n1693 ,n1692);
    or g3283(n1785 ,n1691 ,n1642);
    or g3284(n1784 ,n1690 ,n1718);
    or g3285(n1783 ,n1719 ,n1720);
    or g3286(n1782 ,n1721 ,n1723);
    or g3287(n1781 ,n1702 ,n1622);
    or g3288(n1780 ,n1726 ,n1671);
    or g3289(n1779 ,n1703 ,n1635);
    or g3290(n1778 ,n1664 ,n1677);
    or g3291(n1777 ,n1624 ,n1727);
    or g3292(n1776 ,n1685 ,n1684);
    or g3293(n1775 ,n1696 ,n1694);
    or g3294(n1774 ,n1711 ,n1682);
    or g3295(n1773 ,n1676 ,n1675);
    or g3296(n1772 ,n1668 ,n1655);
    or g3297(n1771 ,n1667 ,n1673);
    or g3298(n1770 ,n1665 ,n1669);
    or g3299(n1769 ,n1672 ,n1647);
    or g3300(n1798 ,n1018 ,n1735);
    not g3301(n1768 ,n1767);
    not g3302(n1765 ,n1764);
    or g3303(n1763 ,n1725 ,n1688);
    or g3304(n1762 ,n1662 ,n1674);
    or g3305(n1761 ,n1623 ,n1625);
    or g3306(n1760 ,n1678 ,n1683);
    or g3307(n1759 ,n1627 ,n1660);
    or g3308(n1758 ,n1698 ,n1697);
    or g3309(n1757 ,n1636 ,n1657);
    or g3310(n1756 ,n1658 ,n1661);
    or g3311(n1755 ,n1680 ,n1679);
    or g3312(n1754 ,n1714 ,n1650);
    or g3313(n1753 ,n1626 ,n1621);
    or g3314(n1752 ,n1705 ,n1646);
    or g3315(n1751 ,n1649 ,n1687);
    or g3316(n1750 ,n1707 ,n1641);
    or g3317(n1749 ,n1639 ,n1656);
    or g3318(n1748 ,n1637 ,n1654);
    or g3319(n1747 ,n1634 ,n1724);
    or g3320(n1746 ,n1631 ,n1704);
    or g3321(n1745 ,n1633 ,n1632);
    or g3322(n1744 ,n1629 ,n1659);
    or g3323(n1743 ,n1640 ,n1695);
    or g3324(n1742 ,n1648 ,n1643);
    or g3325(n1741 ,n1628 ,n1645);
    or g3326(n1740 ,n1653 ,n1708);
    or g3327(n1739 ,n1732 ,n1728);
    or g3328(n1738 ,n1732 ,n1730);
    nor g3329(n1737 ,n1600 ,n1731);
    nor g3330(n1736 ,n1605 ,n1732);
    nor g3331(n1767 ,n1717 ,n1732);
    or g3332(n1766 ,n814 ,n1734);
    nor g3333(n1764 ,n811 ,n1722);
    not g3334(n1734 ,n1733);
    not g3335(n1731 ,n1730);
    not g3336(n1729 ,n1728);
    xnor g3337(n1727 ,n6[8] ,n921);
    xnor g3338(n1726 ,n6[27] ,n899);
    xnor g3339(n1725 ,n6[7] ,n887);
    xnor g3340(n1724 ,n6[28] ,n1273);
    xnor g3341(n1723 ,n6[30] ,n902);
    or g3342(n1722 ,n872 ,n1602);
    xnor g3343(n1721 ,n6[31] ,n908);
    xnor g3344(n1720 ,n6[6] ,n1270);
    xnor g3345(n1719 ,n6[7] ,n1241);
    xnor g3346(n1718 ,n6[8] ,n897);
    nor g3347(n1717 ,n33[2] ,n1603);
    or g3348(n1716 ,n33[2] ,n1601);
    xnor g3349(n1715 ,n6[18] ,n1281);
    xnor g3350(n1714 ,n6[15] ,n935);
    xnor g3351(n1713 ,n6[14] ,n1255);
    xnor g3352(n1712 ,n6[16] ,n1246);
    xnor g3353(n1711 ,n6[21] ,n1249);
    xnor g3354(n1710 ,n6[7] ,n1292);
    xnor g3355(n1709 ,n6[17] ,n924);
    xnor g3356(n1708 ,n6[30] ,n917);
    xnor g3357(n1707 ,n6[27] ,n1291);
    xnor g3358(n1706 ,n6[29] ,n1243);
    xnor g3359(n1705 ,n6[11] ,n1244);
    xnor g3360(n1704 ,n6[22] ,n928);
    xnor g3361(n1703 ,n6[29] ,n1263);
    xnor g3362(n1702 ,n6[21] ,n1296);
    xnor g3363(n1701 ,n6[21] ,n1288);
    xnor g3364(n1700 ,n6[20] ,n926);
    xnor g3365(n1699 ,n6[15] ,n892);
    xnor g3366(n1698 ,n6[19] ,n1261);
    xnor g3367(n1697 ,n6[18] ,n1223);
    xnor g3368(n1696 ,n6[17] ,n1233);
    xnor g3369(n1695 ,n6[24] ,n1278);
    xnor g3370(n1694 ,n6[16] ,n1224);
    xnor g3371(n1693 ,n6[13] ,n1247);
    xnor g3372(n1692 ,n6[12] ,n1257);
    xnor g3373(n1691 ,n6[11] ,n1248);
    xnor g3374(n1690 ,n6[9] ,n903);
    xnor g3375(n1689 ,n6[28] ,n1286);
    or g3376(n1735 ,n33[2] ,n1604);
    nor g3377(n1733 ,n33[2] ,n1593);
    nor g3378(n1732 ,n872 ,n1601);
    nor g3379(n1730 ,n33[2] ,n1602);
    nor g3380(n1728 ,n1221 ,n1606);
    xnor g3381(n1688 ,n6[6] ,n1254);
    xnor g3382(n1687 ,n6[24] ,n1264);
    xnor g3383(n1686 ,n6[22] ,n1232);
    xnor g3384(n1685 ,n6[7] ,n1272);
    xnor g3385(n1684 ,n6[6] ,n1295);
    xnor g3386(n1683 ,n6[14] ,n1280);
    xnor g3387(n1682 ,n6[20] ,n913);
    xnor g3388(n1681 ,n6[19] ,n1260);
    xnor g3389(n1680 ,n6[17] ,n900);
    xnor g3390(n1679 ,n6[16] ,n886);
    xnor g3391(n1678 ,n6[15] ,n1250);
    xnor g3392(n1677 ,n6[22] ,n1293);
    xnor g3393(n1676 ,n6[13] ,n1256);
    xnor g3394(n1675 ,n6[12] ,n880);
    xnor g3395(n1674 ,n6[28] ,n874);
    xnor g3396(n1673 ,n6[10] ,n1290);
    xnor g3397(n1672 ,n6[25] ,n929);
    xnor g3398(n1671 ,n6[26] ,n1230);
    xnor g3399(n1670 ,n6[24] ,n1242);
    xnor g3400(n1669 ,n6[26] ,n894);
    xnor g3401(n1668 ,n6[31] ,n1245);
    xnor g3402(n1667 ,n6[11] ,n1236);
    xnor g3403(n1666 ,n6[23] ,n1225);
    xnor g3404(n1665 ,n6[27] ,n1271);
    xnor g3405(n1664 ,n6[23] ,n1279);
    xnor g3406(n1663 ,n6[23] ,n1285);
    xnor g3407(n1662 ,n6[29] ,n882);
    xnor g3408(n1661 ,n6[30] ,n1239);
    xnor g3409(n1660 ,n6[16] ,n1238);
    xnor g3410(n1659 ,n6[14] ,n925);
    xnor g3411(n1658 ,n6[31] ,n1258);
    xnor g3412(n1657 ,n6[10] ,n1267);
    xnor g3413(n1656 ,n6[8] ,n909);
    xnor g3414(n1655 ,n6[30] ,n918);
    xnor g3415(n1654 ,n6[26] ,n1235);
    xnor g3416(n1653 ,n6[31] ,n1253);
    xnor g3417(n1652 ,n6[8] ,n1226);
    xnor g3418(n1651 ,n6[6] ,n1240);
    xnor g3419(n1650 ,n6[14] ,n1284);
    xnor g3420(n1649 ,n6[25] ,n1252);
    xnor g3421(n1648 ,n6[19] ,n1265);
    xnor g3422(n1647 ,n6[24] ,n1294);
    xnor g3423(n1646 ,n6[10] ,n916);
    xnor g3424(n1645 ,n6[20] ,n901);
    xnor g3425(n1644 ,n6[22] ,n1266);
    xnor g3426(n1643 ,n6[18] ,n884);
    xnor g3427(n1642 ,n6[10] ,n1229);
    xnor g3428(n1641 ,n6[26] ,n890);
    xnor g3429(n1640 ,n6[25] ,n1268);
    xnor g3430(n1639 ,n6[9] ,n920);
    xnor g3431(n1638 ,n6[25] ,n1251);
    xnor g3432(n1637 ,n6[27] ,n1275);
    xnor g3433(n1636 ,n6[11] ,n1274);
    xnor g3434(n1635 ,n6[28] ,n1237);
    xnor g3435(n1634 ,n6[29] ,n1262);
    xnor g3436(n1633 ,n6[13] ,n1287);
    xnor g3437(n1632 ,n6[12] ,n1297);
    xnor g3438(n1631 ,n6[23] ,n1231);
    xnor g3439(n1630 ,n6[9] ,n1276);
    xnor g3440(n1629 ,n6[15] ,n1283);
    xnor g3441(n1628 ,n6[21] ,n1227);
    xnor g3442(n1627 ,n6[17] ,n934);
    xnor g3443(n1626 ,n6[13] ,n1269);
    xnor g3444(n1625 ,n6[18] ,n1277);
    xnor g3445(n1624 ,n6[9] ,n1282);
    xnor g3446(n1623 ,n6[19] ,n1228);
    xnor g3447(n1622 ,n6[20] ,n1289);
    xnor g3448(n1621 ,n6[12] ,n1234);
    nor g3449(n1620 ,n1259 ,n813);
    nor g3450(n1619 ,n1546 ,n814);
    nor g3451(n1618 ,n953 ,n799);
    nor g3452(n1617 ,n1410 ,n814);
    nor g3453(n1616 ,n1396 ,n813);
    nor g3454(n1615 ,n1380 ,n810);
    nor g3455(n1614 ,n1304 ,n810);
    nor g3456(n1613 ,n943 ,n814);
    nor g3457(n1612 ,n1335 ,n799);
    nor g3458(n1611 ,n888 ,n839);
    nor g3459(n1610 ,n1003 ,n813);
    nor g3460(n1609 ,n1301 ,n813);
    nor g3461(n1608 ,n1377 ,n814);
    nor g3462(n1607 ,n1348 ,n810);
    not g3463(n1606 ,n1605);
    not g3464(n1604 ,n1603);
    not g3465(n1602 ,n1601);
    nor g3466(n1600 ,n2 ,n3);
    nor g3467(n1599 ,n1528 ,n813);
    nor g3468(n1598 ,n951 ,n814);
    nor g3469(n1597 ,n1341 ,n814);
    nor g3470(n1596 ,n949 ,n814);
    nor g3471(n1595 ,n1343 ,n810);
    nor g3472(n1594 ,n1299 ,n813);
    or g3473(n1593 ,n1221 ,n1222);
    nor g3474(n1592 ,n1222 ,n813);
    nor g3475(n1591 ,n1401 ,n813);
    nor g3476(n1590 ,n1221 ,n810);
    nor g3477(n1605 ,n33[1] ,n33[2]);
    nor g3478(n1603 ,n1222 ,n33[0]);
    nor g3479(n1601 ,n33[0] ,n33[1]);
    not g3480(n1589 ,n10[8]);
    not g3481(n1588 ,n23[31]);
    not g3482(n1587 ,n21[1]);
    not g3483(n1586 ,n10[27]);
    not g3484(n1585 ,n9[8]);
    not g3485(n1584 ,n11[31]);
    not g3486(n1583 ,n24[23]);
    not g3487(n1582 ,n22[30]);
    not g3488(n1581 ,n11[24]);
    not g3489(n1580 ,n130);
    not g3490(n1579 ,n9[7]);
    not g3491(n1578 ,n11[14]);
    not g3492(n1577 ,n21[21]);
    not g3493(n1576 ,n22[17]);
    not g3494(n1575 ,n9[18]);
    not g3495(n1574 ,n9[28]);
    not g3496(n1573 ,n9[4]);
    not g3497(n1572 ,n21[14]);
    not g3498(n1571 ,n11[13]);
    not g3499(n1570 ,n21[29]);
    not g3500(n1569 ,n22[10]);
    not g3501(n1568 ,n9[24]);
    not g3502(n1567 ,n21[16]);
    not g3503(n1566 ,n11[2]);
    not g3504(n1565 ,n23[14]);
    not g3505(n1564 ,n11[12]);
    not g3506(n1563 ,n10[14]);
    not g3507(n1562 ,n11[23]);
    not g3508(n1561 ,n9[13]);
    not g3509(n1560 ,n9[27]);
    not g3510(n1559 ,n22[24]);
    not g3511(n1558 ,n21[18]);
    not g3512(n1557 ,n9[26]);
    not g3513(n1556 ,n10[6]);
    not g3514(n1555 ,n24[11]);
    not g3515(n1554 ,n22[7]);
    not g3516(n1553 ,n24[19]);
    not g3517(n1552 ,n23[16]);
    not g3518(n1551 ,n10[3]);
    not g3519(n1550 ,n11[15]);
    not g3520(n1549 ,n22[25]);
    not g3521(n1548 ,n22[15]);
    not g3522(n1547 ,n22[16]);
    not g3523(n1546 ,n36[0]);
    not g3524(n1545 ,n11[22]);
    not g3525(n1544 ,n10[23]);
    not g3526(n1543 ,n24[31]);
    not g3527(n1542 ,n10[19]);
    not g3528(n1541 ,n11[0]);
    not g3529(n1540 ,n9[5]);
    not g3530(n1539 ,n24[16]);
    not g3531(n1538 ,n11[20]);
    not g3532(n1537 ,n9[23]);
    not g3533(n1536 ,n11[18]);
    not g3534(n1535 ,n24[18]);
    not g3535(n1534 ,n9[16]);
    not g3536(n1533 ,n9[3]);
    not g3537(n1532 ,n23[2]);
    not g3538(n1531 ,n9[6]);
    not g3539(n1530 ,n10[30]);
    not g3540(n1529 ,n24[12]);
    not g3541(n1528 ,n36[2]);
    not g3542(n1527 ,n22[19]);
    not g3543(n1526 ,n21[7]);
    not g3544(n1525 ,n23[8]);
    not g3545(n1524 ,n14);
    not g3546(n1523 ,n23[22]);
    not g3547(n1522 ,n9[22]);
    not g3548(n1521 ,n23[24]);
    not g3549(n1520 ,n131);
    not g3550(n1519 ,n24[7]);
    not g3551(n1518 ,n11[9]);
    not g3552(n1517 ,n10[5]);
    not g3553(n1516 ,n21[9]);
    not g3554(n1515 ,n22[9]);
    not g3555(n1514 ,n11[4]);
    not g3556(n1513 ,n23[19]);
    not g3557(n1512 ,n10[18]);
    not g3558(n1511 ,n9[25]);
    not g3559(n1510 ,n22[14]);
    not g3560(n1509 ,n22[11]);
    not g3561(n1508 ,n10[31]);
    not g3562(n1507 ,n21[22]);
    not g3563(n1506 ,n23[20]);
    not g3564(n1505 ,n23[6]);
    not g3565(n1504 ,n21[15]);
    not g3566(n1503 ,n10[16]);
    not g3567(n1502 ,n10[0]);
    not g3568(n1501 ,n23[21]);
    not g3569(n1500 ,n24[22]);
    not g3570(n1499 ,n10[10]);
    not g3571(n1498 ,n23[11]);
    not g3572(n1497 ,n128);
    not g3573(n1496 ,n23[1]);
    not g3574(n1495 ,n22[20]);
    not g3575(n1494 ,n10[21]);
    not g3576(n1493 ,n9[0]);
    not g3577(n1492 ,n11[6]);
    not g3578(n1491 ,n11[5]);
    not g3579(n1490 ,n24[3]);
    not g3580(n1489 ,n11[27]);
    not g3581(n1488 ,n21[30]);
    not g3582(n1487 ,n21[20]);
    not g3583(n1486 ,n21[5]);
    not g3584(n1485 ,n22[2]);
    not g3585(n1484 ,n11[10]);
    not g3586(n1483 ,n9[11]);
    not g3587(n1482 ,n22[3]);
    not g3588(n1481 ,n24[13]);
    not g3589(n1480 ,n10[12]);
    not g3590(n1479 ,n22[29]);
    not g3591(n1478 ,n24[21]);
    not g3592(n1477 ,n21[28]);
    not g3593(n1476 ,n9[2]);
    not g3594(n1475 ,n23[10]);
    not g3595(n1474 ,n15);
    not g3596(n1473 ,n9[20]);
    not g3597(n1472 ,n9[1]);
    not g3598(n1471 ,n22[1]);
    not g3599(n1470 ,n10[1]);
    not g3600(n1469 ,n9[31]);
    not g3601(n1468 ,n21[12]);
    not g3602(n1467 ,n21[10]);
    not g3603(n1466 ,n23[13]);
    not g3604(n1465 ,n11[11]);
    not g3605(n1464 ,n24[1]);
    not g3606(n1463 ,n21[26]);
    not g3607(n1462 ,n10[22]);
    not g3608(n1461 ,n22[6]);
    not g3609(n1460 ,n129);
    not g3610(n1459 ,n10[11]);
    not g3611(n1458 ,n22[28]);
    not g3612(n1457 ,n11[19]);
    not g3613(n1456 ,n23[12]);
    not g3614(n1455 ,n11[21]);
    not g3615(n1454 ,n11[8]);
    not g3616(n1453 ,n11[26]);
    not g3617(n1452 ,n9[17]);
    not g3618(n1451 ,n10[20]);
    not g3619(n1450 ,n22[27]);
    not g3620(n1449 ,n24[5]);
    not g3621(n1448 ,n21[27]);
    not g3622(n1447 ,n10[15]);
    not g3623(n1446 ,n10[7]);
    not g3624(n1445 ,n9[12]);
    not g3625(n1444 ,n21[8]);
    not g3626(n1443 ,n21[3]);
    not g3627(n1442 ,n9[10]);
    not g3628(n1441 ,n23[30]);
    not g3629(n1440 ,n11[17]);
    not g3630(n1439 ,n24[25]);
    not g3631(n1438 ,n24[4]);
    not g3632(n1437 ,n24[29]);
    not g3633(n1436 ,n10[9]);
    not g3634(n1435 ,n22[31]);
    not g3635(n1434 ,n21[6]);
    not g3636(n1433 ,n10[25]);
    not g3637(n1432 ,n9[30]);
    not g3638(n1431 ,n24[17]);
    not g3639(n1430 ,n24[26]);
    not g3640(n1429 ,n11[29]);
    not g3641(n1428 ,n23[5]);
    not g3642(n1427 ,n21[23]);
    not g3643(n1426 ,n22[21]);
    not g3644(n1425 ,n23[9]);
    not g3645(n1424 ,n24[20]);
    not g3646(n1423 ,n23[17]);
    not g3647(n1422 ,n24[30]);
    not g3648(n1421 ,n24[15]);
    not g3649(n1420 ,n10[29]);
    not g3650(n1419 ,n10[2]);
    not g3651(n1418 ,n21[4]);
    not g3652(n1417 ,n23[3]);
    not g3653(n1416 ,n9[14]);
    not g3654(n1415 ,n22[5]);
    not g3655(n1414 ,n24[24]);
    not g3656(n1413 ,n22[18]);
    not g3657(n1412 ,n23[15]);
    not g3658(n1411 ,n11[28]);
    not g3659(n1410 ,n35[1]);
    not g3660(n1409 ,n25[26]);
    not g3661(n1408 ,n28[13]);
    not g3662(n1407 ,n28[15]);
    not g3663(n1406 ,n27[19]);
    not g3664(n1405 ,n26[29]);
    not g3665(n1404 ,n28[24]);
    not g3666(n1403 ,n28[10]);
    not g3667(n1402 ,n28[27]);
    not g3668(n1401 ,n34[4]);
    not g3669(n1400 ,n26[28]);
    not g3670(n1399 ,n28[28]);
    not g3671(n1398 ,n26[16]);
    not g3672(n1397 ,n28[31]);
    not g3673(n1396 ,n34[6]);
    not g3674(n1395 ,n26[9]);
    not g3675(n1394 ,n28[4]);
    not g3676(n1393 ,n27[1]);
    not g3677(n1392 ,n25[1]);
    not g3678(n1391 ,n26[3]);
    not g3679(n1390 ,n25[7]);
    not g3680(n1389 ,n27[5]);
    not g3681(n1388 ,n25[3]);
    not g3682(n1387 ,n25[10]);
    not g3683(n1386 ,n27[23]);
    not g3684(n1385 ,n28[18]);
    not g3685(n1384 ,n25[9]);
    not g3686(n1383 ,n25[6]);
    not g3687(n1382 ,n27[14]);
    not g3688(n1381 ,n26[8]);
    not g3689(n1380 ,n34[7]);
    not g3690(n1379 ,n26[6]);
    not g3691(n1378 ,n27[17]);
    not g3692(n1377 ,n16);
    not g3693(n1376 ,n26[17]);
    not g3694(n1375 ,n27[16]);
    not g3695(n1374 ,n28[19]);
    not g3696(n1373 ,n28[23]);
    not g3697(n1372 ,n28[8]);
    not g3698(n1371 ,n28[26]);
    not g3699(n1370 ,n27[7]);
    not g3700(n1369 ,n25[30]);
    not g3701(n1368 ,n28[5]);
    not g3702(n1367 ,n26[24]);
    not g3703(n1366 ,n27[0]);
    not g3704(n1365 ,n27[26]);
    not g3705(n1364 ,n28[25]);
    not g3706(n1363 ,n26[5]);
    not g3707(n1362 ,n26[7]);
    not g3708(n1361 ,n26[14]);
    not g3709(n1360 ,n28[9]);
    not g3710(n1359 ,n25[21]);
    not g3711(n1358 ,n28[11]);
    not g3712(n1357 ,n25[13]);
    not g3713(n1356 ,n26[11]);
    not g3714(n1355 ,n25[8]);
    not g3715(n1354 ,n27[3]);
    not g3716(n1353 ,n25[11]);
    not g3717(n1352 ,n27[27]);
    not g3718(n1351 ,n25[18]);
    not g3719(n1350 ,n27[24]);
    not g3720(n1349 ,n26[15]);
    not g3721(n1348 ,n34[2]);
    not g3722(n1347 ,n27[22]);
    not g3723(n1346 ,n27[10]);
    not g3724(n1345 ,n26[30]);
    not g3725(n1344 ,n26[22]);
    not g3726(n1343 ,n35[7]);
    not g3727(n1342 ,n25[20]);
    not g3728(n1341 ,n34[3]);
    not g3729(n1340 ,n27[2]);
    not g3730(n1339 ,n27[20]);
    not g3731(n1338 ,n25[17]);
    not g3732(n1337 ,n28[22]);
    not g3733(n1336 ,n26[27]);
    not g3734(n1335 ,n35[3]);
    not g3735(n1334 ,n27[12]);
    not g3736(n1333 ,n28[0]);
    not g3737(n1332 ,n25[28]);
    not g3738(n1331 ,n26[12]);
    not g3739(n1330 ,n25[23]);
    not g3740(n1329 ,n28[3]);
    not g3741(n1328 ,n28[20]);
    not g3742(n1327 ,n25[31]);
    not g3743(n1326 ,n25[2]);
    not g3744(n1325 ,n28[7]);
    not g3745(n1324 ,n26[0]);
    not g3746(n1323 ,n28[29]);
    not g3747(n1322 ,n25[27]);
    not g3748(n1321 ,n26[20]);
    not g3749(n1320 ,n28[17]);
    not g3750(n1319 ,n27[9]);
    not g3751(n1318 ,n26[4]);
    not g3752(n1317 ,n26[21]);
    not g3753(n1316 ,n27[13]);
    not g3754(n1315 ,n27[6]);
    not g3755(n1314 ,n28[6]);
    not g3756(n1313 ,n25[25]);
    not g3757(n1312 ,n27[28]);
    not g3758(n1311 ,n25[22]);
    not g3759(n1310 ,n26[19]);
    not g3760(n1309 ,n27[4]);
    not g3761(n1308 ,n27[11]);
    not g3762(n1307 ,n25[14]);
    not g3763(n1306 ,n27[30]);
    not g3764(n1305 ,n26[31]);
    not g3765(n1304 ,n35[4]);
    not g3766(n1303 ,n25[19]);
    not g3767(n1302 ,n26[23]);
    not g3768(n1301 ,n17);
    not g3769(n1300 ,n26[10]);
    not g3770(n1299 ,n35[2]);
    not g3771(n1298 ,n28[16]);
    not g3772(n1297 ,n31[6]);
    not g3773(n1296 ,n31[15]);
    not g3774(n1295 ,n30[0]);
    not g3775(n1294 ,n31[18]);
    not g3776(n1293 ,n32[16]);
    not g3777(n1292 ,n29[1]);
    not g3778(n1291 ,n29[21]);
    not g3779(n1290 ,n30[4]);
    not g3780(n1289 ,n31[14]);
    not g3781(n1288 ,n32[15]);
    not g3782(n1287 ,n31[7]);
    not g3783(n1286 ,n29[22]);
    not g3784(n1285 ,n31[17]);
    not g3785(n1284 ,n29[8]);
    not g3786(n1283 ,n31[9]);
    not g3787(n1282 ,n30[3]);
    not g3788(n1281 ,n30[12]);
    not g3789(n1280 ,n30[8]);
    not g3790(n1279 ,n32[17]);
    not g3791(n1278 ,n29[18]);
    not g3792(n1277 ,n31[12]);
    not g3793(n1276 ,n29[3]);
    not g3794(n1275 ,n32[21]);
    not g3795(n1274 ,n31[5]);
    not g3796(n1273 ,n32[22]);
    not g3797(n1272 ,n30[1]);
    not g3798(n1271 ,n31[21]);
    not g3799(n1270 ,n32[0]);
    not g3800(n1269 ,n29[7]);
    not g3801(n1268 ,n29[19]);
    not g3802(n1267 ,n31[4]);
    not g3803(n1266 ,n30[16]);
    not g3804(n1265 ,n29[13]);
    not g3805(n1264 ,n32[18]);
    not g3806(n1263 ,n30[23]);
    not g3807(n1262 ,n32[23]);
    not g3808(n1261 ,n32[13]);
    not g3809(n1260 ,n30[13]);
    not g3810(n1259 ,n35[0]);
    not g3811(n1258 ,n31[25]);
    not g3812(n1257 ,n32[6]);
    not g3813(n1256 ,n30[7]);
    not g3814(n1255 ,n32[8]);
    not g3815(n1254 ,n31[0]);
    not g3816(n1253 ,n29[25]);
    not g3817(n1252 ,n32[19]);
    not g3818(n1251 ,n30[19]);
    not g3819(n1250 ,n30[9]);
    not g3820(n1249 ,n30[15]);
    not g3821(n1248 ,n32[5]);
    not g3822(n1247 ,n32[7]);
    not g3823(n1246 ,n29[10]);
    not g3824(n1245 ,n30[25]);
    not g3825(n1244 ,n29[5]);
    not g3826(n1243 ,n29[23]);
    not g3827(n1242 ,n30[18]);
    not g3828(n1241 ,n32[1]);
    not g3829(n1240 ,n29[0]);
    not g3830(n1239 ,n31[24]);
    not g3831(n1238 ,n31[10]);
    not g3832(n1237 ,n30[22]);
    not g3833(n1236 ,n30[5]);
    not g3834(n1235 ,n32[20]);
    not g3835(n1234 ,n29[6]);
    not g3836(n1233 ,n32[11]);
    not g3837(n1232 ,n31[16]);
    not g3838(n1231 ,n29[17]);
    not g3839(n1230 ,n30[20]);
    not g3840(n1229 ,n32[4]);
    not g3841(n1228 ,n31[13]);
    not g3842(n1227 ,n29[15]);
    not g3843(n1226 ,n29[2]);
    not g3844(n1225 ,n30[17]);
    not g3845(n1224 ,n32[10]);
    not g3846(n1223 ,n32[12]);
    not g3847(n1222 ,n33[1]);
    not g3848(n1221 ,n33[0]);
    not g3849(n1220 ,n7[26]);
    not g3850(n1219 ,n4483);
    not g3851(n1218 ,n4585);
    not g3852(n1217 ,n7[11]);
    not g3853(n1216 ,n7[23]);
    not g3854(n1215 ,n4674);
    not g3855(n1214 ,n4562);
    not g3856(n1213 ,n4653);
    not g3857(n1212 ,n4646);
    not g3858(n1211 ,n4683);
    not g3859(n1210 ,n7[18]);
    not g3860(n1209 ,n4667);
    not g3861(n1208 ,n4662);
    not g3862(n1207 ,n4479);
    not g3863(n1206 ,n4666);
    not g3864(n1205 ,n4655);
    not g3865(n1204 ,n4632);
    not g3866(n1203 ,n7[3]);
    not g3867(n1202 ,n4596);
    not g3868(n1201 ,n4620);
    not g3869(n1200 ,n4690);
    not g3870(n1199 ,n4684);
    not g3871(n1198 ,n4563);
    not g3872(n1197 ,n4490);
    not g3873(n1196 ,n4648);
    not g3874(n1195 ,n4657);
    not g3875(n1194 ,n7[21]);
    not g3876(n1193 ,n4634);
    not g3877(n1192 ,n4612);
    not g3878(n1191 ,n4688);
    not g3879(n1190 ,n4480);
    not g3880(n1189 ,n4677);
    not g3881(n1188 ,n4487);
    not g3882(n1187 ,n4616);
    not g3883(n1186 ,n4591);
    not g3884(n1185 ,n4678);
    not g3885(n1184 ,n4572);
    not g3886(n1183 ,n4682);
    not g3887(n1182 ,n7[14]);
    not g3888(n1181 ,n7[16]);
    not g3889(n1180 ,n4608);
    not g3890(n1179 ,n4614);
    not g3891(n1178 ,n7[9]);
    not g3892(n1177 ,n4617);
    not g3893(n1176 ,n4673);
    not g3894(n1175 ,n4582);
    not g3895(n1174 ,n4579);
    not g3896(n1173 ,n7[2]);
    not g3897(n1172 ,n4686);
    not g3898(n1171 ,n6[0]);
    not g3899(n1170 ,n7[22]);
    not g3900(n1169 ,n4671);
    not g3901(n1168 ,n4609);
    not g3902(n1167 ,n7[28]);
    not g3903(n1166 ,n4580);
    not g3904(n1165 ,n4619);
    not g3905(n1164 ,n4560);
    not g3906(n1163 ,n7[30]);
    not g3907(n1162 ,n7[6]);
    not g3908(n1161 ,n4475);
    not g3909(n1160 ,n4638);
    not g3910(n1159 ,n4599);
    not g3911(n1158 ,n4624);
    not g3912(n1157 ,n4477);
    not g3913(n1156 ,n4485);
    not g3914(n1155 ,n4660);
    not g3915(n1154 ,n4470);
    not g3916(n1153 ,n4570);
    not g3917(n1152 ,n4606);
    not g3918(n1151 ,n7[0]);
    not g3919(n1150 ,n4478);
    not g3920(n1149 ,n4597);
    not g3921(n1148 ,n4559);
    not g3922(n1147 ,n4631);
    not g3923(n1146 ,n4564);
    not g3924(n1145 ,n4577);
    not g3925(n1144 ,n4489);
    not g3926(n1143 ,n7[12]);
    not g3927(n1142 ,n4568);
    not g3928(n1141 ,n4578);
    not g3929(n1140 ,n4602);
    not g3930(n1139 ,n4679);
    not g3931(n1138 ,n4566);
    not g3932(n1137 ,n4672);
    not g3933(n1136 ,n7[10]);
    not g3934(n1135 ,n4610);
    not g3935(n1134 ,n4676);
    not g3936(n1133 ,n4571);
    not g3937(n1132 ,n4593);
    not g3938(n1131 ,n7[15]);
    not g3939(n1130 ,n4605);
    not g3940(n1129 ,n4626);
    not g3941(n1128 ,n4656);
    not g3942(n1127 ,n4654);
    not g3943(n1126 ,n4689);
    not g3944(n1125 ,n4491);
    not g3945(n1124 ,n4635);
    not g3946(n1123 ,n6[2]);
    not g3947(n1122 ,n4642);
    not g3948(n1121 ,n4661);
    not g3949(n1120 ,n4630);
    not g3950(n1119 ,n4693);
    not g3951(n1118 ,n4561);
    not g3952(n1117 ,n4607);
    not g3953(n1116 ,n7[1]);
    not g3954(n1115 ,n4481);
    not g3955(n1114 ,n4663);
    not g3956(n1113 ,n4650);
    not g3957(n1112 ,n7[29]);
    not g3958(n1111 ,n4601);
    not g3959(n1110 ,n7[25]);
    not g3960(n1109 ,n4639);
    not g3961(n1108 ,n4625);
    not g3962(n1107 ,n4556);
    not g3963(n1106 ,n4471);
    not g3964(n1105 ,n4685);
    not g3965(n1104 ,n4640);
    not g3966(n1103 ,n4670);
    not g3967(n1102 ,n4658);
    not g3968(n1101 ,n4573);
    not g3969(n1100 ,n4636);
    not g3970(n1099 ,n4629);
    not g3971(n1098 ,n4647);
    not g3972(n1097 ,n4681);
    not g3973(n1096 ,n4627);
    not g3974(n1095 ,n4598);
    not g3975(n1094 ,n4592);
    not g3976(n1093 ,n4484);
    not g3977(n1092 ,n4584);
    not g3978(n1091 ,n4618);
    not g3979(n1090 ,n7[4]);
    not g3980(n1089 ,n4488);
    not g3981(n1088 ,n4643);
    not g3982(n1087 ,n4466);
    not g3983(n1086 ,n4467);
    not g3984(n1085 ,n4595);
    not g3985(n1084 ,n4472);
    not g3986(n1083 ,n4680);
    not g3987(n1082 ,n4486);
    not g3988(n1081 ,n4644);
    not g3989(n1080 ,n4651);
    not g3990(n1079 ,n4569);
    not g3991(n1078 ,n7[8]);
    not g3992(n1077 ,n4659);
    not g3993(n1076 ,n6[3]);
    not g3994(n1075 ,n4581);
    not g3995(n1074 ,n4473);
    not g3996(n1073 ,n4588);
    not g3997(n1072 ,n4649);
    not g3998(n1071 ,n7[13]);
    not g3999(n1070 ,n4645);
    not g4000(n1069 ,n4665);
    not g4001(n1068 ,n4628);
    not g4002(n1067 ,n4637);
    not g4003(n1066 ,n4482);
    not g4004(n1065 ,n4664);
    not g4005(n1064 ,n4558);
    not g4006(n1063 ,n4623);
    not g4007(n1062 ,n7[24]);
    not g4008(n1061 ,n4600);
    not g4009(n1060 ,n4687);
    not g4010(n1059 ,n4574);
    not g4011(n1058 ,n4622);
    not g4012(n1057 ,n4603);
    not g4013(n1056 ,n4589);
    not g4014(n1055 ,n4565);
    not g4015(n1054 ,n4567);
    not g4016(n1053 ,n7[5]);
    not g4017(n1052 ,n6[1]);
    not g4018(n1051 ,n4669);
    not g4019(n1050 ,n4668);
    not g4020(n1049 ,n4476);
    not g4021(n1048 ,n7[7]);
    not g4022(n1047 ,n4641);
    not g4023(n1046 ,n4594);
    not g4024(n1045 ,n4590);
    not g4025(n1044 ,n4474);
    not g4026(n1043 ,n7[20]);
    not g4027(n1042 ,n4692);
    not g4028(n1041 ,n7[31]);
    not g4029(n1040 ,n4604);
    not g4030(n1039 ,n4621);
    not g4031(n1038 ,n4652);
    not g4032(n1037 ,n4587);
    not g4033(n1036 ,n7[27]);
    not g4034(n1035 ,n4583);
    not g4035(n1034 ,n4613);
    not g4036(n1033 ,n7[19]);
    not g4037(n1032 ,n4469);
    not g4038(n1031 ,n4468);
    not g4039(n1030 ,n4675);
    not g4040(n1029 ,n7[17]);
    not g4041(n1028 ,n4691);
    not g4042(n1027 ,n4586);
    not g4043(n1026 ,n4633);
    not g4044(n1025 ,n4557);
    not g4045(n1024 ,n4576);
    not g4046(n1023 ,n4575);
    not g4047(n1022 ,n4611);
    not g4048(n1021 ,n6[4]);
    not g4049(n1020 ,n4615);
    not g4050(n1019 ,n23[7]);
    not g4051(n1018 ,n4);
    not g4052(n1017 ,n21[17]);
    not g4053(n1016 ,n21[19]);
    not g4054(n1015 ,n10[13]);
    not g4055(n1014 ,n22[4]);
    not g4056(n1013 ,n10[26]);
    not g4057(n1012 ,n21[13]);
    not g4058(n1011 ,n24[9]);
    not g4059(n1010 ,n23[27]);
    not g4060(n1009 ,n23[29]);
    not g4061(n1008 ,n9[29]);
    not g4062(n1007 ,n10[28]);
    not g4063(n1006 ,n23[26]);
    not g4064(n1005 ,n23[18]);
    not g4065(n1004 ,n24[8]);
    not g4066(n1003 ,n36[1]);
    not g4067(n1002 ,n21[2]);
    not g4068(n1001 ,n11[30]);
    not g4069(n1000 ,n24[6]);
    not g4070(n999 ,n11[7]);
    not g4071(n998 ,n22[23]);
    not g4072(n997 ,n22[8]);
    not g4073(n996 ,n10[17]);
    not g4074(n995 ,n24[14]);
    not g4075(n994 ,n24[2]);
    not g4076(n993 ,n9[15]);
    not g4077(n992 ,n21[11]);
    not g4078(n991 ,n22[26]);
    not g4079(n990 ,n9[19]);
    not g4080(n989 ,n11[1]);
    not g4081(n988 ,n10[4]);
    not g4082(n987 ,n23[28]);
    not g4083(n986 ,n24[28]);
    not g4084(n985 ,n21[24]);
    not g4085(n984 ,n21[31]);
    not g4086(n983 ,n24[27]);
    not g4087(n982 ,n22[12]);
    not g4088(n981 ,n22[22]);
    not g4089(n980 ,n9[21]);
    not g4090(n979 ,n9[9]);
    not g4091(n978 ,n2);
    not g4092(n977 ,n23[4]);
    not g4093(n976 ,n10[24]);
    not g4094(n975 ,n3);
    not g4095(n974 ,n11[3]);
    not g4096(n973 ,n23[23]);
    not g4097(n972 ,n22[13]);
    not g4098(n971 ,n11[25]);
    not g4099(n970 ,n23[25]);
    not g4100(n969 ,n11[16]);
    not g4101(n968 ,n21[25]);
    not g4102(n967 ,n24[10]);
    not g4103(n966 ,n27[31]);
    not g4104(n965 ,n25[24]);
    not g4105(n964 ,n27[25]);
    not g4106(n963 ,n28[2]);
    not g4107(n962 ,n27[15]);
    not g4108(n961 ,n25[15]);
    not g4109(n960 ,n27[8]);
    not g4110(n959 ,n26[13]);
    not g4111(n958 ,n25[0]);
    not g4112(n957 ,n28[14]);
    not g4113(n956 ,n26[25]);
    not g4114(n955 ,n26[1]);
    not g4115(n954 ,n27[21]);
    not g4116(n953 ,n34[5]);
    not g4117(n952 ,n27[18]);
    not g4118(n951 ,n35[6]);
    not g4119(n950 ,n25[12]);
    not g4120(n949 ,n34[1]);
    not g4121(n948 ,n28[12]);
    not g4122(n947 ,n26[2]);
    not g4123(n946 ,n28[1]);
    not g4124(n945 ,n26[18]);
    not g4125(n944 ,n25[4]);
    not g4126(n943 ,n35[5]);
    not g4127(n942 ,n28[30]);
    not g4128(n941 ,n25[16]);
    not g4129(n940 ,n26[26]);
    not g4130(n939 ,n28[21]);
    not g4131(n938 ,n27[29]);
    not g4132(n937 ,n25[5]);
    not g4133(n936 ,n25[29]);
    not g4134(n935 ,n29[9]);
    not g4135(n934 ,n31[11]);
    not g4136(n933 ,n8[3]);
    not g4137(n932 ,n8[14]);
    not g4138(n931 ,n8[27]);
    not g4139(n930 ,n8[5]);
    not g4140(n929 ,n31[19]);
    not g4141(n928 ,n29[16]);
    not g4142(n927 ,n8[31]);
    not g4143(n926 ,n32[14]);
    not g4144(n925 ,n31[8]);
    not g4145(n924 ,n29[11]);
    not g4146(n923 ,n8[21]);
    not g4147(n922 ,n8[10]);
    not g4148(n921 ,n30[2]);
    not g4149(n920 ,n31[3]);
    not g4150(n919 ,n8[18]);
    not g4151(n918 ,n30[24]);
    not g4152(n917 ,n29[24]);
    not g4153(n916 ,n29[4]);
    not g4154(n915 ,n8[17]);
    not g4155(n914 ,n8[2]);
    not g4156(n913 ,n30[14]);
    not g4157(n912 ,n8[9]);
    not g4158(n911 ,n8[1]);
    not g4159(n910 ,n8[22]);
    not g4160(n909 ,n31[2]);
    not g4161(n908 ,n32[25]);
    not g4162(n907 ,n8[28]);
    not g4163(n906 ,n8[6]);
    not g4164(n905 ,n8[15]);
    not g4165(n904 ,n8[19]);
    not g4166(n903 ,n32[3]);
    not g4167(n902 ,n32[24]);
    not g4168(n901 ,n29[14]);
    not g4169(n900 ,n30[11]);
    not g4170(n899 ,n30[21]);
    not g4171(n898 ,n8[24]);
    not g4172(n897 ,n32[2]);
    not g4173(n896 ,n8[20]);
    not g4174(n895 ,n8[26]);
    not g4175(n894 ,n31[20]);
    not g4176(n893 ,n8[13]);
    not g4177(n892 ,n32[9]);
    not g4178(n891 ,n8[4]);
    not g4179(n890 ,n29[20]);
    not g4180(n889 ,n8[12]);
    not g4181(n888 ,n34[0]);
    not g4182(n887 ,n31[1]);
    not g4183(n886 ,n30[10]);
    not g4184(n885 ,n8[0]);
    not g4185(n884 ,n29[12]);
    not g4186(n883 ,n8[30]);
    not g4187(n882 ,n31[23]);
    not g4188(n881 ,n8[29]);
    not g4189(n880 ,n30[6]);
    not g4190(n879 ,n8[25]);
    not g4191(n878 ,n8[7]);
    not g4192(n877 ,n8[11]);
    not g4193(n876 ,n8[16]);
    not g4194(n875 ,n8[23]);
    not g4195(n874 ,n31[22]);
    not g4196(n873 ,n8[8]);
    not g4197(n872 ,n33[2]);
    not g4198(n871 ,n37[0]);
    not g4199(n870 ,n6[30]);
    not g4200(n869 ,n6[25]);
    not g4201(n868 ,n6[26]);
    not g4202(n867 ,n6[16]);
    not g4203(n866 ,n6[28]);
    not g4204(n865 ,n6[22]);
    not g4205(n864 ,n6[24]);
    not g4206(n863 ,n6[18]);
    not g4207(n862 ,n6[8]);
    not g4208(n861 ,n6[6]);
    not g4209(n860 ,n6[14]);
    not g4210(n859 ,n6[13]);
    not g4211(n858 ,n6[19]);
    not g4212(n857 ,n6[29]);
    not g4213(n856 ,n6[31]);
    not g4214(n855 ,n6[23]);
    not g4215(n854 ,n6[9]);
    not g4216(n853 ,n6[15]);
    not g4217(n852 ,n6[27]);
    not g4218(n851 ,n6[10]);
    not g4219(n850 ,n6[21]);
    not g4220(n849 ,n6[12]);
    not g4221(n848 ,n6[20]);
    not g4222(n847 ,n6[7]);
    not g4223(n846 ,n6[11]);
    not g4224(n845 ,n6[17]);
    not g4225(n844 ,n6[5]);
    not g4226(n814 ,n843);
    not g4227(n813 ,n843);
    not g4228(n843 ,n4465);
    not g4229(n811 ,n842);
    not g4230(n812 ,n842);
    not g4231(n842 ,n4465);
    not g4232(n841 ,n840);
    not g4233(n839 ,n840);
    not g4234(n810 ,n840);
    not g4235(n799 ,n840);
    not g4236(n840 ,n4465);
    not g4237(n809 ,n822);
    not g4238(n822 ,n1873);
    not g4239(n808 ,n815);
    not g4240(n815 ,n1861);
    not g4241(n807 ,n816);
    not g4242(n816 ,n1862);
    not g4243(n806 ,n821);
    not g4244(n821 ,n1872);
    or g4245(n805 ,n6[5] ,n1798);
    or g4246(n804 ,n844 ,n1798);
    or g4247(n803 ,n844 ,n1766);
    or g4248(n802 ,n814 ,n3565);
    or g4249(n801 ,n3494 ,n3562);
    or g4250(n800 ,n3495 ,n3562);
    xor g4251(n4491 ,n6[31] ,n127);
    xor g4252(n4490 ,n6[30] ,n125);
    nor g4253(n127 ,n41 ,n126);
    nor g4254(n4489 ,n124 ,n125);
    not g4255(n126 ,n125);
    nor g4256(n125 ,n50 ,n123);
    nor g4257(n124 ,n6[29] ,n122);
    xor g4258(n4488 ,n6[28] ,n120);
    not g4259(n123 ,n122);
    nor g4260(n122 ,n46 ,n121);
    nor g4261(n4487 ,n119 ,n120);
    xor g4262(n4486 ,n6[26] ,n118);
    xor g4263(n4484 ,n6[24] ,n117);
    not g4264(n121 ,n120);
    nor g4265(n120 ,n48 ,n116);
    nor g4266(n119 ,n6[27] ,n115);
    nor g4267(n4485 ,n114 ,n118);
    nor g4268(n4483 ,n113 ,n117);
    xor g4269(n4482 ,n6[22] ,n112);
    nor g4270(n118 ,n39 ,n111);
    nor g4271(n117 ,n43 ,n109);
    not g4272(n116 ,n115);
    nor g4273(n115 ,n70 ,n111);
    nor g4274(n114 ,n6[25] ,n110);
    nor g4275(n113 ,n6[23] ,n108);
    nor g4276(n4481 ,n107 ,n112);
    nor g4277(n112 ,n53 ,n106);
    not g4278(n111 ,n110);
    nor g4279(n110 ,n79 ,n106);
    not g4280(n109 ,n108);
    nor g4281(n108 ,n69 ,n106);
    nor g4282(n107 ,n6[21] ,n105);
    xor g4283(n4480 ,n6[20] ,n103);
    not g4284(n106 ,n105);
    nor g4285(n105 ,n59 ,n104);
    nor g4286(n4479 ,n102 ,n103);
    xor g4287(n4478 ,n6[18] ,n101);
    xor g4288(n4476 ,n6[16] ,n100);
    not g4289(n104 ,n103);
    nor g4290(n103 ,n61 ,n99);
    nor g4291(n102 ,n6[19] ,n98);
    nor g4292(n4477 ,n96 ,n101);
    nor g4293(n4475 ,n97 ,n100);
    xor g4294(n4474 ,n6[14] ,n95);
    nor g4295(n101 ,n55 ,n94);
    nor g4296(n100 ,n45 ,n92);
    not g4297(n99 ,n98);
    nor g4298(n98 ,n68 ,n94);
    nor g4299(n97 ,n6[15] ,n91);
    nor g4300(n96 ,n6[17] ,n93);
    nor g4301(n4473 ,n90 ,n95);
    nor g4302(n95 ,n56 ,n89);
    not g4303(n94 ,n93);
    nor g4304(n93 ,n80 ,n89);
    not g4305(n92 ,n91);
    nor g4306(n91 ,n71 ,n89);
    nor g4307(n90 ,n6[13] ,n88);
    xor g4308(n4472 ,n6[12] ,n86);
    not g4309(n89 ,n88);
    nor g4310(n88 ,n44 ,n87);
    nor g4311(n4471 ,n85 ,n86);
    xor g4312(n4470 ,n6[10] ,n84);
    not g4313(n87 ,n86);
    nor g4314(n86 ,n60 ,n83);
    nor g4315(n85 ,n6[11] ,n82);
    nor g4316(n4469 ,n81 ,n84);
    nor g4317(n84 ,n52 ,n78);
    not g4318(n83 ,n82);
    nor g4319(n82 ,n67 ,n78);
    nor g4320(n81 ,n6[9] ,n77);
    xor g4321(n4468 ,n6[8] ,n74);
    or g4322(n80 ,n45 ,n73);
    or g4323(n79 ,n43 ,n76);
    not g4324(n78 ,n77);
    nor g4325(n77 ,n54 ,n75);
    nor g4326(n4467 ,n72 ,n74);
    or g4327(n76 ,n57 ,n69);
    not g4328(n75 ,n74);
    nor g4329(n74 ,n63 ,n66);
    or g4330(n73 ,n47 ,n71);
    nor g4331(n72 ,n6[7] ,n65);
    nor g4332(n4466 ,n65 ,n64);
    or g4333(n71 ,n58 ,n56);
    or g4334(n70 ,n42 ,n39);
    or g4335(n69 ,n38 ,n53);
    or g4336(n68 ,n40 ,n55);
    or g4337(n67 ,n51 ,n52);
    not g4338(n66 ,n65);
    nor g4339(n65 ,n49 ,n62);
    nor g4340(n64 ,n6[6] ,n6[5]);
    not g4341(n63 ,n6[7]);
    not g4342(n62 ,n6[5]);
    not g4343(n61 ,n6[19]);
    not g4344(n60 ,n6[11]);
    not g4345(n59 ,n6[20]);
    not g4346(n58 ,n6[14]);
    not g4347(n57 ,n6[24]);
    not g4348(n56 ,n6[13]);
    not g4349(n55 ,n6[17]);
    not g4350(n54 ,n6[8]);
    not g4351(n53 ,n6[21]);
    not g4352(n52 ,n6[9]);
    not g4353(n51 ,n6[10]);
    not g4354(n50 ,n6[29]);
    not g4355(n49 ,n6[6]);
    not g4356(n48 ,n6[27]);
    not g4357(n47 ,n6[16]);
    not g4358(n46 ,n6[28]);
    not g4359(n45 ,n6[15]);
    not g4360(n44 ,n6[12]);
    not g4361(n43 ,n6[23]);
    not g4362(n42 ,n6[26]);
    not g4363(n41 ,n6[30]);
    not g4364(n40 ,n6[18]);
    not g4365(n39 ,n6[25]);
    not g4366(n38 ,n6[22]);
    xor g4367(n4680 ,n34[7] ,n155);
    nor g4368(n4681 ,n154 ,n155);
    nor g4369(n155 ,n138 ,n153);
    nor g4370(n154 ,n34[6] ,n152);
    nor g4371(n4682 ,n151 ,n152);
    not g4372(n153 ,n152);
    nor g4373(n152 ,n137 ,n150);
    nor g4374(n151 ,n34[5] ,n149);
    nor g4375(n4683 ,n148 ,n149);
    not g4376(n150 ,n149);
    nor g4377(n149 ,n132 ,n147);
    nor g4378(n148 ,n34[4] ,n146);
    nor g4379(n4684 ,n145 ,n146);
    not g4380(n147 ,n146);
    nor g4381(n146 ,n133 ,n144);
    nor g4382(n145 ,n34[3] ,n143);
    nor g4383(n4685 ,n142 ,n143);
    not g4384(n144 ,n143);
    nor g4385(n143 ,n135 ,n141);
    nor g4386(n142 ,n34[2] ,n140);
    nor g4387(n4686 ,n140 ,n139);
    not g4388(n141 ,n140);
    nor g4389(n140 ,n134 ,n136);
    nor g4390(n139 ,n34[1] ,n34[0]);
    not g4391(n138 ,n34[6]);
    not g4392(n137 ,n34[5]);
    not g4393(n136 ,n34[0]);
    not g4394(n135 ,n34[2]);
    not g4395(n134 ,n34[1]);
    not g4396(n133 ,n34[3]);
    not g4397(n132 ,n34[4]);
    xor g4398(n4687 ,n35[7] ,n179);
    nor g4399(n4688 ,n178 ,n179);
    nor g4400(n179 ,n162 ,n177);
    nor g4401(n178 ,n35[6] ,n176);
    nor g4402(n4689 ,n175 ,n176);
    not g4403(n177 ,n176);
    nor g4404(n176 ,n161 ,n174);
    nor g4405(n175 ,n35[5] ,n173);
    nor g4406(n4690 ,n172 ,n173);
    not g4407(n174 ,n173);
    nor g4408(n173 ,n156 ,n171);
    nor g4409(n172 ,n35[4] ,n170);
    nor g4410(n4691 ,n169 ,n170);
    not g4411(n171 ,n170);
    nor g4412(n170 ,n157 ,n168);
    nor g4413(n169 ,n35[3] ,n167);
    nor g4414(n4692 ,n166 ,n167);
    not g4415(n168 ,n167);
    nor g4416(n167 ,n159 ,n165);
    nor g4417(n166 ,n35[2] ,n164);
    nor g4418(n4693 ,n164 ,n163);
    not g4419(n165 ,n164);
    nor g4420(n164 ,n158 ,n160);
    nor g4421(n163 ,n35[1] ,n35[0]);
    not g4422(n162 ,n35[6]);
    not g4423(n161 ,n35[5]);
    not g4424(n160 ,n35[0]);
    not g4425(n159 ,n35[2]);
    not g4426(n158 ,n35[1]);
    not g4427(n157 ,n35[3]);
    not g4428(n156 ,n35[4]);
    xor g4429(n4649 ,n21[31] ,n287);
    nor g4430(n4650 ,n286 ,n287);
    nor g4431(n287 ,n210 ,n285);
    nor g4432(n286 ,n21[30] ,n284);
    xor g4433(n4651 ,n21[29] ,n282);
    not g4434(n285 ,n284);
    nor g4435(n284 ,n197 ,n283);
    nor g4436(n4652 ,n281 ,n282);
    not g4437(n283 ,n282);
    nor g4438(n282 ,n208 ,n280);
    nor g4439(n281 ,n21[28] ,n279);
    xor g4440(n4653 ,n21[27] ,n277);
    not g4441(n280 ,n279);
    nor g4442(n279 ,n183 ,n278);
    nor g4443(n4654 ,n276 ,n277);
    xor g4444(n4655 ,n21[25] ,n275);
    not g4445(n278 ,n277);
    nor g4446(n277 ,n195 ,n274);
    nor g4447(n276 ,n21[26] ,n273);
    nor g4448(n4656 ,n272 ,n275);
    nor g4449(n275 ,n193 ,n271);
    not g4450(n274 ,n273);
    nor g4451(n273 ,n216 ,n271);
    nor g4452(n272 ,n21[24] ,n270);
    xor g4453(n4657 ,n21[23] ,n268);
    not g4454(n271 ,n270);
    nor g4455(n270 ,n182 ,n269);
    nor g4456(n4658 ,n267 ,n268);
    xor g4457(n4659 ,n21[21] ,n266);
    xor g4458(n4661 ,n21[19] ,n265);
    not g4459(n269 ,n268);
    nor g4460(n268 ,n209 ,n264);
    nor g4461(n267 ,n21[22] ,n263);
    nor g4462(n4660 ,n262 ,n266);
    nor g4463(n4662 ,n261 ,n265);
    xor g4464(n4663 ,n21[17] ,n260);
    nor g4465(n266 ,n204 ,n257);
    nor g4466(n265 ,n192 ,n259);
    not g4467(n264 ,n263);
    nor g4468(n263 ,n219 ,n257);
    nor g4469(n262 ,n21[20] ,n256);
    nor g4470(n261 ,n21[18] ,n258);
    nor g4471(n4664 ,n255 ,n260);
    nor g4472(n260 ,n188 ,n254);
    not g4473(n259 ,n258);
    nor g4474(n258 ,n217 ,n254);
    not g4475(n257 ,n256);
    nor g4476(n256 ,n227 ,n254);
    nor g4477(n255 ,n21[16] ,n253);
    xor g4478(n4665 ,n21[15] ,n251);
    not g4479(n254 ,n253);
    nor g4480(n253 ,n203 ,n252);
    nor g4481(n4666 ,n250 ,n251);
    xor g4482(n4667 ,n21[13] ,n249);
    xor g4483(n4669 ,n21[11] ,n248);
    or g4484(n252 ,n186 ,n247);
    nor g4485(n251 ,n203 ,n247);
    nor g4486(n250 ,n21[14] ,n246);
    nor g4487(n4668 ,n244 ,n249);
    nor g4488(n4670 ,n245 ,n248);
    xor g4489(n4671 ,n21[9] ,n243);
    nor g4490(n249 ,n191 ,n242);
    nor g4491(n248 ,n189 ,n240);
    not g4492(n247 ,n246);
    nor g4493(n246 ,n218 ,n242);
    nor g4494(n245 ,n21[10] ,n239);
    nor g4495(n244 ,n21[12] ,n241);
    nor g4496(n4672 ,n238 ,n243);
    nor g4497(n243 ,n198 ,n237);
    not g4498(n242 ,n241);
    nor g4499(n241 ,n228 ,n237);
    not g4500(n240 ,n239);
    nor g4501(n239 ,n215 ,n237);
    nor g4502(n238 ,n21[8] ,n236);
    xor g4503(n4673 ,n21[7] ,n235);
    not g4504(n237 ,n236);
    nor g4505(n236 ,n200 ,n234);
    nor g4506(n4674 ,n233 ,n235);
    xor g4507(n4675 ,n21[5] ,n232);
    nor g4508(n235 ,n200 ,n231);
    or g4509(n234 ,n196 ,n231);
    nor g4510(n233 ,n21[6] ,n230);
    nor g4511(n4676 ,n229 ,n232);
    nor g4512(n232 ,n185 ,n226);
    not g4513(n231 ,n230);
    nor g4514(n230 ,n214 ,n226);
    nor g4515(n229 ,n21[4] ,n225);
    xor g4516(n4677 ,n21[3] ,n223);
    or g4517(n228 ,n189 ,n221);
    or g4518(n227 ,n192 ,n224);
    not g4519(n226 ,n225);
    nor g4520(n225 ,n180 ,n222);
    nor g4521(n4678 ,n220 ,n223);
    or g4522(n224 ,n187 ,n217);
    nor g4523(n223 ,n205 ,n213);
    or g4524(n222 ,n205 ,n213);
    or g4525(n221 ,n184 ,n215);
    nor g4526(n220 ,n21[2] ,n212);
    nor g4527(n4679 ,n212 ,n211);
    or g4528(n219 ,n199 ,n204);
    or g4529(n218 ,n181 ,n191);
    or g4530(n217 ,n206 ,n188);
    or g4531(n216 ,n190 ,n193);
    or g4532(n215 ,n201 ,n198);
    or g4533(n214 ,n202 ,n185);
    not g4534(n213 ,n212);
    nor g4535(n212 ,n194 ,n207);
    nor g4536(n211 ,n21[1] ,n21[0]);
    not g4537(n210 ,n21[30]);
    not g4538(n209 ,n21[22]);
    not g4539(n208 ,n21[28]);
    not g4540(n207 ,n21[0]);
    not g4541(n206 ,n21[17]);
    not g4542(n205 ,n21[2]);
    not g4543(n204 ,n21[20]);
    not g4544(n203 ,n21[14]);
    not g4545(n202 ,n21[5]);
    not g4546(n201 ,n21[9]);
    not g4547(n200 ,n21[6]);
    not g4548(n199 ,n21[21]);
    not g4549(n198 ,n21[8]);
    not g4550(n197 ,n21[29]);
    not g4551(n196 ,n21[7]);
    not g4552(n195 ,n21[26]);
    not g4553(n194 ,n21[1]);
    not g4554(n193 ,n21[24]);
    not g4555(n192 ,n21[18]);
    not g4556(n191 ,n21[12]);
    not g4557(n190 ,n21[25]);
    not g4558(n189 ,n21[10]);
    not g4559(n188 ,n21[16]);
    not g4560(n187 ,n21[19]);
    not g4561(n186 ,n21[15]);
    not g4562(n185 ,n21[4]);
    not g4563(n184 ,n21[11]);
    not g4564(n183 ,n21[27]);
    not g4565(n182 ,n21[23]);
    not g4566(n181 ,n21[13]);
    not g4567(n180 ,n21[3]);
    xor g4568(n4618 ,n22[31] ,n395);
    nor g4569(n4619 ,n394 ,n395);
    nor g4570(n395 ,n318 ,n393);
    nor g4571(n394 ,n22[30] ,n392);
    xor g4572(n4620 ,n22[29] ,n390);
    not g4573(n393 ,n392);
    nor g4574(n392 ,n305 ,n391);
    nor g4575(n4621 ,n389 ,n390);
    not g4576(n391 ,n390);
    nor g4577(n390 ,n316 ,n388);
    nor g4578(n389 ,n22[28] ,n387);
    xor g4579(n4622 ,n22[27] ,n385);
    not g4580(n388 ,n387);
    nor g4581(n387 ,n291 ,n386);
    nor g4582(n4623 ,n384 ,n385);
    xor g4583(n4624 ,n22[25] ,n383);
    not g4584(n386 ,n385);
    nor g4585(n385 ,n303 ,n382);
    nor g4586(n384 ,n22[26] ,n381);
    nor g4587(n4625 ,n380 ,n383);
    nor g4588(n383 ,n301 ,n379);
    not g4589(n382 ,n381);
    nor g4590(n381 ,n324 ,n379);
    nor g4591(n380 ,n22[24] ,n378);
    xor g4592(n4626 ,n22[23] ,n376);
    not g4593(n379 ,n378);
    nor g4594(n378 ,n290 ,n377);
    nor g4595(n4627 ,n375 ,n376);
    xor g4596(n4628 ,n22[21] ,n374);
    xor g4597(n4630 ,n22[19] ,n373);
    not g4598(n377 ,n376);
    nor g4599(n376 ,n317 ,n372);
    nor g4600(n375 ,n22[22] ,n371);
    nor g4601(n4629 ,n370 ,n374);
    nor g4602(n4631 ,n369 ,n373);
    xor g4603(n4632 ,n22[17] ,n368);
    nor g4604(n374 ,n312 ,n365);
    nor g4605(n373 ,n300 ,n367);
    not g4606(n372 ,n371);
    nor g4607(n371 ,n327 ,n365);
    nor g4608(n370 ,n22[20] ,n364);
    nor g4609(n369 ,n22[18] ,n366);
    nor g4610(n4633 ,n363 ,n368);
    nor g4611(n368 ,n296 ,n362);
    not g4612(n367 ,n366);
    nor g4613(n366 ,n325 ,n362);
    not g4614(n365 ,n364);
    nor g4615(n364 ,n335 ,n362);
    nor g4616(n363 ,n22[16] ,n361);
    xor g4617(n4634 ,n22[15] ,n359);
    not g4618(n362 ,n361);
    nor g4619(n361 ,n311 ,n360);
    nor g4620(n4635 ,n358 ,n359);
    xor g4621(n4636 ,n22[13] ,n357);
    xor g4622(n4638 ,n22[11] ,n356);
    or g4623(n360 ,n294 ,n355);
    nor g4624(n359 ,n311 ,n355);
    nor g4625(n358 ,n22[14] ,n354);
    nor g4626(n4637 ,n352 ,n357);
    nor g4627(n4639 ,n353 ,n356);
    xor g4628(n4640 ,n22[9] ,n351);
    nor g4629(n357 ,n299 ,n350);
    nor g4630(n356 ,n297 ,n348);
    not g4631(n355 ,n354);
    nor g4632(n354 ,n326 ,n350);
    nor g4633(n353 ,n22[10] ,n347);
    nor g4634(n352 ,n22[12] ,n349);
    nor g4635(n4641 ,n346 ,n351);
    nor g4636(n351 ,n306 ,n345);
    not g4637(n350 ,n349);
    nor g4638(n349 ,n336 ,n345);
    not g4639(n348 ,n347);
    nor g4640(n347 ,n323 ,n345);
    nor g4641(n346 ,n22[8] ,n344);
    xor g4642(n4642 ,n22[7] ,n343);
    not g4643(n345 ,n344);
    nor g4644(n344 ,n308 ,n342);
    nor g4645(n4643 ,n341 ,n343);
    xor g4646(n4644 ,n22[5] ,n340);
    nor g4647(n343 ,n308 ,n339);
    or g4648(n342 ,n304 ,n339);
    nor g4649(n341 ,n22[6] ,n338);
    nor g4650(n4645 ,n337 ,n340);
    nor g4651(n340 ,n293 ,n334);
    not g4652(n339 ,n338);
    nor g4653(n338 ,n322 ,n334);
    nor g4654(n337 ,n22[4] ,n333);
    xor g4655(n4646 ,n22[3] ,n331);
    or g4656(n336 ,n297 ,n329);
    or g4657(n335 ,n300 ,n332);
    not g4658(n334 ,n333);
    nor g4659(n333 ,n288 ,n330);
    nor g4660(n4647 ,n328 ,n331);
    or g4661(n332 ,n295 ,n325);
    nor g4662(n331 ,n313 ,n321);
    or g4663(n330 ,n313 ,n321);
    or g4664(n329 ,n292 ,n323);
    nor g4665(n328 ,n22[2] ,n320);
    nor g4666(n4648 ,n320 ,n319);
    or g4667(n327 ,n307 ,n312);
    or g4668(n326 ,n289 ,n299);
    or g4669(n325 ,n314 ,n296);
    or g4670(n324 ,n298 ,n301);
    or g4671(n323 ,n309 ,n306);
    or g4672(n322 ,n310 ,n293);
    not g4673(n321 ,n320);
    nor g4674(n320 ,n302 ,n315);
    nor g4675(n319 ,n22[1] ,n22[0]);
    not g4676(n318 ,n22[30]);
    not g4677(n317 ,n22[22]);
    not g4678(n316 ,n22[28]);
    not g4679(n315 ,n22[0]);
    not g4680(n314 ,n22[17]);
    not g4681(n313 ,n22[2]);
    not g4682(n312 ,n22[20]);
    not g4683(n311 ,n22[14]);
    not g4684(n310 ,n22[5]);
    not g4685(n309 ,n22[9]);
    not g4686(n308 ,n22[6]);
    not g4687(n307 ,n22[21]);
    not g4688(n306 ,n22[8]);
    not g4689(n305 ,n22[29]);
    not g4690(n304 ,n22[7]);
    not g4691(n303 ,n22[26]);
    not g4692(n302 ,n22[1]);
    not g4693(n301 ,n22[24]);
    not g4694(n300 ,n22[18]);
    not g4695(n299 ,n22[12]);
    not g4696(n298 ,n22[25]);
    not g4697(n297 ,n22[10]);
    not g4698(n296 ,n22[16]);
    not g4699(n295 ,n22[19]);
    not g4700(n294 ,n22[15]);
    not g4701(n293 ,n22[4]);
    not g4702(n292 ,n22[11]);
    not g4703(n291 ,n22[27]);
    not g4704(n290 ,n22[23]);
    not g4705(n289 ,n22[13]);
    not g4706(n288 ,n22[3]);
    xor g4707(n4587 ,n24[31] ,n503);
    nor g4708(n4588 ,n502 ,n503);
    nor g4709(n503 ,n426 ,n501);
    nor g4710(n502 ,n24[30] ,n500);
    xor g4711(n4589 ,n24[29] ,n498);
    not g4712(n501 ,n500);
    nor g4713(n500 ,n413 ,n499);
    nor g4714(n4590 ,n497 ,n498);
    not g4715(n499 ,n498);
    nor g4716(n498 ,n424 ,n496);
    nor g4717(n497 ,n24[28] ,n495);
    xor g4718(n4591 ,n24[27] ,n493);
    not g4719(n496 ,n495);
    nor g4720(n495 ,n399 ,n494);
    nor g4721(n4592 ,n492 ,n493);
    xor g4722(n4593 ,n24[25] ,n491);
    not g4723(n494 ,n493);
    nor g4724(n493 ,n411 ,n490);
    nor g4725(n492 ,n24[26] ,n489);
    nor g4726(n4594 ,n488 ,n491);
    nor g4727(n491 ,n409 ,n487);
    not g4728(n490 ,n489);
    nor g4729(n489 ,n432 ,n487);
    nor g4730(n488 ,n24[24] ,n486);
    xor g4731(n4595 ,n24[23] ,n484);
    not g4732(n487 ,n486);
    nor g4733(n486 ,n398 ,n485);
    nor g4734(n4596 ,n483 ,n484);
    xor g4735(n4597 ,n24[21] ,n482);
    xor g4736(n4599 ,n24[19] ,n481);
    not g4737(n485 ,n484);
    nor g4738(n484 ,n425 ,n480);
    nor g4739(n483 ,n24[22] ,n479);
    nor g4740(n4598 ,n478 ,n482);
    nor g4741(n4600 ,n477 ,n481);
    xor g4742(n4601 ,n24[17] ,n476);
    nor g4743(n482 ,n420 ,n473);
    nor g4744(n481 ,n408 ,n475);
    not g4745(n480 ,n479);
    nor g4746(n479 ,n435 ,n473);
    nor g4747(n478 ,n24[20] ,n472);
    nor g4748(n477 ,n24[18] ,n474);
    nor g4749(n4602 ,n471 ,n476);
    nor g4750(n476 ,n404 ,n470);
    not g4751(n475 ,n474);
    nor g4752(n474 ,n433 ,n470);
    not g4753(n473 ,n472);
    nor g4754(n472 ,n443 ,n470);
    nor g4755(n471 ,n24[16] ,n469);
    xor g4756(n4603 ,n24[15] ,n467);
    not g4757(n470 ,n469);
    nor g4758(n469 ,n419 ,n468);
    nor g4759(n4604 ,n466 ,n467);
    xor g4760(n4605 ,n24[13] ,n465);
    xor g4761(n4607 ,n24[11] ,n464);
    or g4762(n468 ,n402 ,n463);
    nor g4763(n467 ,n419 ,n463);
    nor g4764(n466 ,n24[14] ,n462);
    nor g4765(n4606 ,n460 ,n465);
    nor g4766(n4608 ,n461 ,n464);
    xor g4767(n4609 ,n24[9] ,n459);
    nor g4768(n465 ,n407 ,n458);
    nor g4769(n464 ,n405 ,n456);
    not g4770(n463 ,n462);
    nor g4771(n462 ,n434 ,n458);
    nor g4772(n461 ,n24[10] ,n455);
    nor g4773(n460 ,n24[12] ,n457);
    nor g4774(n4610 ,n454 ,n459);
    nor g4775(n459 ,n414 ,n453);
    not g4776(n458 ,n457);
    nor g4777(n457 ,n444 ,n453);
    not g4778(n456 ,n455);
    nor g4779(n455 ,n431 ,n453);
    nor g4780(n454 ,n24[8] ,n452);
    xor g4781(n4611 ,n24[7] ,n451);
    not g4782(n453 ,n452);
    nor g4783(n452 ,n416 ,n450);
    nor g4784(n4612 ,n449 ,n451);
    xor g4785(n4613 ,n24[5] ,n448);
    nor g4786(n451 ,n416 ,n447);
    or g4787(n450 ,n412 ,n447);
    nor g4788(n449 ,n24[6] ,n446);
    nor g4789(n4614 ,n445 ,n448);
    nor g4790(n448 ,n401 ,n442);
    not g4791(n447 ,n446);
    nor g4792(n446 ,n430 ,n442);
    nor g4793(n445 ,n24[4] ,n441);
    xor g4794(n4615 ,n24[3] ,n439);
    or g4795(n444 ,n405 ,n437);
    or g4796(n443 ,n408 ,n440);
    not g4797(n442 ,n441);
    nor g4798(n441 ,n396 ,n438);
    nor g4799(n4616 ,n436 ,n439);
    or g4800(n440 ,n403 ,n433);
    nor g4801(n439 ,n421 ,n429);
    or g4802(n438 ,n421 ,n429);
    or g4803(n437 ,n400 ,n431);
    nor g4804(n436 ,n24[2] ,n428);
    nor g4805(n4617 ,n428 ,n427);
    or g4806(n435 ,n415 ,n420);
    or g4807(n434 ,n397 ,n407);
    or g4808(n433 ,n422 ,n404);
    or g4809(n432 ,n406 ,n409);
    or g4810(n431 ,n417 ,n414);
    or g4811(n430 ,n418 ,n401);
    not g4812(n429 ,n428);
    nor g4813(n428 ,n410 ,n423);
    nor g4814(n427 ,n24[1] ,n24[0]);
    not g4815(n426 ,n24[30]);
    not g4816(n425 ,n24[22]);
    not g4817(n424 ,n24[28]);
    not g4818(n423 ,n24[0]);
    not g4819(n422 ,n24[17]);
    not g4820(n421 ,n24[2]);
    not g4821(n420 ,n24[20]);
    not g4822(n419 ,n24[14]);
    not g4823(n418 ,n24[5]);
    not g4824(n417 ,n24[9]);
    not g4825(n416 ,n24[6]);
    not g4826(n415 ,n24[21]);
    not g4827(n414 ,n24[8]);
    not g4828(n413 ,n24[29]);
    not g4829(n412 ,n24[7]);
    not g4830(n411 ,n24[26]);
    not g4831(n410 ,n24[1]);
    not g4832(n409 ,n24[24]);
    not g4833(n408 ,n24[18]);
    not g4834(n407 ,n24[12]);
    not g4835(n406 ,n24[25]);
    not g4836(n405 ,n24[10]);
    not g4837(n404 ,n24[16]);
    not g4838(n403 ,n24[19]);
    not g4839(n402 ,n24[15]);
    not g4840(n401 ,n24[4]);
    not g4841(n400 ,n24[11]);
    not g4842(n399 ,n24[27]);
    not g4843(n398 ,n24[23]);
    not g4844(n397 ,n24[13]);
    not g4845(n396 ,n24[3]);
    xor g4846(n4556 ,n23[31] ,n611);
    nor g4847(n4557 ,n610 ,n611);
    nor g4848(n611 ,n534 ,n609);
    nor g4849(n610 ,n23[30] ,n608);
    xor g4850(n4558 ,n23[29] ,n606);
    not g4851(n609 ,n608);
    nor g4852(n608 ,n521 ,n607);
    nor g4853(n4559 ,n605 ,n606);
    not g4854(n607 ,n606);
    nor g4855(n606 ,n532 ,n604);
    nor g4856(n605 ,n23[28] ,n603);
    xor g4857(n4560 ,n23[27] ,n601);
    not g4858(n604 ,n603);
    nor g4859(n603 ,n507 ,n602);
    nor g4860(n4561 ,n600 ,n601);
    xor g4861(n4562 ,n23[25] ,n599);
    not g4862(n602 ,n601);
    nor g4863(n601 ,n519 ,n598);
    nor g4864(n600 ,n23[26] ,n597);
    nor g4865(n4563 ,n596 ,n599);
    nor g4866(n599 ,n517 ,n595);
    not g4867(n598 ,n597);
    nor g4868(n597 ,n540 ,n595);
    nor g4869(n596 ,n23[24] ,n594);
    xor g4870(n4564 ,n23[23] ,n592);
    not g4871(n595 ,n594);
    nor g4872(n594 ,n506 ,n593);
    nor g4873(n4565 ,n591 ,n592);
    xor g4874(n4566 ,n23[21] ,n590);
    xor g4875(n4568 ,n23[19] ,n589);
    not g4876(n593 ,n592);
    nor g4877(n592 ,n533 ,n588);
    nor g4878(n591 ,n23[22] ,n587);
    nor g4879(n4567 ,n586 ,n590);
    nor g4880(n4569 ,n585 ,n589);
    xor g4881(n4570 ,n23[17] ,n584);
    nor g4882(n590 ,n528 ,n581);
    nor g4883(n589 ,n516 ,n583);
    not g4884(n588 ,n587);
    nor g4885(n587 ,n543 ,n581);
    nor g4886(n586 ,n23[20] ,n580);
    nor g4887(n585 ,n23[18] ,n582);
    nor g4888(n4571 ,n579 ,n584);
    nor g4889(n584 ,n512 ,n578);
    not g4890(n583 ,n582);
    nor g4891(n582 ,n541 ,n578);
    not g4892(n581 ,n580);
    nor g4893(n580 ,n551 ,n578);
    nor g4894(n579 ,n23[16] ,n577);
    xor g4895(n4572 ,n23[15] ,n575);
    not g4896(n578 ,n577);
    nor g4897(n577 ,n527 ,n576);
    nor g4898(n4573 ,n574 ,n575);
    xor g4899(n4574 ,n23[13] ,n573);
    xor g4900(n4576 ,n23[11] ,n572);
    or g4901(n576 ,n510 ,n571);
    nor g4902(n575 ,n527 ,n571);
    nor g4903(n574 ,n23[14] ,n570);
    nor g4904(n4575 ,n568 ,n573);
    nor g4905(n4577 ,n569 ,n572);
    xor g4906(n4578 ,n23[9] ,n567);
    nor g4907(n573 ,n515 ,n566);
    nor g4908(n572 ,n513 ,n564);
    not g4909(n571 ,n570);
    nor g4910(n570 ,n542 ,n566);
    nor g4911(n569 ,n23[10] ,n563);
    nor g4912(n568 ,n23[12] ,n565);
    nor g4913(n4579 ,n562 ,n567);
    nor g4914(n567 ,n522 ,n561);
    not g4915(n566 ,n565);
    nor g4916(n565 ,n552 ,n561);
    not g4917(n564 ,n563);
    nor g4918(n563 ,n539 ,n561);
    nor g4919(n562 ,n23[8] ,n560);
    xor g4920(n4580 ,n23[7] ,n559);
    not g4921(n561 ,n560);
    nor g4922(n560 ,n524 ,n558);
    nor g4923(n4581 ,n557 ,n559);
    xor g4924(n4582 ,n23[5] ,n556);
    nor g4925(n559 ,n524 ,n555);
    or g4926(n558 ,n520 ,n555);
    nor g4927(n557 ,n23[6] ,n554);
    nor g4928(n4583 ,n553 ,n556);
    nor g4929(n556 ,n509 ,n550);
    not g4930(n555 ,n554);
    nor g4931(n554 ,n538 ,n550);
    nor g4932(n553 ,n23[4] ,n549);
    xor g4933(n4584 ,n23[3] ,n547);
    or g4934(n552 ,n513 ,n545);
    or g4935(n551 ,n516 ,n548);
    not g4936(n550 ,n549);
    nor g4937(n549 ,n504 ,n546);
    nor g4938(n4585 ,n544 ,n547);
    or g4939(n548 ,n511 ,n541);
    nor g4940(n547 ,n529 ,n537);
    or g4941(n546 ,n529 ,n537);
    or g4942(n545 ,n508 ,n539);
    nor g4943(n544 ,n23[2] ,n536);
    nor g4944(n4586 ,n536 ,n535);
    or g4945(n543 ,n523 ,n528);
    or g4946(n542 ,n505 ,n515);
    or g4947(n541 ,n530 ,n512);
    or g4948(n540 ,n514 ,n517);
    or g4949(n539 ,n525 ,n522);
    or g4950(n538 ,n526 ,n509);
    not g4951(n537 ,n536);
    nor g4952(n536 ,n518 ,n531);
    nor g4953(n535 ,n23[1] ,n23[0]);
    not g4954(n534 ,n23[30]);
    not g4955(n533 ,n23[22]);
    not g4956(n532 ,n23[28]);
    not g4957(n531 ,n23[0]);
    not g4958(n530 ,n23[17]);
    not g4959(n529 ,n23[2]);
    not g4960(n528 ,n23[20]);
    not g4961(n527 ,n23[14]);
    not g4962(n526 ,n23[5]);
    not g4963(n525 ,n23[9]);
    not g4964(n524 ,n23[6]);
    not g4965(n523 ,n23[21]);
    not g4966(n522 ,n23[8]);
    not g4967(n521 ,n23[29]);
    not g4968(n520 ,n23[7]);
    not g4969(n519 ,n23[26]);
    not g4970(n518 ,n23[1]);
    not g4971(n517 ,n23[24]);
    not g4972(n516 ,n23[18]);
    not g4973(n515 ,n23[12]);
    not g4974(n514 ,n23[25]);
    not g4975(n513 ,n23[10]);
    not g4976(n512 ,n23[16]);
    not g4977(n511 ,n23[19]);
    not g4978(n510 ,n23[15]);
    not g4979(n509 ,n23[4]);
    not g4980(n508 ,n23[11]);
    not g4981(n507 ,n23[27]);
    not g4982(n506 ,n23[23]);
    not g4983(n505 ,n23[13]);
    not g4984(n504 ,n23[3]);
    nor g4985(n37[0] ,n703 ,n798);
    nor g4986(n798 ,n743 ,n797);
    nor g4987(n797 ,n746 ,n796);
    nor g4988(n796 ,n768 ,n795);
    nor g4989(n795 ,n748 ,n794);
    nor g4990(n794 ,n739 ,n793);
    nor g4991(n793 ,n763 ,n792);
    nor g4992(n792 ,n755 ,n791);
    nor g4993(n791 ,n750 ,n790);
    nor g4994(n790 ,n745 ,n789);
    nor g4995(n789 ,n741 ,n788);
    nor g4996(n788 ,n761 ,n787);
    nor g4997(n787 ,n765 ,n786);
    nor g4998(n786 ,n760 ,n785);
    nor g4999(n785 ,n757 ,n784);
    nor g5000(n784 ,n738 ,n783);
    nor g5001(n783 ,n749 ,n782);
    nor g5002(n782 ,n747 ,n781);
    nor g5003(n781 ,n744 ,n780);
    nor g5004(n780 ,n742 ,n779);
    nor g5005(n779 ,n740 ,n778);
    nor g5006(n778 ,n753 ,n777);
    nor g5007(n777 ,n767 ,n776);
    nor g5008(n776 ,n766 ,n775);
    nor g5009(n775 ,n764 ,n774);
    nor g5010(n774 ,n762 ,n773);
    nor g5011(n773 ,n759 ,n772);
    nor g5012(n772 ,n758 ,n771);
    nor g5013(n771 ,n756 ,n770);
    nor g5014(n770 ,n754 ,n769);
    nor g5015(n769 ,n752 ,n751);
    or g5016(n768 ,n716 ,n708);
    or g5017(n767 ,n734 ,n732);
    or g5018(n766 ,n729 ,n728);
    or g5019(n765 ,n723 ,n707);
    or g5020(n764 ,n724 ,n722);
    or g5021(n763 ,n720 ,n714);
    or g5022(n762 ,n719 ,n717);
    or g5023(n761 ,n733 ,n730);
    or g5024(n760 ,n713 ,n712);
    or g5025(n759 ,n725 ,n721);
    or g5026(n758 ,n710 ,n709);
    or g5027(n757 ,n690 ,n684);
    or g5028(n756 ,n735 ,n691);
    or g5029(n755 ,n705 ,n701);
    or g5030(n754 ,n731 ,n704);
    or g5031(n753 ,n675 ,n737);
    nor g5032(n752 ,n706 ,n699);
    or g5033(n751 ,n697 ,n702);
    or g5034(n750 ,n695 ,n692);
    or g5035(n749 ,n696 ,n694);
    or g5036(n748 ,n693 ,n715);
    or g5037(n747 ,n711 ,n689);
    or g5038(n746 ,n688 ,n727);
    or g5039(n745 ,n686 ,n685);
    or g5040(n744 ,n687 ,n718);
    or g5041(n743 ,n681 ,n726);
    or g5042(n742 ,n683 ,n682);
    or g5043(n741 ,n679 ,n676);
    or g5044(n740 ,n680 ,n678);
    or g5045(n739 ,n677 ,n736);
    or g5046(n738 ,n700 ,n698);
    nor g5047(n737 ,n613 ,n4534);
    nor g5048(n736 ,n632 ,n4550);
    nor g5049(n735 ,n673 ,n4496);
    nor g5050(n734 ,n634 ,n4502);
    nor g5051(n733 ,n627 ,n4545);
    nor g5052(n732 ,n669 ,n4501);
    nor g5053(n731 ,n618 ,n4527);
    nor g5054(n730 ,n661 ,n4544);
    nor g5055(n729 ,n646 ,n4533);
    nor g5056(n728 ,n654 ,n4532);
    nor g5057(n727 ,n640 ,n4521);
    nor g5058(n726 ,n636 ,n4554);
    nor g5059(n725 ,n668 ,n4498);
    nor g5060(n724 ,n652 ,n4500);
    nor g5061(n723 ,n629 ,n4512);
    nor g5062(n722 ,n612 ,n4499);
    nor g5063(n721 ,n660 ,n4497);
    nor g5064(n720 ,n659 ,n4518);
    nor g5065(n719 ,n649 ,n4531);
    nor g5066(n718 ,n648 ,n4505);
    nor g5067(n717 ,n656 ,n4530);
    nor g5068(n716 ,n666 ,n4553);
    nor g5069(n715 ,n619 ,n4519);
    nor g5070(n714 ,n638 ,n4517);
    nor g5071(n713 ,n658 ,n4543);
    nor g5072(n712 ,n622 ,n4542);
    nor g5073(n711 ,n631 ,n4539);
    nor g5074(n710 ,n642 ,n4529);
    nor g5075(n709 ,n662 ,n4528);
    nor g5076(n708 ,n639 ,n4552);
    nor g5077(n707 ,n635 ,n4511);
    nor g5078(n706 ,n667 ,n4525);
    nor g5079(n705 ,n617 ,n4549);
    nor g5080(n704 ,n615 ,n4526);
    nor g5081(n703 ,n655 ,n4523);
    nor g5082(n702 ,n643 ,n4493);
    nor g5083(n701 ,n653 ,n4548);
    nor g5084(n700 ,n623 ,n4541);
    nor g5085(n699 ,n674 ,n4524);
    nor g5086(n698 ,n663 ,n4540);
    nor g5087(n697 ,n633 ,n4494);
    nor g5088(n696 ,n621 ,n4508);
    nor g5089(n695 ,n664 ,n4516);
    nor g5090(n694 ,n620 ,n4507);
    nor g5091(n693 ,n641 ,n4520);
    nor g5092(n692 ,n651 ,n4515);
    nor g5093(n691 ,n665 ,n4495);
    nor g5094(n690 ,n637 ,n4510);
    nor g5095(n689 ,n650 ,n4538);
    nor g5096(n688 ,n671 ,n4522);
    nor g5097(n687 ,n614 ,n4506);
    nor g5098(n686 ,n630 ,n4547);
    nor g5099(n685 ,n628 ,n4546);
    nor g5100(n684 ,n657 ,n4509);
    nor g5101(n683 ,n616 ,n4537);
    nor g5102(n682 ,n670 ,n4536);
    nor g5103(n681 ,n626 ,n4555);
    nor g5104(n680 ,n645 ,n4504);
    nor g5105(n679 ,n624 ,n4514);
    nor g5106(n678 ,n644 ,n4503);
    nor g5107(n677 ,n647 ,n4551);
    nor g5108(n676 ,n625 ,n4513);
    nor g5109(n675 ,n672 ,n4535);
    not g5110(n674 ,n4492);
    not g5111(n673 ,n4528);
    not g5112(n672 ,n4503);
    not g5113(n671 ,n4554);
    not g5114(n670 ,n4504);
    not g5115(n669 ,n4533);
    not g5116(n668 ,n4530);
    not g5117(n667 ,n4493);
    not g5118(n666 ,n4521);
    not g5119(n665 ,n4527);
    not g5120(n664 ,n4548);
    not g5121(n663 ,n4508);
    not g5122(n662 ,n4496);
    not g5123(n661 ,n4512);
    not g5124(n660 ,n4529);
    not g5125(n659 ,n4550);
    not g5126(n658 ,n4511);
    not g5127(n657 ,n4541);
    not g5128(n656 ,n4498);
    not g5129(n655 ,n4555);
    not g5130(n654 ,n4500);
    not g5131(n653 ,n4516);
    not g5132(n652 ,n4532);
    not g5133(n651 ,n4547);
    not g5134(n650 ,n4506);
    not g5135(n649 ,n4499);
    not g5136(n648 ,n4537);
    not g5137(n647 ,n4519);
    not g5138(n646 ,n4501);
    not g5139(n645 ,n4536);
    not g5140(n644 ,n4535);
    not g5141(n643 ,n4525);
    not g5142(n642 ,n4497);
    not g5143(n641 ,n4552);
    not g5144(n640 ,n4553);
    not g5145(n639 ,n4520);
    not g5146(n638 ,n4549);
    not g5147(n637 ,n4542);
    not g5148(n636 ,n4522);
    not g5149(n635 ,n4543);
    not g5150(n634 ,n4534);
    not g5151(n633 ,n4526);
    not g5152(n632 ,n4518);
    not g5153(n631 ,n4507);
    not g5154(n630 ,n4515);
    not g5155(n629 ,n4544);
    not g5156(n628 ,n4514);
    not g5157(n627 ,n4513);
    not g5158(n626 ,n4523);
    not g5159(n625 ,n4545);
    not g5160(n624 ,n4546);
    not g5161(n623 ,n4509);
    not g5162(n622 ,n4510);
    not g5163(n621 ,n4540);
    not g5164(n620 ,n4539);
    not g5165(n619 ,n4551);
    not g5166(n618 ,n4495);
    not g5167(n617 ,n4517);
    not g5168(n616 ,n4505);
    not g5169(n615 ,n4494);
    not g5170(n614 ,n4538);
    not g5171(n613 ,n4502);
    not g5172(n612 ,n4531);
endmodule
