module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n11);
    input [63:0] n0;
    input [31:0] n1;
    input [3:0] n2;
    input n3;
    input [1:0] n4;
    input [5:0] n5;
    output [63:0] n6;
    output [31:0] n7;
    output n8, n9, n10, n11;
    output [5:0] n12;
    output [7:0] n13;
    wire [63:0] n0;
    wire [31:0] n1;
    wire [3:0] n2;
    wire n3;
    wire [1:0] n4;
    wire [5:0] n5;
    wire [63:0] n6;
    wire [31:0] n7;
    wire n8, n9, n10, n11;
    wire [5:0] n12;
    wire [7:0] n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133;
    wire n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
    wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
    wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157;
    wire n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165;
    wire n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
    wire n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
    wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
    wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
    wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
    wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
    wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
    wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
    wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
    wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
    wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
    wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
    wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
    wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277;
    wire n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285;
    wire n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293;
    wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
    wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
    wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
    wire n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325;
    wire n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333;
    wire n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
    wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
    wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357;
    wire n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365;
    wire n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373;
    wire n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
    wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
    wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397;
    wire n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405;
    wire n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413;
    wire n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
    wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
    wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437;
    wire n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
    wire n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453;
    wire n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
    wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
    wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477;
    wire n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485;
    wire n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493;
    wire n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
    wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
    wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
    wire n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;
    wire n2526, n2527;
    buf g0(n13[4], 1'b0);
    buf g1(n13[5], 1'b0);
    buf g2(n13[6], 1'b0);
    buf g3(n13[7], 1'b0);
    buf g4(n12[0], 1'b0);
    buf g5(n12[1], 1'b0);
    buf g6(n12[2], 1'b0);
    not g7(n2374 ,n2425);
    not g8(n2373 ,n2411);
    not g9(n2372 ,n2396);
    not g10(n2371 ,n2397);
    not g11(n2370 ,n2410);
    or g12(n10 ,n2494 ,n2368);
    or g13(n8 ,n2377 ,n2369);
    nor g14(n2369 ,n2367 ,n2364);
    nor g15(n2368 ,n2366 ,n2365);
    or g16(n2367 ,n2363 ,n2428);
    or g17(n2366 ,n2362 ,n3);
    or g18(n2364 ,n2493 ,n2376);
    not g19(n2363 ,n2426);
    not g20(n2362 ,n2428);
    nor g21(n2410 ,n2348 ,n2361);
    nor g22(n2396 ,n2346 ,n2360);
    nor g23(n2397 ,n2339 ,n2358);
    nor g24(n2411 ,n2340 ,n2359);
    or g25(n2361 ,n2321 ,n2356);
    or g26(n2360 ,n2328 ,n2355);
    or g27(n2359 ,n2312 ,n2354);
    or g28(n2358 ,n2306 ,n2357);
    or g29(n2357 ,n2334 ,n2353);
    or g30(n2356 ,n2325 ,n2351);
    or g31(n2355 ,n2326 ,n2352);
    or g32(n2354 ,n2309 ,n2350);
    or g33(n2353 ,n2345 ,n2344);
    or g34(n2352 ,n2343 ,n2342);
    or g35(n2351 ,n2341 ,n2347);
    or g36(n2350 ,n2338 ,n2349);
    or g37(n2349 ,n2336 ,n2335);
    or g38(n2348 ,n2330 ,n2308);
    or g39(n2347 ,n2329 ,n2313);
    or g40(n2346 ,n2333 ,n2331);
    or g41(n2345 ,n2332 ,n2327);
    or g42(n2344 ,n2323 ,n2319);
    or g43(n2343 ,n2324 ,n2337);
    or g44(n2342 ,n2318 ,n2317);
    or g45(n2341 ,n2311 ,n2322);
    or g46(n2340 ,n2316 ,n2314);
    or g47(n2339 ,n2315 ,n2310);
    or g48(n2338 ,n2307 ,n2320);
    xor g49(n2337 ,n0[30] ,n1[30]);
    xor g50(n2336 ,n0[9] ,n1[9]);
    xor g51(n2335 ,n0[8] ,n1[8]);
    xor g52(n2334 ,n0[22] ,n1[22]);
    xor g53(n2333 ,n0[27] ,n1[27]);
    xor g54(n2332 ,n0[19] ,n1[19]);
    xor g55(n2331 ,n0[26] ,n1[26]);
    xor g56(n2330 ,n0[2] ,n1[2]);
    xor g57(n2329 ,n0[5] ,n1[5]);
    xor g58(n2328 ,n0[24] ,n1[24]);
    xor g59(n2327 ,n0[18] ,n1[18]);
    xor g60(n2326 ,n0[25] ,n1[25]);
    xor g61(n2325 ,n0[3] ,n1[3]);
    xor g62(n2324 ,n0[31] ,n1[31]);
    xor g63(n2323 ,n0[17] ,n1[17]);
    xor g64(n2322 ,n0[6] ,n1[6]);
    not g65(n2321 ,n2425);
    xor g66(n2320 ,n0[10] ,n1[10]);
    xor g67(n2319 ,n0[16] ,n1[16]);
    xor g68(n2318 ,n0[29] ,n1[29]);
    xor g69(n2317 ,n0[28] ,n1[28]);
    xor g70(n2316 ,n0[14] ,n1[14]);
    xor g71(n2315 ,n0[23] ,n1[23]);
    xor g72(n2314 ,n0[13] ,n1[13]);
    xor g73(n2313 ,n0[4] ,n1[4]);
    xor g74(n2312 ,n0[15] ,n1[15]);
    xor g75(n2311 ,n0[7] ,n1[7]);
    xor g76(n2310 ,n0[21] ,n1[21]);
    xor g77(n2309 ,n0[12] ,n1[12]);
    xor g78(n2308 ,n0[1] ,n1[1]);
    xor g79(n2307 ,n0[11] ,n1[11]);
    xor g80(n2306 ,n0[20] ,n1[20]);
    xnor g81(n2425 ,n0[0] ,n1[0]);
    nor g82(n2424 ,n2305 ,n2304);
    or g83(n2423 ,n2304 ,n4[1]);
    not g84(n2305 ,n4[1]);
    not g85(n2304 ,n4[0]);
    not g86(n2444 ,n0[48]);
    not g87(n2429 ,n0[63]);
    not g88(n2430 ,n0[62]);
    not g89(n2431 ,n0[61]);
    not g90(n2432 ,n0[60]);
    not g91(n2433 ,n0[59]);
    not g92(n2434 ,n0[58]);
    not g93(n2435 ,n0[57]);
    not g94(n2436 ,n0[56]);
    not g95(n2437 ,n0[55]);
    not g96(n2438 ,n0[54]);
    not g97(n2439 ,n0[53]);
    not g98(n2440 ,n0[52]);
    not g99(n2441 ,n0[51]);
    not g100(n2442 ,n0[50]);
    not g101(n2443 ,n0[49]);
    not g102(n2492 ,n0[0]);
    not g103(n2445 ,n0[47]);
    not g104(n2446 ,n0[46]);
    not g105(n2447 ,n0[45]);
    not g106(n2448 ,n0[44]);
    not g107(n2449 ,n0[43]);
    not g108(n2450 ,n0[42]);
    not g109(n2451 ,n0[41]);
    not g110(n2452 ,n0[40]);
    not g111(n2453 ,n0[39]);
    not g112(n2454 ,n0[38]);
    not g113(n2455 ,n0[37]);
    not g114(n2456 ,n0[36]);
    not g115(n2457 ,n0[35]);
    not g116(n2458 ,n0[34]);
    not g117(n2459 ,n0[33]);
    not g118(n2476 ,n0[16]);
    not g119(n2461 ,n0[31]);
    not g120(n2462 ,n0[30]);
    not g121(n2463 ,n0[29]);
    not g122(n2464 ,n0[28]);
    not g123(n2465 ,n0[27]);
    not g124(n2466 ,n0[26]);
    not g125(n2467 ,n0[25]);
    not g126(n2468 ,n0[24]);
    not g127(n2469 ,n0[23]);
    not g128(n2470 ,n0[22]);
    not g129(n2471 ,n0[21]);
    not g130(n2472 ,n0[20]);
    not g131(n2473 ,n0[19]);
    not g132(n2474 ,n0[18]);
    not g133(n2475 ,n0[17]);
    not g134(n2460 ,n0[32]);
    not g135(n2477 ,n0[15]);
    not g136(n2478 ,n0[14]);
    not g137(n2479 ,n0[13]);
    not g138(n2480 ,n0[12]);
    not g139(n2481 ,n0[11]);
    not g140(n2482 ,n0[10]);
    not g141(n2483 ,n0[9]);
    not g142(n2484 ,n0[8]);
    not g143(n2485 ,n0[7]);
    not g144(n2486 ,n0[6]);
    not g145(n2487 ,n0[5]);
    not g146(n2488 ,n0[4]);
    not g147(n2489 ,n0[3]);
    not g148(n2490 ,n0[2]);
    not g149(n2491 ,n0[1]);
    or g150(n9 ,n2498 ,n2303);
    nor g151(n2303 ,n3 ,n2302);
    or g152(n2302 ,n2375 ,n2426);
    or g153(n13[2] ,n2496 ,n2300);
    or g154(n2426 ,n2301 ,n2297);
    or g155(n13[1] ,n2497 ,n2299);
    or g156(n13[0] ,n2495 ,n2298);
    or g157(n2301 ,n2295 ,n2414);
    nor g158(n2300 ,n2293 ,n2376);
    nor g159(n2299 ,n2295 ,n2376);
    nor g160(n2298 ,n2296 ,n2376);
    nor g161(n13[3] ,n2294 ,n2376);
    not g162(n2296 ,n2414);
    not g163(n2295 ,n2413);
    not g164(n2294 ,n2412);
    not g165(n2293 ,n2398);
    nor g166(n2377 ,n3 ,n2292);
    or g167(n2292 ,n2290 ,n2291);
    nor g168(n2291 ,n2274 ,n2289);
    nor g169(n2290 ,n2022 ,n2287);
    or g170(n12[3] ,n1824 ,n2288);
    or g171(n2289 ,n2285 ,n2286);
    nor g172(n2288 ,n2376 ,n2280);
    or g173(n2287 ,n2242 ,n2281);
    nor g174(n2286 ,n1355 ,n2283);
    nor g175(n2285 ,n1351 ,n2284);
    or g176(n12[4] ,n1825 ,n2282);
    nor g177(n2284 ,n2205 ,n2278);
    nor g178(n2283 ,n2258 ,n2275);
    nor g179(n2493 ,n2206 ,n2279);
    nor g180(n2282 ,n2376 ,n2276);
    nor g181(n2281 ,n1351 ,n2277);
    nor g182(n2280 ,n2399 ,n2273);
    or g183(n2279 ,n2223 ,n2272);
    or g184(n2278 ,n2249 ,n2270);
    nor g185(n2277 ,n2132 ,n2269);
    nor g186(n2276 ,n2221 ,n2265);
    or g187(n2275 ,n2154 ,n2268);
    or g188(n2274 ,n2264 ,n2266);
    nor g189(n12[5] ,n2376 ,n2271);
    nor g190(n2273 ,n2401 ,n2267);
    not g191(n2272 ,n2271);
    or g192(n2270 ,n2224 ,n2257);
    or g193(n2269 ,n2131 ,n2263);
    or g194(n2268 ,n2162 ,n2256);
    nor g195(n2271 ,n2221 ,n2261);
    nor g196(n2267 ,n2402 ,n2260);
    nor g197(n2266 ,n1352 ,n2262);
    nor g198(n2265 ,n2222 ,n2261);
    or g199(n2264 ,n2[0] ,n2259);
    or g200(n2263 ,n2199 ,n2252);
    nor g201(n2262 ,n2117 ,n2250);
    or g202(n7[3] ,n2000 ,n2255);
    or g203(n7[2] ,n1999 ,n2254);
    or g204(n7[1] ,n1998 ,n2253);
    or g205(n7[6] ,n1997 ,n2248);
    nor g206(n2260 ,n2403 ,n2243);
    nor g207(n2259 ,n1356 ,n2251);
    or g208(n2258 ,n2246 ,n2155);
    or g209(n2257 ,n2153 ,n2247);
    or g210(n2256 ,n2146 ,n2245);
    or g211(n7[4] ,n2207 ,n2244);
    or g212(n2261 ,n2402 ,n2403);
    or g213(n7[11] ,n2063 ,n2241);
    or g214(n2255 ,n2238 ,n2180);
    or g215(n2254 ,n2237 ,n2179);
    or g216(n2253 ,n2236 ,n2176);
    or g217(n2252 ,n2233 ,n2231);
    or g218(n7[12] ,n2064 ,n2234);
    nor g219(n2251 ,n1793 ,n2230);
    or g220(n2250 ,n2018 ,n2228);
    or g221(n2249 ,n2226 ,n2225);
    or g222(n2248 ,n2214 ,n2156);
    or g223(n2247 ,n2211 ,n2219);
    or g224(n2246 ,n1424 ,n2217);
    or g225(n2245 ,n2216 ,n2215);
    or g226(n7[5] ,n2098 ,n2232);
    or g227(n2244 ,n2091 ,n2239);
    or g228(n7[0] ,n2094 ,n2235);
    or g229(n7[15] ,n2012 ,n2240);
    or g230(n7[14] ,n2087 ,n2213);
    or g231(n7[13] ,n2083 ,n2212);
    or g232(n7[9] ,n2005 ,n2229);
    or g233(n7[8] ,n2075 ,n2208);
    or g234(n7[10] ,n2006 ,n2227);
    or g235(n7[7] ,n2003 ,n2218);
    nor g236(n2243 ,n2404 ,n2220);
    or g237(n2242 ,n2210 ,n2209);
    xnor g238(n2403 ,n1[4] ,n2177);
    or g239(n2241 ,n1987 ,n2174);
    or g240(n2240 ,n2108 ,n2181);
    or g241(n2239 ,n2069 ,n2203);
    or g242(n2238 ,n1809 ,n2188);
    or g243(n2237 ,n1806 ,n2187);
    or g244(n2236 ,n1804 ,n2186);
    or g245(n2235 ,n2202 ,n2103);
    or g246(n2234 ,n1989 ,n2175);
    or g247(n2233 ,n2198 ,n2197);
    or g248(n2232 ,n2204 ,n2136);
    or g249(n2231 ,n2196 ,n2195);
    or g250(n2230 ,n2194 ,n2193);
    or g251(n2229 ,n2116 ,n2172);
    or g252(n2228 ,n2017 ,n2192);
    or g253(n2227 ,n2118 ,n2173);
    or g254(n2226 ,n2171 ,n2170);
    or g255(n2225 ,n2169 ,n2168);
    or g256(n2224 ,n2167 ,n2191);
    not g257(n2223 ,n2222);
    nor g258(n2220 ,n2178 ,n2405);
    or g259(n2219 ,n2164 ,n2163);
    or g260(n2218 ,n2189 ,n2157);
    or g261(n2217 ,n1422 ,n2183);
    or g262(n2216 ,n2161 ,n2160);
    or g263(n2215 ,n2159 ,n2158);
    or g264(n2214 ,n1771 ,n2182);
    or g265(n2213 ,n2084 ,n2185);
    or g266(n2212 ,n2010 ,n2184);
    or g267(n2211 ,n2166 ,n2165);
    nor g268(n2210 ,n1356 ,n2201);
    nor g269(n2209 ,n1355 ,n2200);
    or g270(n2208 ,n2007 ,n2190);
    nor g271(n2207 ,n1914 ,n2177);
    or g272(n2206 ,n2406 ,n2400);
    or g273(n2205 ,n2151 ,n2152);
    nor g274(n2222 ,n2404 ,n2405);
    or g275(n2221 ,n2399 ,n2401);
    or g276(n7[17] ,n1813 ,n2070);
    or g277(n2204 ,n1816 ,n2111);
    or g278(n7[16] ,n1812 ,n2068);
    or g279(n2203 ,n1811 ,n2110);
    or g280(n7[23] ,n1781 ,n2061);
    or g281(n7[18] ,n1817 ,n2071);
    or g282(n2202 ,n1802 ,n2104);
    nor g283(n2201 ,n1423 ,n2134);
    nor g284(n2200 ,n1897 ,n2133);
    or g285(n2199 ,n2130 ,n2129);
    or g286(n2198 ,n2128 ,n2127);
    or g287(n2197 ,n2126 ,n2125);
    or g288(n2196 ,n2124 ,n2123);
    or g289(n2195 ,n2121 ,n2122);
    or g290(n7[22] ,n1778 ,n2049);
    or g291(n2194 ,n1425 ,n2120);
    or g292(n2193 ,n1518 ,n2119);
    or g293(n2192 ,n2115 ,n2114);
    or g294(n2191 ,n2054 ,n2113);
    or g295(n2190 ,n1779 ,n2112);
    or g296(n7[21] ,n1774 ,n2047);
    or g297(n2189 ,n1775 ,n2100);
    or g298(n7[20] ,n1772 ,n2046);
    or g299(n7[19] ,n1769 ,n2072);
    or g300(n2188 ,n1864 ,n2109);
    or g301(n2187 ,n1863 ,n2107);
    or g302(n2186 ,n1862 ,n2106);
    or g303(n2185 ,n2011 ,n2105);
    or g304(n2184 ,n1710 ,n2135);
    or g305(n2183 ,n1698 ,n2147);
    or g306(n2182 ,n1849 ,n2099);
    or g307(n2181 ,n2089 ,n2085);
    or g308(n2180 ,n2090 ,n2097);
    or g309(n2179 ,n2088 ,n2096);
    not g310(n2178 ,n2406);
    or g311(n2176 ,n2086 ,n2095);
    or g312(n2175 ,n2082 ,n2081);
    or g313(n2174 ,n2080 ,n2079);
    or g314(n2173 ,n2078 ,n2077);
    or g315(n2172 ,n2076 ,n2074);
    or g316(n2171 ,n2139 ,n2060);
    or g317(n2170 ,n2140 ,n2059);
    or g318(n2169 ,n2058 ,n2057);
    or g319(n2168 ,n2056 ,n2067);
    or g320(n2167 ,n2102 ,n2055);
    or g321(n2166 ,n2138 ,n2150);
    or g322(n2165 ,n2149 ,n2142);
    or g323(n2164 ,n2137 ,n2053);
    or g324(n2163 ,n2148 ,n2052);
    or g325(n2162 ,n2066 ,n2051);
    or g326(n2161 ,n2141 ,n2050);
    or g327(n2160 ,n2145 ,n2062);
    or g328(n2159 ,n2144 ,n2143);
    or g329(n2158 ,n2048 ,n2065);
    or g330(n2157 ,n2101 ,n2093);
    or g331(n2156 ,n2073 ,n2092);
    xnor g332(n2155 ,n1[12] ,n1924);
    xnor g333(n2154 ,n1[9] ,n1929);
    xnor g334(n2153 ,n1[9] ,n1948);
    xnor g335(n2152 ,n1[1] ,n1937);
    xnor g336(n2151 ,n1[3] ,n1934);
    xnor g337(n2400 ,n1[0] ,n2039);
    xnor g338(n2405 ,n1[2] ,n2040);
    xnor g339(n2399 ,n1[7] ,n1932);
    xnor g340(n2404 ,n1[3] ,n2043);
    xnor g341(n2406 ,n1[1] ,n2044);
    xnor g342(n2402 ,n1[5] ,n2045);
    xnor g343(n2401 ,n1[6] ,n1933);
    xnor g344(n2177 ,n1467 ,n1955);
    or g345(n7[25] ,n2032 ,n1785);
    nor g346(n2150 ,n1092 ,n1945);
    nor g347(n2149 ,n1091 ,n1921);
    nor g348(n2148 ,n1094 ,n1950);
    nor g349(n2147 ,n1093 ,n1954);
    nor g350(n2146 ,n1092 ,n1926);
    nor g351(n2145 ,n1091 ,n1923);
    nor g352(n2144 ,n1095 ,n2042);
    nor g353(n2143 ,n1036 ,n1928);
    nor g354(n2142 ,n1036 ,n1947);
    nor g355(n2141 ,n1090 ,n1931);
    nor g356(n2140 ,n1085 ,n1939);
    nor g357(n2139 ,n1029 ,n1943);
    nor g358(n2138 ,n1082 ,n1936);
    nor g359(n2137 ,n1027 ,n1941);
    or g360(n2136 ,n1814 ,n1981);
    or g361(n2135 ,n1798 ,n1979);
    or g362(n2134 ,n1745 ,n1990);
    or g363(n2133 ,n1696 ,n1988);
    or g364(n2132 ,n1978 ,n1977);
    or g365(n2131 ,n1976 ,n1975);
    or g366(n2130 ,n1026 ,n1974);
    or g367(n2129 ,n1973 ,n1972);
    or g368(n2128 ,n1971 ,n1919);
    or g369(n2127 ,n1970 ,n1969);
    or g370(n2126 ,n1918 ,n1968);
    or g371(n2125 ,n1966 ,n1967);
    or g372(n2124 ,n1965 ,n1917);
    or g373(n2123 ,n1964 ,n1963);
    or g374(n2122 ,n1960 ,n1959);
    or g375(n2121 ,n1961 ,n1962);
    or g376(n2120 ,n1427 ,n1986);
    or g377(n2119 ,n1517 ,n2021);
    or g378(n2118 ,n1791 ,n1985);
    or g379(n2117 ,n2020 ,n2019);
    or g380(n2116 ,n1784 ,n1984);
    or g381(n2115 ,n2016 ,n2015);
    or g382(n2114 ,n2014 ,n2013);
    or g383(n2113 ,n1958 ,n1957);
    or g384(n2112 ,n1777 ,n1956);
    or g385(n2111 ,n2002 ,n1815);
    or g386(n7[30] ,n2037 ,n1795);
    or g387(n2110 ,n1736 ,n2038);
    or g388(n2109 ,n1728 ,n1994);
    or g389(n2108 ,n1865 ,n1995);
    or g390(n2107 ,n1740 ,n1993);
    or g391(n2106 ,n1563 ,n1992);
    or g392(n2105 ,n1861 ,n1991);
    or g393(n2104 ,n2004 ,n1801);
    or g394(n2103 ,n1880 ,n1980);
    or g395(n7[29] ,n2034 ,n1794);
    or g396(n7[27] ,n2035 ,n1789);
    or g397(n7[26] ,n2033 ,n1818);
    or g398(n7[28] ,n2036 ,n1792);
    or g399(n7[24] ,n2031 ,n1782);
    nor g400(n2102 ,n1095 ,n1952);
    nor g401(n2101 ,n1415 ,n1951);
    or g402(n2100 ,n1851 ,n1983);
    or g403(n2099 ,n1750 ,n1982);
    nor g404(n2098 ,n1914 ,n2045);
    nor g405(n2097 ,n1914 ,n2043);
    nor g406(n2096 ,n1914 ,n2040);
    nor g407(n2095 ,n1914 ,n2044);
    nor g408(n2094 ,n1914 ,n2039);
    nor g409(n2093 ,n1914 ,n1932);
    nor g410(n2092 ,n1914 ,n1933);
    nor g411(n2091 ,n1415 ,n1949);
    nor g412(n2090 ,n1415 ,n1944);
    nor g413(n2089 ,n1415 ,n1938);
    nor g414(n2088 ,n1415 ,n1946);
    nor g415(n2087 ,n1415 ,n1940);
    nor g416(n2086 ,n1415 ,n1948);
    nor g417(n2085 ,n1456 ,n2041);
    nor g418(n2084 ,n1456 ,n1922);
    nor g419(n2083 ,n1456 ,n1953);
    nor g420(n2082 ,n1415 ,n1942);
    nor g421(n2081 ,n1456 ,n1924);
    nor g422(n2080 ,n1415 ,n1934);
    nor g423(n2079 ,n1456 ,n1925);
    nor g424(n2078 ,n1415 ,n1935);
    nor g425(n2077 ,n1456 ,n1927);
    nor g426(n2076 ,n1415 ,n1937);
    nor g427(n2075 ,n1456 ,n1930);
    nor g428(n2074 ,n1456 ,n1929);
    or g429(n7[31] ,n1996 ,n1797);
    nor g430(n2073 ,n1415 ,n1920);
    or g431(n2072 ,n2029 ,n1871);
    or g432(n2071 ,n2030 ,n1870);
    or g433(n2070 ,n2028 ,n1868);
    or g434(n2069 ,n2001 ,n1867);
    or g435(n2068 ,n2027 ,n1866);
    nor g436(n2067 ,n1[12] ,n1949);
    nor g437(n2066 ,n1[11] ,n1925);
    nor g438(n2065 ,n1[14] ,n1922);
    or g439(n2064 ,n2009 ,n1858);
    or g440(n2063 ,n2008 ,n1856);
    nor g441(n2062 ,n1[8] ,n1930);
    or g442(n2061 ,n2026 ,n1853);
    nor g443(n2060 ,n1[7] ,n1938);
    nor g444(n2059 ,n1[10] ,n1946);
    nor g445(n2058 ,n1[6] ,n1940);
    nor g446(n2057 ,n1[15] ,n1951);
    nor g447(n2056 ,n1[4] ,n1942);
    nor g448(n2055 ,n1[2] ,n1935);
    or g449(n2054 ,n1915 ,n1916);
    nor g450(n2053 ,n1[14] ,n1920);
    nor g451(n2052 ,n1[11] ,n1944);
    nor g452(n2051 ,n1[10] ,n1927);
    nor g453(n2050 ,n1[13] ,n1953);
    or g454(n2049 ,n2025 ,n1857);
    nor g455(n2048 ,n1[15] ,n2041);
    or g456(n2047 ,n2024 ,n1850);
    or g457(n2046 ,n2023 ,n1848);
    not g458(n2042 ,n2041);
    or g459(n2038 ,n1553 ,n1810);
    nor g460(n2037 ,n1070 ,n1913);
    nor g461(n2036 ,n1134 ,n1913);
    nor g462(n2035 ,n1075 ,n1913);
    nor g463(n2034 ,n1133 ,n1913);
    nor g464(n2033 ,n1131 ,n1913);
    nor g465(n2032 ,n1136 ,n1913);
    nor g466(n2031 ,n1126 ,n1913);
    nor g467(n2030 ,n1056 ,n1913);
    nor g468(n2029 ,n1119 ,n1913);
    nor g469(n2028 ,n1120 ,n1913);
    nor g470(n2027 ,n1058 ,n1913);
    nor g471(n2026 ,n1122 ,n1913);
    nor g472(n2025 ,n1059 ,n1913);
    nor g473(n2024 ,n1057 ,n1913);
    nor g474(n2023 ,n1121 ,n1913);
    or g475(n2022 ,n1118 ,n1899);
    or g476(n2021 ,n1790 ,n1894);
    or g477(n2020 ,n1827 ,n1893);
    or g478(n2019 ,n1892 ,n1891);
    or g479(n2018 ,n1890 ,n1889);
    or g480(n2017 ,n1787 ,n1786);
    or g481(n2016 ,n1888 ,n1887);
    or g482(n2015 ,n1886 ,n1885);
    or g483(n2014 ,n1884 ,n1883);
    or g484(n2013 ,n1882 ,n1881);
    nor g485(n2012 ,n1095 ,n1913);
    nor g486(n2011 ,n1091 ,n1913);
    nor g487(n2010 ,n1093 ,n1913);
    nor g488(n2009 ,n1094 ,n1913);
    nor g489(n2008 ,n1092 ,n1913);
    nor g490(n2007 ,n1090 ,n1913);
    nor g491(n2006 ,n1036 ,n1913);
    nor g492(n2005 ,n1089 ,n1913);
    nor g493(n2004 ,n1032 ,n1913);
    nor g494(n2003 ,n1085 ,n1913);
    nor g495(n2002 ,n1083 ,n1913);
    nor g496(n2001 ,n1029 ,n1913);
    nor g497(n2000 ,n1028 ,n1913);
    nor g498(n1999 ,n1082 ,n1913);
    nor g499(n1998 ,n1084 ,n1913);
    nor g500(n1997 ,n1027 ,n1913);
    nor g501(n1996 ,n1129 ,n1913);
    or g502(n1995 ,n1707 ,n1807);
    or g503(n1994 ,n1552 ,n1808);
    or g504(n1993 ,n1743 ,n1805);
    or g505(n1992 ,n1550 ,n1803);
    or g506(n1991 ,n1732 ,n1799);
    or g507(n1990 ,n1152 ,n1898);
    or g508(n1989 ,n1733 ,n1796);
    or g509(n1988 ,n1195 ,n1896);
    or g510(n1987 ,n1562 ,n1800);
    or g511(n1986 ,n1171 ,n1895);
    or g512(n1985 ,n1788 ,n1855);
    or g513(n1984 ,n1854 ,n1783);
    or g514(n1983 ,n1559 ,n1773);
    or g515(n1982 ,n1738 ,n1770);
    or g516(n1981 ,n1869 ,n1822);
    or g517(n1980 ,n1860 ,n1821);
    or g518(n1979 ,n1859 ,n1820);
    or g519(n1978 ,n1901 ,n1911);
    or g520(n1977 ,n1847 ,n1844);
    or g521(n1976 ,n1843 ,n1842);
    or g522(n1975 ,n1841 ,n1910);
    or g523(n1974 ,n1872 ,n1909);
    or g524(n1973 ,n1873 ,n1879);
    or g525(n1972 ,n1840 ,n1826);
    or g526(n1971 ,n1908 ,n1839);
    or g527(n1970 ,n1907 ,n1838);
    or g528(n1969 ,n1837 ,n1878);
    or g529(n1968 ,n1875 ,n1874);
    or g530(n1967 ,n1912 ,n1835);
    or g531(n1966 ,n1906 ,n1836);
    or g532(n1965 ,n1834 ,n1905);
    or g533(n1964 ,n1833 ,n1830);
    or g534(n1963 ,n1877 ,n1846);
    or g535(n1962 ,n1831 ,n1845);
    or g536(n1961 ,n1832 ,n1904);
    or g537(n1960 ,n1829 ,n1903);
    or g538(n1959 ,n1876 ,n1828);
    or g539(n1958 ,n1902 ,n1900);
    or g540(n1957 ,n1780 ,n1776);
    or g541(n1956 ,n1852 ,n1819);
    nor g542(n2494 ,n1078 ,n1823);
    xnor g543(n1955 ,n1230 ,n1470);
    xnor g544(n2045 ,n1480 ,n1479);
    xnor g545(n2044 ,n1482 ,n1469);
    xnor g546(n2043 ,n1477 ,n1478);
    xnor g547(n2041 ,n1566 ,n1575);
    xnor g548(n2040 ,n1468 ,n1475);
    xnor g549(n2039 ,n1484 ,n1483);
    not g550(n1954 ,n1953);
    not g551(n1952 ,n1951);
    not g552(n1950 ,n1949);
    not g553(n1947 ,n1946);
    not g554(n1945 ,n1944);
    not g555(n1943 ,n1942);
    not g556(n1941 ,n1940);
    not g557(n1939 ,n1938);
    not g558(n1936 ,n1935);
    not g559(n1931 ,n1930);
    not g560(n1928 ,n1927);
    not g561(n1926 ,n1925);
    not g562(n1923 ,n1922);
    not g563(n1921 ,n1920);
    xor g564(n6[42] ,n1635 ,n0[42]);
    xor g565(n6[43] ,n1689 ,n0[43]);
    xor g566(n6[55] ,n1686 ,n0[55]);
    xor g567(n6[45] ,n1684 ,n0[45]);
    xor g568(n6[46] ,n1670 ,n0[46]);
    xor g569(n6[47] ,n1675 ,n0[47]);
    xor g570(n6[48] ,n1671 ,n0[48]);
    xor g571(n6[49] ,n1668 ,n0[49]);
    xor g572(n6[33] ,n1665 ,n0[33]);
    xnor g573(n1919 ,n1029 ,n1583);
    xnor g574(n1918 ,n1082 ,n1604);
    xnor g575(n1917 ,n1027 ,n1587);
    xnor g576(n1916 ,n1[5] ,n1589);
    xor g577(n6[2] ,n1660 ,n0[2]);
    xor g578(n6[1] ,n1662 ,n0[1]);
    xor g579(n6[3] ,n1658 ,n0[3]);
    xor g580(n6[50] ,n1666 ,n0[50]);
    xor g581(n6[34] ,n1663 ,n0[34]);
    xor g582(n6[44] ,n1693 ,n0[44]);
    xor g583(n6[5] ,n1654 ,n0[5]);
    xor g584(n6[35] ,n1659 ,n0[35]);
    xor g585(n6[51] ,n1657 ,n0[51]);
    xor g586(n6[4] ,n1656 ,n0[4]);
    xor g587(n6[7] ,n1650 ,n0[7]);
    xor g588(n6[6] ,n1653 ,n0[6]);
    xor g589(n6[36] ,n1655 ,n0[36]);
    xor g590(n6[59] ,n1645 ,n0[59]);
    xor g591(n6[37] ,n1651 ,n0[37]);
    xor g592(n6[38] ,n1649 ,n0[38]);
    xor g593(n6[58] ,n1661 ,n0[58]);
    xor g594(n6[52] ,n1652 ,n0[52]);
    xor g595(n6[57] ,n1673 ,n0[57]);
    xnor g596(n1915 ,n1[13] ,n1606);
    xor g597(n6[16] ,n1631 ,n0[16]);
    xor g598(n6[17] ,n1682 ,n0[17]);
    xor g599(n6[15] ,n1633 ,n0[15]);
    xor g600(n6[13] ,n1639 ,n0[13]);
    xor g601(n6[14] ,n1636 ,n0[14]);
    xor g602(n6[39] ,n1642 ,n0[39]);
    xor g603(n6[12] ,n1640 ,n0[12]);
    xor g604(n6[10] ,n1644 ,n0[10]);
    xor g605(n6[9] ,n1646 ,n0[9]);
    xor g606(n6[8] ,n1648 ,n0[8]);
    xor g607(n6[62] ,n1647 ,n0[62]);
    xor g608(n6[11] ,n1643 ,n0[11]);
    xor g609(n6[61] ,n1677 ,n0[61]);
    xor g610(n6[31] ,n1680 ,n0[31]);
    xor g611(n6[63] ,n1637 ,n0[63]);
    xor g612(n6[30] ,n1669 ,n0[30]);
    xor g613(n6[29] ,n1672 ,n0[29]);
    xor g614(n6[60] ,n1691 ,n0[60]);
    xor g615(n6[56] ,n1679 ,n0[56]);
    xor g616(n6[28] ,n1674 ,n0[28]);
    xor g617(n6[27] ,n1676 ,n0[27]);
    xor g618(n6[26] ,n1678 ,n0[26]);
    xor g619(n6[25] ,n1688 ,n0[25]);
    xor g620(n6[24] ,n1681 ,n0[24]);
    xor g621(n6[23] ,n1683 ,n0[23]);
    xor g622(n6[22] ,n1685 ,n0[22]);
    xor g623(n6[21] ,n1694 ,n0[21]);
    xor g624(n6[19] ,n1690 ,n0[19]);
    xor g625(n6[53] ,n1641 ,n0[53]);
    xor g626(n6[20] ,n1692 ,n0[20]);
    xor g627(n6[18] ,n1687 ,n0[18]);
    xor g628(n6[40] ,n1638 ,n0[40]);
    xor g629(n6[32] ,n1667 ,n0[32]);
    xor g630(n6[0] ,n1664 ,n0[0]);
    xor g631(n6[54] ,n1634 ,n0[54]);
    xor g632(n6[41] ,n1632 ,n0[41]);
    xnor g633(n1953 ,n1476 ,n1272);
    xnor g634(n1951 ,n0[63] ,n1575);
    xnor g635(n1949 ,n0[60] ,n1576);
    xnor g636(n1948 ,n0[57] ,n1567);
    xnor g637(n1946 ,n0[58] ,n1573);
    xnor g638(n1944 ,n0[59] ,n1571);
    xnor g639(n1942 ,n0[4] ,n1570);
    xnor g640(n1940 ,n0[6] ,n1569);
    xnor g641(n1938 ,n0[7] ,n1566);
    xnor g642(n1937 ,n0[1] ,n1574);
    xnor g643(n1935 ,n0[2] ,n1572);
    xnor g644(n1934 ,n0[3] ,n1565);
    xnor g645(n1933 ,n1471 ,n1481);
    xnor g646(n1932 ,n1473 ,n1472);
    xnor g647(n1930 ,n1474 ,n1357);
    xnor g648(n1929 ,n1567 ,n1574);
    xnor g649(n1927 ,n1572 ,n1573);
    xnor g650(n1925 ,n1565 ,n1571);
    xnor g651(n1924 ,n1570 ,n1576);
    xnor g652(n1922 ,n1569 ,n1568);
    xnor g653(n1920 ,n0[62] ,n1568);
    nor g654(n1912 ,n1093 ,n1611);
    nor g655(n2495 ,n1080 ,n1768);
    nor g656(n2496 ,n1077 ,n1768);
    nor g657(n1911 ,n1[20] ,n1597);
    nor g658(n1910 ,n1059 ,n1581);
    nor g659(n1909 ,n1121 ,n1596);
    nor g660(n1908 ,n1120 ,n1618);
    nor g661(n1907 ,n1058 ,n1617);
    nor g662(n1906 ,n1057 ,n1586);
    nor g663(n1905 ,n1119 ,n1598);
    nor g664(n1904 ,n1122 ,n1577);
    nor g665(n1903 ,n1056 ,n1602);
    nor g666(n1902 ,n1090 ,n1593);
    nor g667(n1901 ,n1[11] ,n1591);
    nor g668(n1900 ,n1032 ,n1595);
    nor g669(n1899 ,n1394 ,n1521);
    or g670(n1898 ,n1248 ,n1746);
    or g671(n1897 ,n1249 ,n1695);
    or g672(n1896 ,n1321 ,n1697);
    or g673(n1895 ,n1314 ,n1747);
    or g674(n1894 ,n1516 ,n1515);
    or g675(n1893 ,n1514 ,n1513);
    or g676(n1892 ,n1512 ,n1511);
    or g677(n1891 ,n1522 ,n1510);
    or g678(n1890 ,n1509 ,n1508);
    or g679(n1889 ,n1524 ,n1507);
    or g680(n1888 ,n1519 ,n1525);
    or g681(n1887 ,n1506 ,n1505);
    or g682(n1886 ,n1504 ,n1503);
    or g683(n1885 ,n1494 ,n1502);
    or g684(n1884 ,n1501 ,n1500);
    or g685(n1883 ,n1493 ,n1499);
    or g686(n1882 ,n1495 ,n1498);
    or g687(n1881 ,n1497 ,n1496);
    nor g688(n1880 ,n1050 ,n1523);
    nor g689(n1879 ,n1095 ,n1620);
    nor g690(n1878 ,n1092 ,n1590);
    nor g691(n2497 ,n1137 ,n1768);
    nor g692(n1877 ,n1094 ,n1609);
    nor g693(n1876 ,n1091 ,n1614);
    nor g694(n1875 ,n1036 ,n1626);
    nor g695(n1874 ,n1089 ,n1624);
    nor g696(n2498 ,n1361 ,n1768);
    nor g697(n1873 ,n1032 ,n1623);
    nor g698(n1872 ,n1085 ,n1628);
    nor g699(n1871 ,n1414 ,n1608);
    nor g700(n1870 ,n1414 ,n1605);
    nor g701(n1869 ,n1414 ,n1585);
    nor g702(n1868 ,n1414 ,n1601);
    nor g703(n1867 ,n1414 ,n1597);
    nor g704(n1866 ,n1414 ,n1622);
    nor g705(n1865 ,n1414 ,n1621);
    nor g706(n1864 ,n1414 ,n1599);
    nor g707(n1863 ,n1414 ,n1603);
    nor g708(n1862 ,n1414 ,n1619);
    nor g709(n1861 ,n1414 ,n1615);
    nor g710(n1860 ,n1414 ,n1616);
    nor g711(n1859 ,n1414 ,n1612);
    nor g712(n1858 ,n1414 ,n1610);
    nor g713(n1857 ,n1414 ,n1588);
    nor g714(n1856 ,n1414 ,n1591);
    nor g715(n1855 ,n1414 ,n1627);
    nor g716(n1854 ,n1414 ,n1625);
    nor g717(n1853 ,n1414 ,n1629);
    nor g718(n1852 ,n1414 ,n1613);
    nor g719(n1851 ,n1414 ,n1578);
    nor g720(n1850 ,n1414 ,n1580);
    nor g721(n1849 ,n1414 ,n1582);
    nor g722(n1848 ,n1414 ,n1584);
    nor g723(n1847 ,n1028 ,n1607);
    nor g724(n1846 ,n1083 ,n1579);
    nor g725(n1845 ,n1084 ,n1600);
    or g726(n2376 ,n3 ,n2375);
    or g727(n1914 ,n1055 ,n2375);
    nor g728(n1913 ,n1055 ,n1630);
    nor g729(n1844 ,n1[16] ,n1616);
    nor g730(n1843 ,n1[13] ,n1612);
    nor g731(n1842 ,n1[7] ,n1629);
    nor g732(n1841 ,n1[15] ,n1621);
    nor g733(n1840 ,n1[1] ,n1601);
    nor g734(n1839 ,n1[22] ,n1582);
    nor g735(n1838 ,n1[14] ,n1615);
    nor g736(n1837 ,n1[12] ,n1610);
    nor g737(n1836 ,n1[9] ,n1625);
    nor g738(n1835 ,n1[21] ,n1585);
    nor g739(n1834 ,n1[23] ,n1578);
    nor g740(n1833 ,n1[18] ,n1603);
    nor g741(n1832 ,n1[5] ,n1580);
    nor g742(n1831 ,n1[3] ,n1608);
    nor g743(n1830 ,n1[10] ,n1627);
    nor g744(n1829 ,n1[19] ,n1599);
    nor g745(n1828 ,n1[17] ,n1619);
    or g746(n1827 ,n1488 ,n1526);
    nor g747(n1826 ,n1[0] ,n1622);
    nor g748(n1825 ,n1205 ,n1768);
    nor g749(n1824 ,n1316 ,n1768);
    nor g750(n1822 ,n1415 ,n1606);
    nor g751(n1821 ,n1415 ,n1592);
    nor g752(n1820 ,n1415 ,n1589);
    nor g753(n1819 ,n1415 ,n1594);
    or g754(n1818 ,n1717 ,n1537);
    or g755(n1817 ,n1704 ,n1558);
    or g756(n1816 ,n1760 ,n1699);
    or g757(n1815 ,n1767 ,n1748);
    or g758(n1814 ,n1735 ,n1557);
    or g759(n1813 ,n1705 ,n1556);
    or g760(n1812 ,n1706 ,n1555);
    or g761(n1811 ,n1739 ,n1759);
    or g762(n1810 ,n1766 ,n1700);
    or g763(n1809 ,n1765 ,n1749);
    or g764(n1808 ,n1742 ,n1758);
    or g765(n1807 ,n1564 ,n1551);
    or g766(n1806 ,n1764 ,n1757);
    or g767(n1805 ,n1729 ,n1554);
    or g768(n1804 ,n1744 ,n1756);
    or g769(n1803 ,n1763 ,n1730);
    or g770(n1802 ,n1762 ,n1549);
    or g771(n1801 ,n1755 ,n1701);
    or g772(n1800 ,n1709 ,n1536);
    or g773(n1799 ,n1708 ,n1548);
    or g774(n1798 ,n1561 ,n1544);
    or g775(n1797 ,n1711 ,n1540);
    or g776(n1796 ,n1712 ,n1543);
    or g777(n1795 ,n1721 ,n1547);
    or g778(n1794 ,n1713 ,n1538);
    or g779(n1793 ,n1489 ,n1485);
    or g780(n1792 ,n1715 ,n1542);
    or g781(n1791 ,n1722 ,n1541);
    or g782(n1790 ,n1490 ,n1487);
    or g783(n1789 ,n1716 ,n1539);
    or g784(n1788 ,n1731 ,n1753);
    or g785(n1787 ,n1492 ,n1491);
    or g786(n1786 ,n1520 ,n1486);
    or g787(n1785 ,n1714 ,n1535);
    or g788(n1784 ,n1752 ,n1534);
    or g789(n1783 ,n1718 ,n1560);
    or g790(n1782 ,n1719 ,n1533);
    or g791(n1781 ,n1720 ,n1532);
    nor g792(n1780 ,n1[8] ,n1592);
    or g793(n1779 ,n1724 ,n1546);
    or g794(n1778 ,n1723 ,n1531);
    or g795(n1777 ,n1734 ,n1751);
    nor g796(n1776 ,n1[0] ,n1594);
    or g797(n1775 ,n1754 ,n1545);
    or g798(n1774 ,n1725 ,n1530);
    or g799(n1773 ,n1737 ,n1702);
    or g800(n1772 ,n1726 ,n1529);
    or g801(n1771 ,n1761 ,n1703);
    or g802(n1770 ,n1741 ,n1528);
    or g803(n1769 ,n1727 ,n1527);
    nor g804(n1767 ,n1066 ,n1466);
    nor g805(n1766 ,n1071 ,n1466);
    nor g806(n1765 ,n1073 ,n1466);
    nor g807(n1764 ,n1128 ,n1466);
    nor g808(n1763 ,n1062 ,n1466);
    nor g809(n1762 ,n1063 ,n1466);
    nor g810(n1761 ,n1067 ,n1466);
    nor g811(n1760 ,n1135 ,n1457);
    nor g812(n1759 ,n1065 ,n1457);
    nor g813(n1758 ,n1069 ,n1457);
    nor g814(n1757 ,n1068 ,n1457);
    nor g815(n1756 ,n1125 ,n1457);
    nor g816(n1755 ,n1074 ,n1457);
    nor g817(n1754 ,n1127 ,n1457);
    nor g818(n1753 ,n1130 ,n1457);
    nor g819(n1752 ,n1072 ,n1457);
    nor g820(n1751 ,n1064 ,n1457);
    nor g821(n1750 ,n1132 ,n1457);
    nor g822(n1749 ,n1339 ,n1455);
    nor g823(n1748 ,n1336 ,n1455);
    or g824(n1747 ,n1158 ,n1398);
    or g825(n1746 ,n1192 ,n1396);
    or g826(n1745 ,n1177 ,n1397);
    nor g827(n1744 ,n1031 ,n1413);
    nor g828(n1743 ,n1030 ,n1413);
    nor g829(n1742 ,n1086 ,n1413);
    nor g830(n1741 ,n1086 ,n1455);
    nor g831(n1740 ,n1031 ,n1455);
    nor g832(n1739 ,n1030 ,n1455);
    nor g833(n1738 ,n1033 ,n1413);
    nor g834(n1737 ,n1034 ,n1413);
    nor g835(n1736 ,n1088 ,n1413);
    nor g836(n1735 ,n1087 ,n1413);
    nor g837(n1734 ,n1088 ,n1455);
    nor g838(n1733 ,n1033 ,n1455);
    nor g839(n1732 ,n1034 ,n1455);
    nor g840(n1731 ,n1087 ,n1455);
    nor g841(n1730 ,n1038 ,n1456);
    nor g842(n1729 ,n1035 ,n1456);
    nor g843(n1728 ,n1037 ,n1456);
    nor g844(n1727 ,n1039 ,n1413);
    nor g845(n1726 ,n1040 ,n1413);
    nor g846(n1725 ,n1044 ,n1413);
    nor g847(n1724 ,n1046 ,n1413);
    nor g848(n1723 ,n1111 ,n1413);
    nor g849(n1722 ,n1109 ,n1413);
    nor g850(n1721 ,n1042 ,n1413);
    nor g851(n1720 ,n1110 ,n1413);
    nor g852(n1719 ,n1048 ,n1413);
    nor g853(n1718 ,n1106 ,n1413);
    nor g854(n1717 ,n1108 ,n1413);
    nor g855(n1716 ,n1101 ,n1413);
    nor g856(n1715 ,n1100 ,n1413);
    nor g857(n1714 ,n1097 ,n1413);
    nor g858(n1713 ,n1105 ,n1413);
    nor g859(n1712 ,n1102 ,n1413);
    nor g860(n1711 ,n1047 ,n1413);
    nor g861(n1710 ,n1113 ,n1413);
    nor g862(n1709 ,n1041 ,n1413);
    nor g863(n1708 ,n1103 ,n1413);
    nor g864(n1707 ,n1112 ,n1413);
    nor g865(n1706 ,n1043 ,n1413);
    nor g866(n1705 ,n1049 ,n1413);
    nor g867(n1704 ,n1045 ,n1413);
    nor g868(n1703 ,n1107 ,n1456);
    nor g869(n1702 ,n1099 ,n1456);
    nor g870(n1701 ,n1098 ,n1456);
    nor g871(n1700 ,n1096 ,n1456);
    nor g872(n1699 ,n1104 ,n1456);
    or g873(n1698 ,n1428 ,n1418);
    or g874(n1697 ,n1419 ,n1426);
    or g875(n1696 ,n1421 ,n1420);
    or g876(n1695 ,n1142 ,n1395);
    nor g877(n1694 ,n1053 ,n1458);
    nor g878(n1693 ,n1114 ,n1461);
    nor g879(n1692 ,n1114 ,n1458);
    nor g880(n1691 ,n1114 ,n1463);
    nor g881(n1690 ,n1115 ,n1458);
    nor g882(n1689 ,n1115 ,n1461);
    nor g883(n1688 ,n1054 ,n1460);
    nor g884(n1687 ,n1117 ,n1458);
    nor g885(n1686 ,n1052 ,n1462);
    nor g886(n1685 ,n1116 ,n1458);
    nor g887(n1684 ,n1053 ,n1461);
    nor g888(n1683 ,n1052 ,n1458);
    nor g889(n1682 ,n1054 ,n1458);
    nor g890(n1681 ,n1051 ,n1460);
    nor g891(n1680 ,n1052 ,n1460);
    nor g892(n1679 ,n1051 ,n1463);
    nor g893(n1678 ,n1117 ,n1460);
    nor g894(n1677 ,n1053 ,n1463);
    nor g895(n1676 ,n1115 ,n1460);
    nor g896(n1675 ,n1052 ,n1461);
    nor g897(n1674 ,n1114 ,n1460);
    nor g898(n1673 ,n1054 ,n1463);
    nor g899(n1672 ,n1053 ,n1460);
    nor g900(n1671 ,n1051 ,n1462);
    nor g901(n1670 ,n1116 ,n1461);
    nor g902(n1669 ,n1116 ,n1460);
    nor g903(n1668 ,n1054 ,n1462);
    nor g904(n1667 ,n1051 ,n1464);
    nor g905(n1666 ,n1117 ,n1462);
    nor g906(n1665 ,n1054 ,n1464);
    nor g907(n1664 ,n1051 ,n1465);
    nor g908(n1663 ,n1117 ,n1464);
    nor g909(n1662 ,n1054 ,n1465);
    nor g910(n1661 ,n1117 ,n1463);
    nor g911(n1660 ,n1117 ,n1465);
    nor g912(n1659 ,n1115 ,n1464);
    nor g913(n1658 ,n1115 ,n1465);
    nor g914(n1657 ,n1115 ,n1462);
    nor g915(n1656 ,n1114 ,n1465);
    nor g916(n1655 ,n1114 ,n1464);
    nor g917(n1654 ,n1053 ,n1465);
    nor g918(n1653 ,n1116 ,n1465);
    nor g919(n1652 ,n1114 ,n1462);
    nor g920(n1651 ,n1053 ,n1464);
    nor g921(n1650 ,n1052 ,n1465);
    nor g922(n1649 ,n1116 ,n1464);
    nor g923(n1648 ,n1051 ,n1459);
    nor g924(n1647 ,n1116 ,n1463);
    nor g925(n1646 ,n1054 ,n1459);
    nor g926(n1645 ,n1115 ,n1463);
    nor g927(n1644 ,n1117 ,n1459);
    nor g928(n1643 ,n1115 ,n1459);
    nor g929(n1642 ,n1052 ,n1464);
    nor g930(n1641 ,n1053 ,n1462);
    nor g931(n1640 ,n1114 ,n1459);
    nor g932(n1639 ,n1053 ,n1459);
    nor g933(n1638 ,n1051 ,n1461);
    nor g934(n1637 ,n1052 ,n1463);
    nor g935(n1636 ,n1116 ,n1459);
    nor g936(n1635 ,n1117 ,n1461);
    nor g937(n1634 ,n1116 ,n1462);
    nor g938(n1633 ,n1052 ,n1459);
    nor g939(n1632 ,n1054 ,n1461);
    nor g940(n1631 ,n1051 ,n1458);
    or g941(n2375 ,n1173 ,n1417);
    or g942(n1768 ,n3 ,n1439);
    not g943(n11 ,n1630);
    not g944(n1629 ,n1628);
    not g945(n1627 ,n1626);
    not g946(n1625 ,n1624);
    not g947(n1623 ,n1622);
    not g948(n1621 ,n1620);
    not g949(n1619 ,n1618);
    not g950(n1617 ,n1616);
    not g951(n1615 ,n1614);
    not g952(n1612 ,n1611);
    not g953(n1610 ,n1609);
    not g954(n1608 ,n1607);
    not g955(n1605 ,n1604);
    not g956(n1603 ,n1602);
    not g957(n1601 ,n1600);
    not g958(n1599 ,n1598);
    not g959(n1597 ,n1596);
    not g960(n1595 ,n1594);
    not g961(n1593 ,n1592);
    not g962(n1591 ,n1590);
    not g963(n1588 ,n1587);
    not g964(n1586 ,n1585);
    not g965(n1584 ,n1583);
    not g966(n1582 ,n1581);
    not g967(n1580 ,n1579);
    not g968(n1578 ,n1577);
    nor g969(n1564 ,n1341 ,n1455);
    nor g970(n1563 ,n1331 ,n1455);
    nor g971(n1562 ,n1342 ,n1455);
    nor g972(n1561 ,n1333 ,n1455);
    nor g973(n1560 ,n1337 ,n1455);
    nor g974(n1559 ,n1344 ,n1455);
    nor g975(n1558 ,n1353 ,n1411);
    nor g976(n1557 ,n1342 ,n1411);
    nor g977(n1556 ,n1360 ,n1411);
    nor g978(n1555 ,n1347 ,n1411);
    nor g979(n1554 ,n1336 ,n1411);
    nor g980(n1553 ,n1337 ,n1411);
    nor g981(n1552 ,n1344 ,n1411);
    nor g982(n1551 ,n1366 ,n1411);
    nor g983(n1550 ,n1339 ,n1411);
    nor g984(n1549 ,n1331 ,n1411);
    nor g985(n1548 ,n1266 ,n1411);
    nor g986(n1547 ,n1251 ,n1411);
    nor g987(n1546 ,n1255 ,n1411);
    nor g988(n1545 ,n1341 ,n1411);
    nor g989(n1544 ,n1274 ,n1411);
    nor g990(n1543 ,n1258 ,n1411);
    nor g991(n1542 ,n1253 ,n1411);
    nor g992(n1541 ,n1256 ,n1411);
    nor g993(n1540 ,n1280 ,n1411);
    nor g994(n1539 ,n1286 ,n1411);
    nor g995(n1538 ,n1278 ,n1411);
    nor g996(n1537 ,n1260 ,n1411);
    nor g997(n1536 ,n1288 ,n1411);
    nor g998(n1535 ,n1282 ,n1411);
    nor g999(n1534 ,n1276 ,n1411);
    nor g1000(n1533 ,n1262 ,n1411);
    nor g1001(n1532 ,n1359 ,n1411);
    nor g1002(n1531 ,n1349 ,n1411);
    nor g1003(n1530 ,n1284 ,n1411);
    nor g1004(n1529 ,n1264 ,n1411);
    nor g1005(n1528 ,n1333 ,n1411);
    nor g1006(n1527 ,n1364 ,n1411);
    or g1007(n1526 ,n1389 ,n1435);
    or g1008(n1525 ,n1390 ,n1438);
    or g1009(n1524 ,n1374 ,n1387);
    nor g1010(n1523 ,n1454 ,n1412);
    or g1011(n1522 ,n1386 ,n1378);
    or g1012(n1521 ,n1362 ,n1453);
    xnor g1013(n1520 ,n1[17] ,n1360);
    or g1014(n1519 ,n1371 ,n1445);
    or g1015(n1518 ,n1377 ,n1429);
    or g1016(n1517 ,n1431 ,n1404);
    or g1017(n1516 ,n1392 ,n1381);
    or g1018(n1515 ,n1393 ,n1432);
    or g1019(n1514 ,n1388 ,n1376);
    or g1020(n1513 ,n1373 ,n1447);
    or g1021(n1512 ,n1452 ,n1441);
    or g1022(n1511 ,n1448 ,n1434);
    or g1023(n1510 ,n1380 ,n1408);
    or g1024(n1509 ,n1391 ,n1443);
    or g1025(n1508 ,n1379 ,n1430);
    or g1026(n1507 ,n1437 ,n1406);
    or g1027(n1506 ,n1369 ,n1382);
    or g1028(n1505 ,n1384 ,n1436);
    or g1029(n1504 ,n1400 ,n1375);
    or g1030(n1503 ,n1368 ,n1433);
    or g1031(n1502 ,n1449 ,n1405);
    or g1032(n1501 ,n1383 ,n1450);
    or g1033(n1500 ,n1367 ,n1444);
    or g1034(n1499 ,n1401 ,n1402);
    or g1035(n1498 ,n1446 ,n1403);
    or g1036(n1497 ,n1385 ,n1442);
    or g1037(n1496 ,n1372 ,n1409);
    or g1038(n1495 ,n1451 ,n1407);
    or g1039(n1494 ,n1370 ,n1440);
    or g1040(n1493 ,n1410 ,n1399);
    xnor g1041(n1492 ,n1[23] ,n1359);
    xnor g1042(n1491 ,n1[18] ,n1353);
    xnor g1043(n1490 ,n1[15] ,n1341);
    xnor g1044(n1489 ,n1[9] ,n1337);
    xnor g1045(n1488 ,n1[4] ,n1337);
    xnor g1046(n1487 ,n1[5] ,n1336);
    xnor g1047(n1486 ,n1[10] ,n1256);
    xnor g1048(n1485 ,n1[3] ,n1339);
    xnor g1049(n1484 ,n1333 ,n1336);
    xnor g1050(n1483 ,n1337 ,n1331);
    xnor g1051(n1482 ,n1266 ,n1258);
    xnor g1052(n1481 ,n1235 ,n1236);
    xnor g1053(n1480 ,n1238 ,n1237);
    xnor g1054(n1479 ,n1239 ,n1242);
    nor g1055(n1630 ,n1350 ,n1416);
    xnor g1056(n1478 ,n1253 ,n1262);
    xnor g1057(n1477 ,n1251 ,n1260);
    xnor g1058(n1476 ,n1268 ,n1267);
    xnor g1059(n1475 ,n1264 ,n1347);
    xnor g1060(n1474 ,n1219 ,n1270);
    xnor g1061(n1473 ,n1297 ,n1232);
    xnor g1062(n1472 ,n1231 ,n1300);
    xnor g1063(n1471 ,n1229 ,n1234);
    xnor g1064(n1470 ,n0[37] ,n1208);
    xnor g1065(n1469 ,n1256 ,n1255);
    xnor g1066(n1468 ,n1349 ,n1353);
    xnor g1067(n1467 ,n0[36] ,n1243);
    xnor g1068(n1628 ,n0[55] ,n1298);
    xnor g1069(n1626 ,n0[58] ,n1210);
    xnor g1070(n1624 ,n0[57] ,n1216);
    xnor g1071(n1622 ,n1048 ,n1269);
    xnor g1072(n1620 ,n0[63] ,n1213);
    xnor g1073(n1618 ,n0[17] ,n1227);
    xnor g1074(n1616 ,n1043 ,n1271);
    xnor g1075(n1614 ,n0[62] ,n1209);
    xnor g1076(n1613 ,n1228 ,n1098);
    xnor g1077(n1611 ,n0[61] ,n1215);
    xnor g1078(n1609 ,n0[60] ,n1214);
    xnor g1079(n1607 ,n0[51] ,n1294);
    xnor g1080(n1606 ,n1224 ,n1272);
    xnor g1081(n1604 ,n0[50] ,n1293);
    xnor g1082(n1602 ,n0[58] ,n1221);
    xnor g1083(n1600 ,n0[49] ,n1292);
    xnor g1084(n1598 ,n0[59] ,n1245);
    xnor g1085(n1596 ,n0[44] ,n1226);
    xnor g1086(n1594 ,n1270 ,n1269);
    xnor g1087(n1592 ,n1271 ,n1357);
    xnor g1088(n1590 ,n0[59] ,n1212);
    xnor g1089(n1589 ,n1301 ,n1268);
    xnor g1090(n1587 ,n0[54] ,n1299);
    xnor g1091(n1585 ,n1031 ,n1267);
    xnor g1092(n1583 ,n0[52] ,n1295);
    xnor g1093(n1581 ,n0[46] ,n1290);
    xnor g1094(n1579 ,n0[53] ,n1289);
    xnor g1095(n1577 ,n0[47] ,n1291);
    xnor g1096(n1576 ,n0[44] ,n1296);
    xnor g1097(n1575 ,n0[47] ,n1244);
    xnor g1098(n1574 ,n0[49] ,n1218);
    xnor g1099(n1573 ,n0[42] ,n1222);
    xnor g1100(n1572 ,n0[50] ,n1220);
    xnor g1101(n1571 ,n0[43] ,n1240);
    xnor g1102(n1570 ,n0[52] ,n1217);
    xnor g1103(n1569 ,n0[54] ,n1225);
    xnor g1104(n1568 ,n0[46] ,n1241);
    xnor g1105(n1567 ,n0[41] ,n1233);
    xnor g1106(n1566 ,n0[55] ,n1223);
    xnor g1107(n1565 ,n0[51] ,n1211);
    not g1108(n1455 ,n1454);
    nor g1109(n1453 ,n1141 ,n1302);
    nor g1110(n1452 ,n1136 ,n1281);
    nor g1111(n1451 ,n1133 ,n1277);
    nor g1112(n1450 ,n1075 ,n1285);
    nor g1113(n1449 ,n1129 ,n1279);
    nor g1114(n1448 ,n1131 ,n1259);
    nor g1115(n1447 ,n1126 ,n1261);
    nor g1116(n1446 ,n1134 ,n1252);
    nor g1117(n1445 ,n1070 ,n1250);
    nor g1118(n1444 ,n1057 ,n1283);
    nor g1119(n1443 ,n1119 ,n1363);
    nor g1120(n1442 ,n1058 ,n1346);
    nor g1121(n1441 ,n1059 ,n1348);
    nor g1122(n1440 ,n1121 ,n1263);
    or g1123(n1439 ,n1118 ,n1352);
    nor g1124(n1438 ,n1093 ,n1273);
    nor g1125(n1437 ,n1095 ,n1365);
    nor g1126(n1436 ,n1092 ,n1287);
    nor g1127(n1435 ,n1089 ,n1275);
    nor g1128(n1434 ,n1094 ,n1257);
    nor g1129(n1433 ,n1091 ,n1265);
    nor g1130(n1432 ,n1085 ,n1345);
    nor g1131(n1431 ,n1093 ,n1334);
    nor g1132(n1430 ,n1090 ,n1254);
    nor g1133(n1429 ,n1092 ,n1343);
    or g1134(n1428 ,n1303 ,n1306);
    or g1135(n1427 ,n1329 ,n1310);
    or g1136(n1426 ,n1326 ,n1318);
    or g1137(n1425 ,n1317 ,n1308);
    or g1138(n1424 ,n1304 ,n1307);
    or g1139(n1423 ,n1325 ,n1309);
    or g1140(n1422 ,n1312 ,n1311);
    or g1141(n1421 ,n1315 ,n1324);
    or g1142(n1420 ,n1323 ,n1322);
    or g1143(n1419 ,n1320 ,n1319);
    or g1144(n1418 ,n1305 ,n1313);
    or g1145(n1466 ,n1199 ,n1356);
    or g1146(n1465 ,n1174 ,n1354);
    or g1147(n1464 ,n1174 ,n1358);
    or g1148(n1463 ,n1207 ,n1358);
    or g1149(n1462 ,n1204 ,n1358);
    or g1150(n1461 ,n1201 ,n1358);
    or g1151(n1460 ,n1207 ,n1354);
    or g1152(n1459 ,n1201 ,n1354);
    or g1153(n1458 ,n1204 ,n1354);
    or g1154(n1457 ,n1199 ,n1355);
    or g1155(n1456 ,n1200 ,n1355);
    nor g1156(n1454 ,n1200 ,n1356);
    not g1157(n1417 ,n1416);
    not g1158(n1413 ,n1412);
    nor g1159(n1410 ,n1[14] ,n1266);
    nor g1160(n1409 ,n1032 ,n1332);
    nor g1161(n1408 ,n1028 ,n1345);
    nor g1162(n1407 ,n1083 ,n1343);
    nor g1163(n1406 ,n1084 ,n1338);
    nor g1164(n1405 ,n1027 ,n1334);
    nor g1165(n1404 ,n1084 ,n1332);
    nor g1166(n1403 ,n1082 ,n1335);
    nor g1167(n1402 ,n1085 ,n1340);
    nor g1168(n1401 ,n1[26] ,n1260);
    nor g1169(n1400 ,n1[28] ,n1253);
    nor g1170(n1399 ,n1[0] ,n1331);
    or g1171(n1398 ,n1182 ,n1330);
    or g1172(n1397 ,n1[7] ,n1246);
    or g1173(n1396 ,n1191 ,n1247);
    or g1174(n1395 ,n1[11] ,n1327);
    or g1175(n1394 ,n2427 ,n1352);
    nor g1176(n1393 ,n1[11] ,n1342);
    nor g1177(n1392 ,n1[7] ,n1344);
    nor g1178(n1391 ,n1[1] ,n1339);
    nor g1179(n1390 ,n1[11] ,n1288);
    nor g1180(n1389 ,n1[15] ,n1366);
    nor g1181(n1388 ,n1[21] ,n1284);
    nor g1182(n1387 ,n1[9] ,n1276);
    nor g1183(n1386 ,n1[6] ,n1333);
    nor g1184(n1385 ,n1[29] ,n1278);
    nor g1185(n1384 ,n1[30] ,n1251);
    nor g1186(n1383 ,n1[2] ,n1336);
    nor g1187(n1382 ,n1[5] ,n1342);
    nor g1188(n1381 ,n1[1] ,n1331);
    nor g1189(n1380 ,n1[12] ,n1258);
    nor g1190(n1379 ,n1[19] ,n1364);
    nor g1191(n1378 ,n1[3] ,n1344);
    nor g1192(n1377 ,n1[13] ,n1333);
    nor g1193(n1376 ,n1[20] ,n1264);
    nor g1194(n1375 ,n1[7] ,n1341);
    nor g1195(n1374 ,n1[22] ,n1349);
    nor g1196(n1373 ,n1[25] ,n1282);
    nor g1197(n1372 ,n1[27] ,n1286);
    nor g1198(n1371 ,n1[13] ,n1274);
    nor g1199(n1370 ,n1[8] ,n1255);
    nor g1200(n1369 ,n1[16] ,n1347);
    nor g1201(n1368 ,n1[24] ,n1262);
    nor g1202(n1367 ,n1[31] ,n1280);
    nor g1203(n1416 ,n2[3] ,n1328);
    or g1204(n1415 ,n1200 ,n1351);
    or g1205(n1414 ,n1199 ,n1351);
    nor g1206(n1412 ,n1199 ,n1352);
    or g1207(n1411 ,n1200 ,n1352);
    not g1208(n1366 ,n1365);
    not g1209(n1364 ,n1363);
    not g1210(n1361 ,n1362);
    not g1211(n1351 ,n1350);
    not g1212(n1349 ,n1348);
    not g1213(n1347 ,n1346);
    not g1214(n1344 ,n1345);
    not g1215(n1342 ,n1343);
    not g1216(n1341 ,n1340);
    not g1217(n1339 ,n1338);
    not g1218(n1336 ,n1335);
    not g1219(n1333 ,n1334);
    not g1220(n1331 ,n1332);
    or g1221(n1330 ,n1170 ,n1153);
    or g1222(n1329 ,n2374 ,n1167);
    nor g1223(n1328 ,n1118 ,n1173);
    or g1224(n1327 ,n1188 ,n1143);
    or g1225(n1326 ,n1178 ,n1148);
    or g1226(n1325 ,n1198 ,n1145);
    or g1227(n1324 ,n1190 ,n1150);
    or g1228(n1323 ,n1185 ,n1196);
    or g1229(n1322 ,n1156 ,n1163);
    or g1230(n1321 ,n1187 ,n1186);
    or g1231(n1320 ,n1184 ,n1197);
    or g1232(n1319 ,n1144 ,n1151);
    or g1233(n1318 ,n1160 ,n1172);
    or g1234(n1317 ,n1147 ,n1166);
    nor g1235(n1316 ,n1139 ,n1194);
    or g1236(n1315 ,n1179 ,n1183);
    or g1237(n1314 ,n1168 ,n1165);
    or g1238(n1313 ,n1161 ,n1169);
    or g1239(n1312 ,n1157 ,n1175);
    or g1240(n1311 ,n1146 ,n1193);
    or g1241(n1310 ,n1149 ,n1159);
    or g1242(n1309 ,n1155 ,n1164);
    or g1243(n1308 ,n1181 ,n1162);
    or g1244(n1307 ,n1154 ,n1176);
    xnor g1245(n1306 ,n0[57] ,n1084);
    xnor g1246(n1305 ,n0[56] ,n1032);
    xnor g1247(n1304 ,n1[6] ,n1107);
    xnor g1248(n1303 ,n0[60] ,n1029);
    or g1249(n1302 ,n1140 ,n1206);
    xnor g1250(n1301 ,n0[21] ,n0[5]);
    xnor g1251(n1300 ,n0[57] ,n0[56]);
    xnor g1252(n1299 ,n0[30] ,n0[6]);
    xnor g1253(n1298 ,n0[31] ,n0[7]);
    xnor g1254(n1297 ,n0[59] ,n0[58]);
    xnor g1255(n1296 ,n0[28] ,n0[12]);
    xnor g1256(n1295 ,n0[28] ,n0[4]);
    xnor g1257(n1294 ,n0[27] ,n0[3]);
    xnor g1258(n1293 ,n0[26] ,n0[2]);
    xnor g1259(n1292 ,n0[25] ,n0[1]);
    xnor g1260(n1291 ,n0[23] ,n0[3]);
    xnor g1261(n1290 ,n0[22] ,n0[2]);
    xnor g1262(n1289 ,n0[29] ,n0[5]);
    xnor g1263(n1365 ,n0[15] ,n1043);
    xnor g1264(n1363 ,n0[19] ,n1040);
    nor g1265(n1362 ,n2409 ,n1189);
    xnor g1266(n1360 ,n0[18] ,n0[17]);
    xnor g1267(n1359 ,n0[24] ,n0[23]);
    or g1268(n1358 ,n1079 ,n1203);
    xnor g1269(n1357 ,n1046 ,n1048);
    or g1270(n1356 ,n1124 ,n1202);
    or g1271(n1355 ,n2[2] ,n1202);
    or g1272(n1354 ,n5[5] ,n1203);
    xnor g1273(n1353 ,n1045 ,n1039);
    or g1274(n1352 ,n2[1] ,n1180);
    nor g1275(n1350 ,n1060 ,n1173);
    xnor g1276(n1348 ,n0[22] ,n1110);
    xnor g1277(n1346 ,n0[16] ,n1049);
    xnor g1278(n1345 ,n0[3] ,n1088);
    xnor g1279(n1343 ,n0[5] ,n1033);
    xnor g1280(n1340 ,n0[7] ,n1046);
    xnor g1281(n1338 ,n0[1] ,n1030);
    xnor g1282(n1337 ,n1088 ,n1087);
    xnor g1283(n1335 ,n0[2] ,n1086);
    xnor g1284(n1334 ,n0[6] ,n1034);
    xnor g1285(n1332 ,n1050 ,n0[1]);
    not g1286(n1288 ,n1287);
    not g1287(n1286 ,n1285);
    not g1288(n1284 ,n1283);
    not g1289(n1282 ,n1281);
    not g1290(n1280 ,n1279);
    not g1291(n1278 ,n1277);
    not g1292(n1276 ,n1275);
    not g1293(n1274 ,n1273);
    not g1294(n1266 ,n1265);
    not g1295(n1264 ,n1263);
    not g1296(n1262 ,n1261);
    not g1297(n1260 ,n1259);
    not g1298(n1258 ,n1257);
    not g1299(n1255 ,n1254);
    not g1300(n1253 ,n1252);
    not g1301(n1251 ,n1250);
    xnor g1302(n1249 ,n1[1] ,n1125);
    xnor g1303(n1248 ,n1[4] ,n1071);
    xnor g1304(n1247 ,n1[2] ,n1128);
    xnor g1305(n1246 ,n1[3] ,n1073);
    xnor g1306(n1245 ,n0[43] ,n0[19]);
    xnor g1307(n1244 ,n0[31] ,n0[15]);
    xnor g1308(n1243 ,n0[39] ,n0[38]);
    xnor g1309(n1242 ,n0[41] ,n0[40]);
    xnor g1310(n1241 ,n0[30] ,n0[14]);
    xnor g1311(n1240 ,n0[27] ,n0[11]);
    xnor g1312(n1239 ,n0[43] ,n0[42]);
    xnor g1313(n1238 ,n0[47] ,n0[46]);
    xnor g1314(n1237 ,n0[45] ,n0[44]);
    xnor g1315(n1236 ,n0[49] ,n0[48]);
    xnor g1316(n1235 ,n0[51] ,n0[50]);
    xnor g1317(n1234 ,n0[53] ,n0[52]);
    xnor g1318(n1233 ,n0[25] ,n0[9]);
    xnor g1319(n1232 ,n0[63] ,n0[62]);
    xnor g1320(n1231 ,n0[61] ,n0[60]);
    xnor g1321(n1230 ,n0[35] ,n0[34]);
    xnor g1322(n1229 ,n0[55] ,n0[54]);
    xnor g1323(n1228 ,n0[32] ,n0[8]);
    xnor g1324(n1227 ,n0[57] ,n0[41]);
    xnor g1325(n1226 ,n0[20] ,n0[0]);
    xnor g1326(n1225 ,n0[38] ,n0[22]);
    xnor g1327(n1224 ,n0[61] ,n0[45]);
    xnor g1328(n1223 ,n0[39] ,n0[23]);
    xnor g1329(n1222 ,n0[26] ,n0[10]);
    xnor g1330(n1221 ,n0[42] ,n0[18]);
    xnor g1331(n1220 ,n0[34] ,n0[18]);
    xnor g1332(n1219 ,n0[48] ,n0[40]);
    xnor g1333(n1218 ,n0[33] ,n0[17]);
    xnor g1334(n1217 ,n0[36] ,n0[20]);
    xnor g1335(n1216 ,n0[33] ,n0[9]);
    xnor g1336(n1215 ,n0[37] ,n0[13]);
    xnor g1337(n1214 ,n0[36] ,n0[12]);
    xnor g1338(n1213 ,n0[39] ,n0[15]);
    xnor g1339(n1212 ,n0[35] ,n0[11]);
    xnor g1340(n1211 ,n0[35] ,n0[19]);
    xnor g1341(n1210 ,n0[34] ,n0[10]);
    xnor g1342(n1209 ,n0[38] ,n0[14]);
    xnor g1343(n1208 ,n0[33] ,n0[32]);
    xnor g1344(n1287 ,n0[11] ,n1102);
    xnor g1345(n1285 ,n0[27] ,n1100);
    xnor g1346(n1283 ,n0[21] ,n1111);
    xnor g1347(n1281 ,n0[25] ,n1108);
    xnor g1348(n1279 ,n0[32] ,n1047);
    xnor g1349(n1277 ,n0[29] ,n1042);
    xnor g1350(n1275 ,n0[9] ,n1109);
    xnor g1351(n1273 ,n0[13] ,n1103);
    xnor g1352(n1272 ,n1113 ,n1105);
    xnor g1353(n1271 ,n0[56] ,n0[40]);
    xnor g1354(n1270 ,n0[32] ,n0[16]);
    xnor g1355(n1269 ,n0[48] ,n0[0]);
    xnor g1356(n1268 ,n0[53] ,n0[37]);
    xnor g1357(n1267 ,n0[45] ,n0[21]);
    xnor g1358(n1265 ,n0[14] ,n1112);
    xnor g1359(n1263 ,n0[20] ,n1044);
    xnor g1360(n1261 ,n0[24] ,n1097);
    xnor g1361(n1259 ,n0[26] ,n1101);
    xnor g1362(n1257 ,n0[12] ,n1113);
    xnor g1363(n1256 ,n1109 ,n1041);
    xnor g1364(n1254 ,n0[8] ,n1106);
    xnor g1365(n1252 ,n0[28] ,n1105);
    xnor g1366(n1250 ,n0[30] ,n1047);
    not g1367(n1206 ,n1205);
    nor g1368(n1198 ,n1067 ,n1[6]);
    nor g1369(n1197 ,n1036 ,n2395);
    nor g1370(n1196 ,n1064 ,n1[8]);
    nor g1371(n1195 ,n1074 ,n1[0]);
    nor g1372(n1194 ,n1138 ,n2411);
    nor g1373(n1193 ,n1037 ,n1[3]);
    nor g1374(n1192 ,n1063 ,n1[0]);
    nor g1375(n1191 ,n1062 ,n1[1]);
    nor g1376(n1190 ,n1135 ,n1[5]);
    nor g1377(n1188 ,n1127 ,n1[7]);
    nor g1378(n1187 ,n1065 ,n1[4]);
    nor g1379(n1186 ,n1069 ,n1[3]);
    nor g1380(n1185 ,n1130 ,n1[10]);
    nor g1381(n1184 ,n1068 ,n1[2]);
    nor g1382(n1183 ,n1089 ,n2394);
    nor g1383(n1182 ,n1091 ,n0[7]);
    nor g1384(n1181 ,n1094 ,n0[6]);
    or g1385(n1180 ,n1124 ,n2[3]);
    nor g1386(n1179 ,n1132 ,n1[6]);
    nor g1387(n1178 ,n1072 ,n1[9]);
    nor g1388(n1177 ,n1066 ,n1[5]);
    nor g1389(n1176 ,n1104 ,n1[5]);
    nor g1390(n1175 ,n1099 ,n1[7]);
    or g1391(n1207 ,n1123 ,n1061);
    nor g1392(n1205 ,n1139 ,n1138);
    or g1393(n1204 ,n1123 ,n5[3]);
    nor g1394(n1203 ,n1081 ,n4[1]);
    or g1395(n1202 ,n1076 ,n2[3]);
    or g1396(n1201 ,n1061 ,n5[4]);
    or g1397(n1200 ,n1055 ,n2[0]);
    or g1398(n1199 ,n1118 ,n1055);
    nor g1399(n1172 ,n1082 ,n2387);
    nor g1400(n1171 ,n1090 ,n0[4]);
    nor g1401(n1170 ,n1036 ,n0[5]);
    nor g1402(n1169 ,n1035 ,n1[2]);
    nor g1403(n1168 ,n1087 ,n1[10]);
    nor g1404(n1167 ,n1033 ,n1[12]);
    nor g1405(n1166 ,n1034 ,n1[14]);
    nor g1406(n1165 ,n1088 ,n1[8]);
    nor g1407(n1164 ,n1032 ,n2378);
    nor g1408(n1163 ,n1032 ,n2385);
    nor g1409(n1162 ,n1031 ,n1[2]);
    nor g1410(n1161 ,n1085 ,n0[63]);
    nor g1411(n1160 ,n1085 ,n2392);
    nor g1412(n1159 ,n1086 ,n1[6]);
    nor g1413(n1158 ,n1030 ,n1[4]);
    nor g1414(n1157 ,n1083 ,n0[61]);
    nor g1415(n1156 ,n1090 ,n2393);
    nor g1416(n1155 ,n1027 ,n2384);
    nor g1417(n1154 ,n1028 ,n0[59]);
    nor g1418(n1153 ,n1027 ,n0[3]);
    nor g1419(n1152 ,n1083 ,n2383);
    nor g1420(n1151 ,n1083 ,n2390);
    nor g1421(n1150 ,n1028 ,n2388);
    nor g1422(n1149 ,n1029 ,n0[2]);
    nor g1423(n1148 ,n1029 ,n2389);
    nor g1424(n1147 ,n1082 ,n0[1]);
    nor g1425(n1146 ,n1082 ,n0[58]);
    nor g1426(n1145 ,n1084 ,n2379);
    nor g1427(n1144 ,n1027 ,n2391);
    or g1428(n1143 ,n1[15] ,n1[14]);
    or g1429(n1142 ,n1[13] ,n1[12]);
    or g1430(n1174 ,n5[4] ,n5[3]);
    or g1431(n1173 ,n2[2] ,n2[1]);
    not g1432(n1141 ,n2410);
    not g1433(n1140 ,n2411);
    not g1434(n1139 ,n2396);
    not g1435(n1138 ,n2397);
    not g1436(n1137 ,n2408);
    not g1437(n1136 ,n1[25]);
    not g1438(n1135 ,n2390);
    not g1439(n1134 ,n1[28]);
    not g1440(n1133 ,n1[29]);
    not g1441(n1132 ,n2391);
    not g1442(n1131 ,n1[26]);
    not g1443(n1130 ,n2395);
    not g1444(n1129 ,n1[31]);
    not g1445(n1128 ,n2380);
    not g1446(n1127 ,n2392);
    not g1447(n1126 ,n1[24]);
    not g1448(n1125 ,n2386);
    not g1449(n1124 ,n2[2]);
    not g1450(n1123 ,n5[4]);
    not g1451(n1122 ,n1[23]);
    not g1452(n1121 ,n1[20]);
    not g1453(n1120 ,n1[17]);
    not g1454(n1119 ,n1[19]);
    not g1455(n1118 ,n2[0]);
    not g1456(n1117 ,n2417);
    not g1457(n1116 ,n2421);
    not g1458(n1115 ,n2418);
    not g1459(n1114 ,n2419);
    not g1460(n1113 ,n0[13]);
    not g1461(n1112 ,n0[15]);
    not g1462(n1111 ,n0[22]);
    not g1463(n1110 ,n0[23]);
    not g1464(n1109 ,n0[10]);
    not g1465(n1108 ,n0[26]);
    not g1466(n1107 ,n0[62]);
    not g1467(n1106 ,n0[9]);
    not g1468(n1105 ,n0[29]);
    not g1469(n1104 ,n0[61]);
    not g1470(n1103 ,n0[14]);
    not g1471(n1102 ,n0[12]);
    not g1472(n1101 ,n0[27]);
    not g1473(n1100 ,n0[28]);
    not g1474(n1099 ,n0[63]);
    not g1475(n1098 ,n0[56]);
    not g1476(n1097 ,n0[25]);
    not g1477(n1096 ,n0[60]);
    not g1478(n1095 ,n1[15]);
    not g1479(n1094 ,n1[12]);
    not g1480(n1093 ,n1[13]);
    not g1481(n1092 ,n1[11]);
    not g1482(n1091 ,n1[14]);
    not g1483(n1090 ,n1[8]);
    not g1484(n1089 ,n1[9]);
    not g1485(n1088 ,n0[4]);
    not g1486(n1087 ,n0[5]);
    not g1487(n1086 ,n0[3]);
    not g1488(n1085 ,n1[7]);
    not g1489(n1084 ,n1[1]);
    not g1490(n1083 ,n1[5]);
    not g1491(n1082 ,n1[2]);
    not g1492(n1081 ,n2423);
    not g1493(n1080 ,n2409);
    not g1494(n1079 ,n5[5]);
    not g1495(n1078 ,n2427);
    not g1496(n1077 ,n2407);
    not g1497(n1076 ,n2[1]);
    not g1498(n1075 ,n1[27]);
    not g1499(n1074 ,n2385);
    not g1500(n1073 ,n2381);
    not g1501(n1072 ,n2394);
    not g1502(n1071 ,n2382);
    not g1503(n1070 ,n1[30]);
    not g1504(n1069 ,n2388);
    not g1505(n1068 ,n2387);
    not g1506(n1067 ,n2384);
    not g1507(n1066 ,n2383);
    not g1508(n1065 ,n2389);
    not g1509(n1064 ,n2393);
    not g1510(n1063 ,n2378);
    not g1511(n1062 ,n2379);
    not g1512(n1061 ,n5[3]);
    not g1513(n1060 ,n2[3]);
    not g1514(n1059 ,n1[22]);
    not g1515(n1058 ,n1[16]);
    not g1516(n1057 ,n1[21]);
    not g1517(n1056 ,n1[18]);
    not g1518(n1055 ,n3);
    not g1519(n1054 ,n2416);
    not g1520(n1053 ,n2420);
    not g1521(n1052 ,n2422);
    not g1522(n1051 ,n2415);
    not g1523(n1050 ,n0[0]);
    not g1524(n1049 ,n0[17]);
    not g1525(n1048 ,n0[24]);
    not g1526(n1047 ,n0[31]);
    not g1527(n1046 ,n0[8]);
    not g1528(n1045 ,n0[18]);
    not g1529(n1044 ,n0[21]);
    not g1530(n1043 ,n0[16]);
    not g1531(n1042 ,n0[30]);
    not g1532(n1041 ,n0[11]);
    not g1533(n1040 ,n0[20]);
    not g1534(n1039 ,n0[19]);
    not g1535(n1038 ,n0[57]);
    not g1536(n1037 ,n0[59]);
    not g1537(n1036 ,n1[10]);
    not g1538(n1035 ,n0[58]);
    not g1539(n1034 ,n0[7]);
    not g1540(n1033 ,n0[6]);
    not g1541(n1032 ,n1[0]);
    not g1542(n1031 ,n0[1]);
    not g1543(n1030 ,n0[2]);
    not g1544(n1029 ,n1[4]);
    not g1545(n1028 ,n1[3]);
    not g1546(n1027 ,n1[6]);
    xor g1547(n1026 ,n1090 ,n1613);
    xnor g1548(n2398 ,n54 ,n39);
    nor g1549(n2412 ,n40 ,n54);
    xor g1550(n2413 ,n52 ,n49);
    nor g1551(n54 ,n48 ,n53);
    nor g1552(n53 ,n51 ,n50);
    nor g1553(n52 ,n51 ,n48);
    xor g1554(n2414 ,n37 ,n44);
    nor g1555(n51 ,n47 ,n42);
    not g1556(n50 ,n49);
    nor g1557(n49 ,n38 ,n45);
    nor g1558(n48 ,n46 ,n41);
    not g1559(n47 ,n46);
    nor g1560(n46 ,n27 ,n43);
    not g1561(n45 ,n44);
    xnor g1562(n44 ,n29 ,n35);
    nor g1563(n43 ,n23 ,n36);
    not g1564(n42 ,n41);
    xnor g1565(n41 ,n34 ,n33);
    not g1566(n40 ,n39);
    nor g1567(n39 ,n34 ,n33);
    not g1568(n38 ,n37);
    xnor g1569(n37 ,n2400 ,n28);
    not g1570(n36 ,n35);
    xnor g1571(n35 ,n30 ,n2402);
    nor g1572(n34 ,n26 ,n32);
    nor g1573(n33 ,n25 ,n31);
    nor g1574(n32 ,n21 ,n22);
    nor g1575(n31 ,n17 ,n24);
    xnor g1576(n30 ,n2405 ,n2401);
    xnor g1577(n29 ,n2404 ,n2403);
    xnor g1578(n28 ,n2406 ,n2399);
    nor g1579(n27 ,n20 ,n18);
    nor g1580(n26 ,n15 ,n14);
    nor g1581(n25 ,n16 ,n19);
    nor g1582(n24 ,n2406 ,n2400);
    nor g1583(n23 ,n2404 ,n2403);
    nor g1584(n22 ,n2405 ,n2402);
    not g1585(n21 ,n2401);
    not g1586(n20 ,n2404);
    not g1587(n19 ,n2400);
    not g1588(n18 ,n2403);
    not g1589(n17 ,n2399);
    not g1590(n16 ,n2406);
    not g1591(n15 ,n2405);
    not g1592(n14 ,n2402);
    xnor g1593(n2408 ,n63 ,n66);
    nor g1594(n2407 ,n63 ,n67);
    xor g1595(n2409 ,n2371 ,n64);
    not g1596(n67 ,n66);
    nor g1597(n66 ,n56 ,n65);
    not g1598(n65 ,n64);
    xnor g1599(n64 ,n2370 ,n61);
    nor g1600(n63 ,n60 ,n62);
    nor g1601(n62 ,n55 ,n59);
    xnor g1602(n61 ,n2373 ,n2372);
    nor g1603(n60 ,n57 ,n58);
    nor g1604(n59 ,n2373 ,n2370);
    not g1605(n58 ,n2370);
    not g1606(n57 ,n2373);
    not g1607(n56 ,n2371);
    not g1608(n55 ,n2372);
    or g1609(n2395 ,n466 ,n526);
    xnor g1610(n2394 ,n486 ,n525);
    nor g1611(n526 ,n474 ,n525);
    nor g1612(n525 ,n484 ,n524);
    xnor g1613(n2393 ,n494 ,n523);
    xnor g1614(n2392 ,n504 ,n522);
    nor g1615(n524 ,n490 ,n523);
    nor g1616(n523 ,n520 ,n515);
    nor g1617(n522 ,n496 ,n521);
    xnor g1618(n2391 ,n503 ,n518);
    nor g1619(n521 ,n500 ,n518);
    or g1620(n520 ,n492 ,n519);
    xnor g1621(n2390 ,n502 ,n514);
    nor g1622(n519 ,n505 ,n517);
    nor g1623(n518 ,n510 ,n516);
    not g1624(n517 ,n516);
    nor g1625(n516 ,n498 ,n512);
    or g1626(n515 ,n507 ,n513);
    nor g1627(n514 ,n487 ,n511);
    xnor g1628(n2389 ,n493 ,n508);
    nor g1629(n513 ,n505 ,n509);
    not g1630(n512 ,n511);
    nor g1631(n511 ,n489 ,n508);
    not g1632(n510 ,n509);
    nor g1633(n509 ,n495 ,n506);
    nor g1634(n508 ,n475 ,n501);
    xnor g1635(n2388 ,n485 ,n491);
    nor g1636(n507 ,n497 ,n499);
    nor g1637(n506 ,n488 ,n498);
    or g1638(n505 ,n500 ,n499);
    nor g1639(n504 ,n492 ,n499);
    nor g1640(n503 ,n496 ,n500);
    nor g1641(n502 ,n495 ,n498);
    nor g1642(n501 ,n476 ,n491);
    nor g1643(n500 ,n473 ,n483);
    nor g1644(n499 ,n468 ,n479);
    nor g1645(n498 ,n470 ,n481);
    not g1646(n497 ,n496);
    nor g1647(n496 ,n472 ,n482);
    nor g1648(n495 ,n469 ,n480);
    nor g1649(n494 ,n484 ,n490);
    nor g1650(n493 ,n487 ,n489);
    nor g1651(n492 ,n467 ,n478);
    nor g1652(n491 ,n460 ,n477);
    xnor g1653(n2387 ,n471 ,n461);
    not g1654(n488 ,n487);
    nor g1655(n486 ,n466 ,n474);
    nor g1656(n490 ,n447 ,n465);
    nor g1657(n489 ,n453 ,n463);
    nor g1658(n485 ,n475 ,n476);
    nor g1659(n487 ,n452 ,n462);
    not g1660(n483 ,n482);
    not g1661(n481 ,n480);
    not g1662(n479 ,n478);
    nor g1663(n477 ,n461 ,n459);
    xor g1664(n2386 ,n454 ,n379);
    nor g1665(n484 ,n446 ,n464);
    xnor g1666(n482 ,n443 ,n423);
    xnor g1667(n480 ,n444 ,n424);
    xnor g1668(n478 ,n442 ,n421);
    not g1669(n473 ,n472);
    nor g1670(n476 ,n431 ,n448);
    nor g1671(n475 ,n430 ,n449);
    nor g1672(n474 ,n385 ,n451);
    nor g1673(n472 ,n440 ,n456);
    nor g1674(n471 ,n460 ,n459);
    not g1675(n470 ,n469);
    not g1676(n468 ,n467);
    not g1677(n465 ,n464);
    not g1678(n463 ,n462);
    nor g1679(n469 ,n426 ,n458);
    nor g1680(n467 ,n428 ,n445);
    nor g1681(n466 ,n384 ,n450);
    nor g1682(n464 ,n429 ,n455);
    xnor g1683(n462 ,n425 ,n408);
    nor g1684(n461 ,n432 ,n457);
    nor g1685(n458 ,n395 ,n437);
    nor g1686(n457 ,n380 ,n441);
    nor g1687(n456 ,n424 ,n439);
    nor g1688(n455 ,n421 ,n438);
    nor g1689(n454 ,n432 ,n441);
    nor g1690(n460 ,n416 ,n434);
    nor g1691(n459 ,n417 ,n433);
    not g1692(n453 ,n452);
    not g1693(n451 ,n450);
    not g1694(n449 ,n448);
    not g1695(n447 ,n446);
    nor g1696(n445 ,n423 ,n436);
    xnor g1697(n444 ,n406 ,n393);
    nor g1698(n452 ,n418 ,n427);
    xnor g1699(n443 ,n410 ,n389);
    nor g1700(n450 ,n402 ,n435);
    xnor g1701(n448 ,n405 ,n391);
    xnor g1702(n446 ,n404 ,n422);
    xnor g1703(n442 ,n412 ,n387);
    nor g1704(n440 ,n393 ,n406);
    nor g1705(n439 ,n394 ,n407);
    nor g1706(n438 ,n388 ,n413);
    nor g1707(n437 ,n378 ,n409);
    nor g1708(n436 ,n390 ,n411);
    nor g1709(n435 ,n422 ,n397);
    nor g1710(n441 ,n361 ,n415);
    not g1711(n434 ,n433);
    not g1712(n431 ,n430);
    nor g1713(n429 ,n387 ,n412);
    nor g1714(n428 ,n389 ,n410);
    nor g1715(n427 ,n371 ,n419);
    nor g1716(n426 ,n377 ,n408);
    xnor g1717(n433 ,n386 ,n396);
    xor g1718(n425 ,n378 ,n395);
    nor g1719(n432 ,n360 ,n414);
    nor g1720(n430 ,n374 ,n420);
    nor g1721(n420 ,n373 ,n396);
    nor g1722(n419 ,n366 ,n392);
    nor g1723(n418 ,n367 ,n391);
    nor g1724(n424 ,n350 ,n401);
    nor g1725(n423 ,n339 ,n398);
    nor g1726(n422 ,n338 ,n399);
    nor g1727(n421 ,n349 ,n400);
    not g1728(n417 ,n416);
    not g1729(n415 ,n414);
    not g1730(n413 ,n412);
    not g1731(n411 ,n410);
    not g1732(n409 ,n408);
    not g1733(n407 ,n406);
    xnor g1734(n405 ,n366 ,n371);
    nor g1735(n416 ,n326 ,n403);
    xnor g1736(n414 ,n336 ,n372);
    xnor g1737(n404 ,n368 ,n375);
    xnor g1738(n412 ,n363 ,n382);
    xnor g1739(n410 ,n362 ,n381);
    xnor g1740(n408 ,n365 ,n383);
    xnor g1741(n406 ,n364 ,n370);
    nor g1742(n403 ,n300 ,n372);
    nor g1743(n402 ,n375 ,n368);
    nor g1744(n401 ,n359 ,n383);
    nor g1745(n400 ,n358 ,n381);
    nor g1746(n399 ,n357 ,n382);
    nor g1747(n398 ,n356 ,n370);
    nor g1748(n397 ,n376 ,n369);
    not g1749(n394 ,n393);
    not g1750(n392 ,n391);
    not g1751(n390 ,n389);
    not g1752(n388 ,n387);
    xor g1753(n2385 ,n275 ,n346);
    xnor g1754(n386 ,n342 ,n344);
    xnor g1755(n396 ,n331 ,n263);
    xnor g1756(n395 ,n334 ,n257);
    xnor g1757(n393 ,n337 ,n269);
    xnor g1758(n391 ,n332 ,n313);
    xnor g1759(n389 ,n333 ,n271);
    xnor g1760(n387 ,n335 ,n273);
    not g1761(n385 ,n384);
    not g1762(n380 ,n379);
    not g1763(n378 ,n377);
    not g1764(n376 ,n375);
    nor g1765(n374 ,n344 ,n343);
    nor g1766(n373 ,n345 ,n342);
    nor g1767(n384 ,n283 ,n341);
    nor g1768(n383 ,n324 ,n348);
    nor g1769(n382 ,n320 ,n353);
    nor g1770(n381 ,n328 ,n355);
    nor g1771(n379 ,n276 ,n347);
    nor g1772(n377 ,n321 ,n351);
    nor g1773(n375 ,n323 ,n354);
    not g1774(n369 ,n368);
    not g1775(n367 ,n366);
    xnor g1776(n365 ,n303 ,n243);
    xnor g1777(n364 ,n305 ,n311);
    xnor g1778(n363 ,n309 ,n329);
    xnor g1779(n362 ,n301 ,n307);
    xnor g1780(n372 ,n294 ,n235);
    nor g1781(n371 ,n327 ,n340);
    nor g1782(n370 ,n317 ,n352);
    xnor g1783(n368 ,n295 ,n314);
    xnor g1784(n366 ,n296 ,n290);
    not g1785(n361 ,n360);
    nor g1786(n359 ,n244 ,n304);
    nor g1787(n358 ,n308 ,n302);
    nor g1788(n357 ,n330 ,n310);
    nor g1789(n356 ,n312 ,n306);
    nor g1790(n355 ,n270 ,n319);
    nor g1791(n354 ,n274 ,n315);
    nor g1792(n353 ,n272 ,n316);
    nor g1793(n352 ,n277 ,n318);
    nor g1794(n351 ,n313 ,n297);
    nor g1795(n350 ,n243 ,n303);
    nor g1796(n349 ,n307 ,n301);
    nor g1797(n348 ,n250 ,n322);
    nor g1798(n360 ,n168 ,n325);
    not g1799(n347 ,n346);
    not g1800(n345 ,n344);
    not g1801(n343 ,n342);
    nor g1802(n341 ,n314 ,n287);
    nor g1803(n340 ,n247 ,n298);
    nor g1804(n339 ,n311 ,n305);
    nor g1805(n338 ,n329 ,n309);
    xnor g1806(n337 ,n259 ,n229);
    xnor g1807(n336 ,n253 ,n255);
    xnor g1808(n335 ,n265 ,n225);
    xor g1809(n334 ,n277 ,n241);
    xnor g1810(n333 ,n251 ,n233);
    xnor g1811(n332 ,n267 ,n288);
    xnor g1812(n331 ,n261 ,n247);
    xnor g1813(n346 ,n204 ,n292);
    nor g1814(n344 ,n279 ,n299);
    xnor g1815(n342 ,n278 ,n236);
    not g1816(n330 ,n329);
    nor g1817(n328 ,n229 ,n260);
    nor g1818(n327 ,n264 ,n262);
    nor g1819(n326 ,n254 ,n256);
    nor g1820(n325 ,n133 ,n293);
    nor g1821(n324 ,n245 ,n291);
    nor g1822(n323 ,n225 ,n266);
    nor g1823(n322 ,n246 ,n290);
    nor g1824(n321 ,n268 ,n289);
    nor g1825(n320 ,n233 ,n252);
    nor g1826(n319 ,n230 ,n259);
    nor g1827(n318 ,n242 ,n257);
    nor g1828(n317 ,n241 ,n258);
    nor g1829(n316 ,n234 ,n251);
    nor g1830(n315 ,n226 ,n265);
    nor g1831(n329 ,n171 ,n284);
    not g1832(n312 ,n311);
    not g1833(n310 ,n309);
    not g1834(n308 ,n307);
    not g1835(n306 ,n305);
    not g1836(n304 ,n303);
    not g1837(n302 ,n301);
    nor g1838(n300 ,n253 ,n255);
    nor g1839(n299 ,n235 ,n286);
    nor g1840(n298 ,n263 ,n261);
    nor g1841(n297 ,n267 ,n288);
    xnor g1842(n296 ,n245 ,n250);
    xnor g1843(n295 ,n223 ,n231);
    xnor g1844(n294 ,n201 ,n227);
    nor g1845(n314 ,n174 ,n281);
    nor g1846(n313 ,n239 ,n282);
    nor g1847(n311 ,n158 ,n280);
    xnor g1848(n309 ,n194 ,n238);
    nor g1849(n307 ,n170 ,n285);
    xnor g1850(n305 ,n192 ,n248);
    xnor g1851(n303 ,n191 ,n237);
    xnor g1852(n301 ,n196 ,n249);
    not g1853(n293 ,n292);
    not g1854(n291 ,n290);
    not g1855(n289 ,n288);
    nor g1856(n287 ,n232 ,n224);
    nor g1857(n286 ,n202 ,n228);
    nor g1858(n285 ,n149 ,n248);
    nor g1859(n284 ,n141 ,n249);
    nor g1860(n283 ,n231 ,n223);
    nor g1861(n282 ,n236 ,n240);
    nor g1862(n281 ,n152 ,n238);
    nor g1863(n280 ,n140 ,n237);
    nor g1864(n279 ,n201 ,n227);
    xnor g1865(n278 ,n199 ,n176);
    xnor g1866(n292 ,n0[32] ,n203);
    xnor g1867(n290 ,n197 ,n0[43]);
    xnor g1868(n288 ,n193 ,n178);
    not g1869(n276 ,n275);
    not g1870(n274 ,n273);
    not g1871(n272 ,n271);
    not g1872(n270 ,n269);
    not g1873(n268 ,n267);
    not g1874(n266 ,n265);
    not g1875(n264 ,n263);
    not g1876(n262 ,n261);
    not g1877(n260 ,n259);
    not g1878(n258 ,n257);
    not g1879(n256 ,n255);
    not g1880(n254 ,n253);
    not g1881(n252 ,n251);
    xor g1882(n277 ,n0[44] ,n198);
    xnor g1883(n275 ,n0[0] ,n184);
    xnor g1884(n273 ,n0[31] ,n205);
    xnor g1885(n271 ,n0[30] ,n188);
    xnor g1886(n269 ,n0[29] ,n190);
    xnor g1887(n267 ,n195 ,n0[27]);
    xnor g1888(n265 ,n187 ,n0[47]);
    xnor g1889(n263 ,n183 ,n0[2]);
    xnor g1890(n261 ,n182 ,n0[34]);
    xnor g1891(n259 ,n186 ,n0[45]);
    xnor g1892(n257 ,n181 ,n0[28]);
    xnor g1893(n255 ,n189 ,n0[33]);
    xnor g1894(n253 ,n185 ,n0[1]);
    xnor g1895(n251 ,n180 ,n0[46]);
    not g1896(n246 ,n245);
    not g1897(n244 ,n243);
    not g1898(n242 ,n241);
    nor g1899(n240 ,n176 ,n200);
    nor g1900(n239 ,n177 ,n199);
    nor g1901(n250 ,n157 ,n219);
    nor g1902(n249 ,n164 ,n218);
    nor g1903(n248 ,n172 ,n221);
    nor g1904(n247 ,n166 ,n212);
    nor g1905(n245 ,n167 ,n220);
    nor g1906(n243 ,n169 ,n206);
    nor g1907(n241 ,n160 ,n207);
    not g1908(n234 ,n233);
    not g1909(n232 ,n231);
    not g1910(n230 ,n229);
    not g1911(n228 ,n227);
    not g1912(n226 ,n225);
    not g1913(n224 ,n223);
    nor g1914(n238 ,n173 ,n208);
    nor g1915(n237 ,n161 ,n211);
    nor g1916(n236 ,n159 ,n214);
    nor g1917(n235 ,n155 ,n209);
    nor g1918(n233 ,n162 ,n213);
    nor g1919(n231 ,n132 ,n216);
    nor g1920(n229 ,n163 ,n222);
    nor g1921(n227 ,n156 ,n210);
    nor g1922(n225 ,n165 ,n215);
    nor g1923(n223 ,n175 ,n217);
    nor g1924(n222 ,n130 ,n143);
    nor g1925(n221 ,n93 ,n153);
    nor g1926(n220 ,n90 ,n135);
    nor g1927(n219 ,n88 ,n154);
    nor g1928(n218 ,n99 ,n142);
    nor g1929(n217 ,n124 ,n151);
    nor g1930(n216 ,n125 ,n145);
    nor g1931(n215 ,n98 ,n137);
    nor g1932(n214 ,n128 ,n139);
    nor g1933(n213 ,n129 ,n150);
    nor g1934(n212 ,n89 ,n136);
    nor g1935(n211 ,n94 ,n147);
    nor g1936(n210 ,n127 ,n148);
    nor g1937(n209 ,n126 ,n146);
    nor g1938(n208 ,n131 ,n144);
    nor g1939(n207 ,n92 ,n134);
    nor g1940(n206 ,n179 ,n138);
    xnor g1941(n205 ,n0[39] ,n0[15]);
    xnor g1942(n204 ,n0[24] ,n0[40]);
    xnor g1943(n203 ,n0[48] ,n0[16]);
    not g1944(n202 ,n201);
    not g1945(n200 ,n199);
    xnor g1946(n198 ,n0[60] ,n0[52]);
    xnor g1947(n197 ,n0[59] ,n0[51]);
    xnor g1948(n196 ,n0[22] ,n0[6]);
    xnor g1949(n195 ,n0[35] ,n0[11]);
    xnor g1950(n194 ,n0[23] ,n0[7]);
    xnor g1951(n193 ,n0[19] ,n0[3]);
    xnor g1952(n192 ,n0[21] ,n0[5]);
    xnor g1953(n191 ,n0[20] ,n0[4]);
    xnor g1954(n190 ,n0[37] ,n0[13]);
    xnor g1955(n189 ,n0[41] ,n0[9]);
    xnor g1956(n188 ,n0[38] ,n0[14]);
    xnor g1957(n187 ,n0[63] ,n0[55]);
    xnor g1958(n186 ,n0[61] ,n0[53]);
    xnor g1959(n185 ,n0[25] ,n0[17]);
    xnor g1960(n184 ,n0[56] ,n0[8]);
    xnor g1961(n183 ,n0[26] ,n0[18]);
    xnor g1962(n182 ,n0[42] ,n0[10]);
    xnor g1963(n181 ,n0[36] ,n0[12]);
    xnor g1964(n180 ,n0[62] ,n0[54]);
    xnor g1965(n201 ,n0[57] ,n0[49]);
    xnor g1966(n199 ,n0[58] ,n0[50]);
    not g1967(n179 ,n178);
    not g1968(n177 ,n176);
    nor g1969(n175 ,n115 ,n120);
    nor g1970(n174 ,n73 ,n102);
    nor g1971(n173 ,n70 ,n84);
    nor g1972(n172 ,n111 ,n105);
    nor g1973(n171 ,n118 ,n109);
    nor g1974(n170 ,n121 ,n123);
    nor g1975(n169 ,n107 ,n103);
    nor g1976(n168 ,n104 ,n122);
    nor g1977(n167 ,n100 ,n85);
    nor g1978(n166 ,n86 ,n77);
    nor g1979(n165 ,n71 ,n76);
    nor g1980(n164 ,n74 ,n119);
    nor g1981(n163 ,n78 ,n82);
    nor g1982(n162 ,n117 ,n83);
    nor g1983(n161 ,n113 ,n101);
    nor g1984(n160 ,n108 ,n110);
    nor g1985(n159 ,n69 ,n72);
    nor g1986(n158 ,n79 ,n68);
    nor g1987(n157 ,n80 ,n116);
    nor g1988(n156 ,n81 ,n112);
    nor g1989(n155 ,n75 ,n114);
    nor g1990(n178 ,n95 ,n91);
    nor g1991(n176 ,n96 ,n97);
    nor g1992(n154 ,n0[26] ,n0[18]);
    nor g1993(n153 ,n0[60] ,n0[44]);
    nor g1994(n152 ,n0[23] ,n0[7]);
    nor g1995(n151 ,n0[39] ,n0[15]);
    nor g1996(n150 ,n0[29] ,n0[13]);
    nor g1997(n149 ,n0[21] ,n0[5]);
    nor g1998(n148 ,n0[48] ,n0[16]);
    nor g1999(n147 ,n0[59] ,n0[43]);
    nor g2000(n146 ,n0[56] ,n0[8]);
    nor g2001(n145 ,n0[63] ,n0[47]);
    nor g2002(n144 ,n0[62] ,n0[46]);
    nor g2003(n143 ,n0[28] ,n0[12]);
    nor g2004(n142 ,n0[61] ,n0[45]);
    nor g2005(n141 ,n0[22] ,n0[6]);
    nor g2006(n140 ,n0[20] ,n0[4]);
    nor g2007(n139 ,n0[25] ,n0[1]);
    nor g2008(n138 ,n0[19] ,n0[3]);
    nor g2009(n137 ,n0[30] ,n0[14]);
    nor g2010(n136 ,n0[33] ,n0[9]);
    nor g2011(n135 ,n0[42] ,n0[10]);
    nor g2012(n134 ,n0[27] ,n0[11]);
    nor g2013(n133 ,n0[24] ,n0[40]);
    nor g2014(n132 ,n106 ,n87);
    not g2015(n131 ,n0[54]);
    not g2016(n130 ,n0[36]);
    not g2017(n129 ,n0[37]);
    not g2018(n128 ,n0[17]);
    not g2019(n127 ,n0[32]);
    not g2020(n126 ,n0[0]);
    not g2021(n125 ,n0[55]);
    not g2022(n124 ,n0[31]);
    not g2023(n123 ,n0[5]);
    not g2024(n122 ,n0[40]);
    not g2025(n121 ,n0[21]);
    not g2026(n120 ,n0[15]);
    not g2027(n119 ,n0[45]);
    not g2028(n118 ,n0[22]);
    not g2029(n117 ,n0[29]);
    not g2030(n116 ,n0[18]);
    not g2031(n115 ,n0[39]);
    not g2032(n114 ,n0[8]);
    not g2033(n113 ,n0[59]);
    not g2034(n112 ,n0[16]);
    not g2035(n111 ,n0[60]);
    not g2036(n110 ,n0[11]);
    not g2037(n109 ,n0[6]);
    not g2038(n108 ,n0[27]);
    not g2039(n107 ,n0[19]);
    not g2040(n106 ,n0[63]);
    not g2041(n105 ,n0[44]);
    not g2042(n104 ,n0[24]);
    not g2043(n103 ,n0[3]);
    not g2044(n102 ,n0[7]);
    not g2045(n101 ,n0[43]);
    not g2046(n100 ,n0[42]);
    not g2047(n99 ,n0[53]);
    not g2048(n98 ,n0[38]);
    not g2049(n97 ,n0[49]);
    not g2050(n96 ,n0[57]);
    not g2051(n95 ,n0[58]);
    not g2052(n94 ,n0[51]);
    not g2053(n93 ,n0[52]);
    not g2054(n92 ,n0[35]);
    not g2055(n91 ,n0[50]);
    not g2056(n90 ,n0[34]);
    not g2057(n89 ,n0[41]);
    not g2058(n88 ,n0[2]);
    not g2059(n87 ,n0[47]);
    not g2060(n86 ,n0[33]);
    not g2061(n85 ,n0[10]);
    not g2062(n84 ,n0[46]);
    not g2063(n83 ,n0[13]);
    not g2064(n82 ,n0[12]);
    not g2065(n81 ,n0[48]);
    not g2066(n80 ,n0[26]);
    not g2067(n79 ,n0[20]);
    not g2068(n78 ,n0[28]);
    not g2069(n77 ,n0[9]);
    not g2070(n76 ,n0[14]);
    not g2071(n75 ,n0[56]);
    not g2072(n74 ,n0[61]);
    not g2073(n73 ,n0[23]);
    not g2074(n72 ,n0[1]);
    not g2075(n71 ,n0[30]);
    not g2076(n70 ,n0[62]);
    not g2077(n69 ,n0[25]);
    not g2078(n68 ,n0[4]);
    xnor g2079(n2383 ,n1018 ,n981);
    nor g2080(n2384 ,n982 ,n1018);
    nor g2081(n1018 ,n1017 ,n1009);
    xnor g2082(n2382 ,n1014 ,n1016);
    nor g2083(n1017 ,n1008 ,n1016);
    nor g2084(n1016 ,n1015 ,n1011);
    xnor g2085(n2381 ,n1013 ,n1012);
    nor g2086(n1015 ,n1012 ,n1010);
    xnor g2087(n2380 ,n1006 ,n999);
    nor g2088(n1014 ,n1009 ,n1008);
    nor g2089(n1013 ,n1011 ,n1010);
    nor g2090(n1012 ,n1004 ,n1007);
    nor g2091(n1011 ,n997 ,n1001);
    nor g2092(n1010 ,n998 ,n1000);
    nor g2093(n1009 ,n987 ,n1002);
    nor g2094(n1008 ,n986 ,n1003);
    nor g2095(n1007 ,n999 ,n1005);
    nor g2096(n1006 ,n1004 ,n1005);
    nor g2097(n1005 ,n994 ,n993);
    nor g2098(n1004 ,n995 ,n992);
    not g2099(n1003 ,n1002);
    nor g2100(n1002 ,n979 ,n996);
    not g2101(n1001 ,n1000);
    xnor g2102(n1000 ,n985 ,n988);
    xnor g2103(n2379 ,n989 ,n969);
    nor g2104(n999 ,n983 ,n991);
    not g2105(n998 ,n997);
    nor g2106(n997 ,n968 ,n990);
    nor g2107(n996 ,n977 ,n988);
    not g2108(n995 ,n994);
    xnor g2109(n994 ,n974 ,n955);
    not g2110(n993 ,n992);
    xnor g2111(n992 ,n975 ,n978);
    nor g2112(n991 ,n969 ,n984);
    nor g2113(n990 ,n973 ,n978);
    nor g2114(n989 ,n983 ,n984);
    nor g2115(n988 ,n972 ,n976);
    not g2116(n987 ,n986);
    nor g2117(n986 ,n981 ,n980);
    xnor g2118(n985 ,n960 ,n945);
    not g2119(n982 ,n981);
    nor g2120(n980 ,n905 ,n967);
    nor g2121(n979 ,n945 ,n961);
    nor g2122(n984 ,n965 ,n962);
    nor g2123(n983 ,n964 ,n963);
    nor g2124(n981 ,n906 ,n966);
    nor g2125(n977 ,n946 ,n960);
    nor g2126(n976 ,n955 ,n971);
    xor g2127(n2378 ,n952 ,n846);
    xnor g2128(n975 ,n953 ,n947);
    xnor g2129(n974 ,n895 ,n950);
    nor g2130(n978 ,n958 ,n970);
    nor g2131(n973 ,n948 ,n954);
    nor g2132(n972 ,n896 ,n950);
    nor g2133(n971 ,n895 ,n951);
    nor g2134(n970 ,n924 ,n959);
    nor g2135(n969 ,n949 ,n957);
    nor g2136(n968 ,n947 ,n953);
    not g2137(n967 ,n966);
    nor g2138(n966 ,n936 ,n956);
    not g2139(n965 ,n964);
    xnor g2140(n964 ,n941 ,n917);
    not g2141(n963 ,n962);
    xnor g2142(n962 ,n940 ,n937);
    not g2143(n961 ,n960);
    xnor g2144(n960 ,n939 ,n943);
    nor g2145(n959 ,n923 ,n937);
    nor g2146(n958 ,n922 ,n938);
    nor g2147(n957 ,n931 ,n944);
    nor g2148(n956 ,n935 ,n943);
    nor g2149(n955 ,n928 ,n942);
    not g2150(n954 ,n953);
    xnor g2151(n953 ,n925 ,n904);
    xnor g2152(n952 ,n929 ,n931);
    not g2153(n951 ,n950);
    xnor g2154(n950 ,n926 ,n897);
    nor g2155(n949 ,n847 ,n930);
    not g2156(n948 ,n947);
    nor g2157(n947 ,n898 ,n933);
    not g2158(n946 ,n945);
    nor g2159(n945 ,n918 ,n932);
    nor g2160(n944 ,n846 ,n929);
    nor g2161(n943 ,n919 ,n927);
    nor g2162(n942 ,n917 ,n934);
    xnor g2163(n941 ,n914 ,n908);
    xnor g2164(n940 ,n924 ,n922);
    xnor g2165(n939 ,n912 ,n910);
    not g2166(n938 ,n937);
    xnor g2167(n937 ,n907 ,n916);
    nor g2168(n936 ,n910 ,n913);
    nor g2169(n935 ,n911 ,n912);
    nor g2170(n934 ,n909 ,n915);
    nor g2171(n933 ,n900 ,n916);
    nor g2172(n932 ,n904 ,n920);
    not g2173(n930 ,n929);
    nor g2174(n928 ,n908 ,n914);
    nor g2175(n927 ,n897 ,n921);
    xnor g2176(n926 ,n893 ,n891);
    xnor g2177(n925 ,n902 ,n869);
    xnor g2178(n931 ,n889 ,n854);
    xnor g2179(n929 ,n888 ,n848);
    not g2180(n923 ,n922);
    nor g2181(n921 ,n894 ,n892);
    nor g2182(n920 ,n870 ,n903);
    nor g2183(n919 ,n893 ,n891);
    nor g2184(n918 ,n869 ,n902);
    nor g2185(n924 ,n882 ,n901);
    nor g2186(n922 ,n885 ,n899);
    not g2187(n915 ,n914);
    not g2188(n913 ,n912);
    not g2189(n911 ,n910);
    not g2190(n909 ,n908);
    xnor g2191(n907 ,n878 ,n831);
    xnor g2192(n917 ,n874 ,n821);
    xnor g2193(n916 ,n873 ,n827);
    xnor g2194(n914 ,n871 ,n823);
    xnor g2195(n912 ,n887 ,n841);
    nor g2196(n910 ,n883 ,n890);
    xnor g2197(n908 ,n872 ,n838);
    not g2198(n906 ,n905);
    not g2199(n903 ,n902);
    nor g2200(n901 ,n858 ,n886);
    nor g2201(n900 ,n832 ,n878);
    nor g2202(n899 ,n859 ,n876);
    nor g2203(n898 ,n831 ,n879);
    nor g2204(n905 ,n842 ,n887);
    nor g2205(n904 ,n861 ,n875);
    nor g2206(n902 ,n863 ,n880);
    not g2207(n896 ,n895);
    not g2208(n894 ,n893);
    not g2209(n892 ,n891);
    nor g2210(n890 ,n802 ,n884);
    xnor g2211(n889 ,n852 ,n858);
    xor g2212(n888 ,n859 ,n850);
    nor g2213(n897 ,n864 ,n881);
    xnor g2214(n895 ,n845 ,n856);
    xnor g2215(n893 ,n844 ,n803);
    nor g2216(n891 ,n860 ,n877);
    nor g2217(n886 ,n852 ,n854);
    nor g2218(n885 ,n851 ,n849);
    nor g2219(n884 ,n799 ,n856);
    nor g2220(n883 ,n798 ,n857);
    nor g2221(n882 ,n853 ,n855);
    nor g2222(n881 ,n838 ,n868);
    nor g2223(n880 ,n843 ,n867);
    nor g2224(n887 ,n833 ,n862);
    not g2225(n879 ,n878);
    nor g2226(n877 ,n839 ,n865);
    nor g2227(n876 ,n850 ,n848);
    nor g2228(n875 ,n840 ,n866);
    xnor g2229(n874 ,n819 ,n839);
    xnor g2230(n873 ,n825 ,n843);
    xnor g2231(n872 ,n829 ,n817);
    xnor g2232(n871 ,n836 ,n840);
    xnor g2233(n878 ,n816 ,n759);
    not g2234(n870 ,n869);
    nor g2235(n868 ,n830 ,n818);
    nor g2236(n867 ,n826 ,n828);
    nor g2237(n866 ,n824 ,n837);
    nor g2238(n865 ,n822 ,n820);
    nor g2239(n864 ,n829 ,n817);
    nor g2240(n863 ,n825 ,n827);
    nor g2241(n862 ,n803 ,n834);
    nor g2242(n861 ,n823 ,n836);
    nor g2243(n860 ,n821 ,n819);
    nor g2244(n869 ,n810 ,n835);
    not g2245(n857 ,n856);
    not g2246(n855 ,n854);
    not g2247(n853 ,n852);
    not g2248(n851 ,n850);
    not g2249(n849 ,n848);
    not g2250(n847 ,n846);
    xnor g2251(n845 ,n798 ,n802);
    xnor g2252(n844 ,n813 ,n800);
    xor g2253(n859 ,n796 ,n739);
    xnor g2254(n858 ,n797 ,n755);
    xnor g2255(n856 ,n815 ,n760);
    xnor g2256(n854 ,n793 ,n713);
    xnor g2257(n852 ,n792 ,n717);
    xnor g2258(n850 ,n794 ,n721);
    xnor g2259(n848 ,n795 ,n735);
    xnor g2260(n846 ,n791 ,n757);
    not g2261(n842 ,n841);
    not g2262(n837 ,n836);
    nor g2263(n835 ,n759 ,n809);
    nor g2264(n834 ,n801 ,n814);
    nor g2265(n833 ,n800 ,n813);
    nor g2266(n843 ,n789 ,n808);
    nor g2267(n841 ,n761 ,n815);
    nor g2268(n840 ,n787 ,n806);
    nor g2269(n839 ,n786 ,n805);
    nor g2270(n838 ,n790 ,n811);
    nor g2271(n836 ,n788 ,n812);
    not g2272(n832 ,n831);
    not g2273(n830 ,n829);
    not g2274(n828 ,n827);
    not g2275(n826 ,n825);
    not g2276(n824 ,n823);
    not g2277(n822 ,n821);
    not g2278(n820 ,n819);
    not g2279(n818 ,n817);
    xnor g2280(n816 ,n776 ,n706);
    nor g2281(n831 ,n783 ,n807);
    xnor g2282(n829 ,n763 ,n694);
    xnor g2283(n827 ,n767 ,n709);
    xnor g2284(n825 ,n768 ,n704);
    xnor g2285(n823 ,n766 ,n710);
    xnor g2286(n821 ,n765 ,n691);
    xnor g2287(n819 ,n764 ,n692);
    nor g2288(n817 ,n785 ,n804);
    not g2289(n814 ,n813);
    nor g2290(n812 ,n736 ,n774);
    nor g2291(n811 ,n737 ,n781);
    nor g2292(n810 ,n706 ,n777);
    nor g2293(n809 ,n707 ,n776);
    nor g2294(n808 ,n738 ,n769);
    nor g2295(n807 ,n762 ,n784);
    nor g2296(n806 ,n742 ,n772);
    nor g2297(n805 ,n740 ,n770);
    nor g2298(n804 ,n741 ,n782);
    nor g2299(n815 ,n747 ,n779);
    nor g2300(n813 ,n746 ,n778);
    not g2301(n801 ,n800);
    not g2302(n799 ,n798);
    xor g2303(n797 ,n762 ,n715);
    xnor g2304(n796 ,n725 ,n723);
    xnor g2305(n795 ,n719 ,n727);
    xor g2306(n794 ,n742 ,n731);
    xor g2307(n793 ,n738 ,n711);
    xor g2308(n792 ,n741 ,n733);
    xor g2309(n791 ,n737 ,n729);
    nor g2310(n803 ,n743 ,n773);
    nor g2311(n802 ,n745 ,n775);
    nor g2312(n800 ,n744 ,n771);
    nor g2313(n798 ,n748 ,n780);
    nor g2314(n790 ,n758 ,n730);
    nor g2315(n789 ,n712 ,n714);
    nor g2316(n788 ,n720 ,n728);
    nor g2317(n787 ,n722 ,n732);
    nor g2318(n786 ,n726 ,n724);
    nor g2319(n785 ,n734 ,n718);
    nor g2320(n784 ,n715 ,n756);
    nor g2321(n783 ,n716 ,n755);
    nor g2322(n782 ,n733 ,n717);
    nor g2323(n781 ,n757 ,n729);
    nor g2324(n780 ,n710 ,n754);
    nor g2325(n779 ,n692 ,n753);
    nor g2326(n778 ,n709 ,n751);
    not g2327(n777 ,n776);
    nor g2328(n775 ,n693 ,n752);
    nor g2329(n774 ,n719 ,n727);
    nor g2330(n773 ,n694 ,n749);
    nor g2331(n772 ,n721 ,n731);
    nor g2332(n771 ,n691 ,n750);
    nor g2333(n770 ,n725 ,n723);
    nor g2334(n769 ,n711 ,n713);
    xnor g2335(n768 ,n702 ,n693);
    xnor g2336(n767 ,n677 ,n696);
    xnor g2337(n766 ,n681 ,n700);
    xnor g2338(n765 ,n685 ,n683);
    xnor g2339(n764 ,n687 ,n698);
    xnor g2340(n763 ,n689 ,n679);
    xnor g2341(n776 ,n633 ,n708);
    not g2342(n761 ,n760);
    not g2343(n758 ,n757);
    not g2344(n756 ,n755);
    nor g2345(n754 ,n701 ,n682);
    nor g2346(n753 ,n699 ,n688);
    nor g2347(n752 ,n705 ,n703);
    nor g2348(n751 ,n697 ,n678);
    nor g2349(n750 ,n684 ,n686);
    nor g2350(n749 ,n680 ,n690);
    nor g2351(n748 ,n700 ,n681);
    nor g2352(n747 ,n698 ,n687);
    nor g2353(n746 ,n696 ,n677);
    nor g2354(n745 ,n704 ,n702);
    nor g2355(n744 ,n683 ,n685);
    nor g2356(n743 ,n679 ,n689);
    xor g2357(n762 ,n2435 ,n650);
    nor g2358(n760 ,n634 ,n708);
    nor g2359(n759 ,n624 ,n695);
    xnor g2360(n757 ,n2489 ,n656);
    xnor g2361(n755 ,n645 ,n655);
    not g2362(n740 ,n739);
    not g2363(n736 ,n735);
    not g2364(n734 ,n733);
    not g2365(n732 ,n731);
    not g2366(n730 ,n729);
    not g2367(n728 ,n727);
    not g2368(n726 ,n725);
    not g2369(n724 ,n723);
    not g2370(n722 ,n721);
    not g2371(n720 ,n719);
    not g2372(n718 ,n717);
    not g2373(n716 ,n715);
    not g2374(n714 ,n713);
    not g2375(n712 ,n711);
    xor g2376(n742 ,n2461 ,n652);
    xor g2377(n741 ,n2486 ,n653);
    xnor g2378(n739 ,n2473 ,n637);
    xor g2379(n738 ,n2456 ,n648);
    xor g2380(n737 ,n2450 ,n644);
    xnor g2381(n735 ,n2468 ,n643);
    xnor g2382(n733 ,n2430 ,n646);
    xnor g2383(n731 ,n2445 ,n636);
    xnor g2384(n729 ,n2443 ,n651);
    xnor g2385(n727 ,n2439 ,n647);
    xnor g2386(n725 ,n2459 ,n638);
    xnor g2387(n723 ,n2441 ,n639);
    xnor g2388(n721 ,n2452 ,n640);
    xnor g2389(n719 ,n2470 ,n641);
    xnor g2390(n717 ,n2454 ,n635);
    xnor g2391(n715 ,n2487 ,n654);
    xnor g2392(n713 ,n2447 ,n642);
    xnor g2393(n711 ,n2448 ,n649);
    not g2394(n707 ,n706);
    not g2395(n705 ,n704);
    not g2396(n703 ,n702);
    not g2397(n701 ,n700);
    not g2398(n699 ,n698);
    not g2399(n697 ,n696);
    nor g2400(n695 ,n602 ,n655);
    nor g2401(n710 ,n629 ,n674);
    nor g2402(n709 ,n619 ,n666);
    nor g2403(n708 ,n621 ,n665);
    nor g2404(n706 ,n613 ,n675);
    nor g2405(n704 ,n614 ,n670);
    nor g2406(n702 ,n622 ,n668);
    nor g2407(n700 ,n620 ,n671);
    nor g2408(n698 ,n618 ,n676);
    nor g2409(n696 ,n627 ,n660);
    not g2410(n690 ,n689);
    not g2411(n688 ,n687);
    not g2412(n686 ,n685);
    not g2413(n684 ,n683);
    not g2414(n682 ,n681);
    not g2415(n680 ,n679);
    not g2416(n678 ,n677);
    nor g2417(n694 ,n625 ,n661);
    nor g2418(n693 ,n630 ,n662);
    nor g2419(n692 ,n626 ,n672);
    nor g2420(n691 ,n628 ,n657);
    nor g2421(n689 ,n632 ,n658);
    nor g2422(n687 ,n601 ,n659);
    nor g2423(n685 ,n616 ,n673);
    nor g2424(n683 ,n615 ,n664);
    nor g2425(n681 ,n631 ,n667);
    nor g2426(n679 ,n617 ,n663);
    nor g2427(n677 ,n623 ,n669);
    nor g2428(n676 ,n588 ,n599);
    nor g2429(n675 ,n552 ,n603);
    nor g2430(n674 ,n590 ,n592);
    nor g2431(n673 ,n557 ,n597);
    nor g2432(n672 ,n556 ,n591);
    nor g2433(n671 ,n586 ,n594);
    nor g2434(n670 ,n553 ,n600);
    nor g2435(n669 ,n551 ,n593);
    nor g2436(n668 ,n548 ,n612);
    nor g2437(n667 ,n583 ,n609);
    nor g2438(n666 ,n587 ,n608);
    nor g2439(n665 ,n580 ,n610);
    nor g2440(n664 ,n582 ,n595);
    nor g2441(n663 ,n555 ,n598);
    nor g2442(n662 ,n584 ,n605);
    nor g2443(n661 ,n549 ,n611);
    nor g2444(n660 ,n581 ,n596);
    nor g2445(n659 ,n589 ,n606);
    nor g2446(n658 ,n558 ,n607);
    nor g2447(n657 ,n554 ,n604);
    xnor g2448(n656 ,n2484 ,n2472);
    xnor g2449(n654 ,n2491 ,n2460);
    xnor g2450(n653 ,n2432 ,n2477);
    xnor g2451(n652 ,n2478 ,n2462);
    xnor g2452(n651 ,n2488 ,n2442);
    xnor g2453(n650 ,n2476 ,n2475);
    xnor g2454(n649 ,n2466 ,n2429);
    xnor g2455(n648 ,n2455 ,n2433);
    xnor g2456(n647 ,n2436 ,n2492);
    xnor g2457(n646 ,n2479 ,n2457);
    xnor g2458(n645 ,n2483 ,n2482);
    xnor g2459(n644 ,n2480 ,n2449);
    xnor g2460(n643 ,n2490 ,n2431);
    xnor g2461(n642 ,n2467 ,n2446);
    xnor g2462(n641 ,n2485 ,n2469);
    xnor g2463(n640 ,n2465 ,n2451);
    xnor g2464(n639 ,n2440 ,n2434);
    xnor g2465(n638 ,n2463 ,n2458);
    xnor g2466(n637 ,n2474 ,n2471);
    xnor g2467(n636 ,n2481 ,n2444);
    xnor g2468(n635 ,n2464 ,n2453);
    xnor g2469(n655 ,n2437 ,n2438);
    not g2470(n634 ,n633);
    nor g2471(n632 ,n529 ,n544);
    nor g2472(n631 ,n563 ,n575);
    nor g2473(n630 ,n569 ,n534);
    nor g2474(n629 ,n565 ,n570);
    nor g2475(n628 ,n567 ,n543);
    nor g2476(n627 ,n559 ,n566);
    nor g2477(n626 ,n533 ,n577);
    nor g2478(n625 ,n545 ,n564);
    nor g2479(n624 ,n578 ,n546);
    nor g2480(n623 ,n568 ,n561);
    nor g2481(n622 ,n535 ,n572);
    nor g2482(n621 ,n531 ,n560);
    nor g2483(n620 ,n539 ,n573);
    nor g2484(n619 ,n530 ,n532);
    nor g2485(n618 ,n541 ,n574);
    nor g2486(n617 ,n547 ,n537);
    nor g2487(n616 ,n576 ,n571);
    nor g2488(n615 ,n536 ,n538);
    nor g2489(n614 ,n528 ,n579);
    nor g2490(n613 ,n527 ,n562);
    nor g2491(n633 ,n585 ,n550);
    nor g2492(n612 ,n2466 ,n2448);
    nor g2493(n611 ,n2490 ,n2468);
    nor g2494(n610 ,n2436 ,n2439);
    nor g2495(n609 ,n2434 ,n2441);
    nor g2496(n608 ,n2464 ,n2454);
    nor g2497(n607 ,n2465 ,n2452);
    nor g2498(n606 ,n2488 ,n2443);
    nor g2499(n605 ,n2463 ,n2459);
    nor g2500(n604 ,n2433 ,n2456);
    nor g2501(n603 ,n2491 ,n2487);
    nor g2502(n602 ,n2483 ,n2482);
    nor g2503(n601 ,n542 ,n540);
    nor g2504(n600 ,n2478 ,n2462);
    nor g2505(n599 ,n2480 ,n2450);
    nor g2506(n598 ,n2435 ,n2476);
    nor g2507(n597 ,n2474 ,n2473);
    nor g2508(n596 ,n2485 ,n2470);
    nor g2509(n595 ,n2489 ,n2484);
    nor g2510(n594 ,n2467 ,n2447);
    nor g2511(n593 ,n2481 ,n2445);
    nor g2512(n592 ,n2479 ,n2430);
    nor g2513(n591 ,n2486 ,n2432);
    not g2514(n590 ,n2457);
    not g2515(n589 ,n2442);
    not g2516(n588 ,n2449);
    not g2517(n587 ,n2453);
    not g2518(n586 ,n2446);
    not g2519(n585 ,n2437);
    not g2520(n584 ,n2458);
    not g2521(n583 ,n2440);
    not g2522(n582 ,n2472);
    not g2523(n581 ,n2469);
    not g2524(n580 ,n2492);
    not g2525(n579 ,n2462);
    not g2526(n578 ,n2483);
    not g2527(n577 ,n2432);
    not g2528(n576 ,n2474);
    not g2529(n575 ,n2441);
    not g2530(n574 ,n2450);
    not g2531(n573 ,n2447);
    not g2532(n572 ,n2448);
    not g2533(n571 ,n2473);
    not g2534(n570 ,n2430);
    not g2535(n569 ,n2463);
    not g2536(n568 ,n2481);
    not g2537(n567 ,n2433);
    not g2538(n566 ,n2470);
    not g2539(n565 ,n2479);
    not g2540(n564 ,n2468);
    not g2541(n563 ,n2434);
    not g2542(n562 ,n2487);
    not g2543(n561 ,n2445);
    not g2544(n560 ,n2439);
    not g2545(n559 ,n2485);
    not g2546(n558 ,n2451);
    not g2547(n557 ,n2471);
    not g2548(n556 ,n2477);
    not g2549(n555 ,n2475);
    not g2550(n554 ,n2455);
    not g2551(n553 ,n2461);
    not g2552(n552 ,n2460);
    not g2553(n551 ,n2444);
    not g2554(n550 ,n2438);
    not g2555(n549 ,n2431);
    not g2556(n548 ,n2429);
    not g2557(n547 ,n2435);
    not g2558(n546 ,n2482);
    not g2559(n545 ,n2490);
    not g2560(n544 ,n2452);
    not g2561(n543 ,n2456);
    not g2562(n542 ,n2488);
    not g2563(n541 ,n2480);
    not g2564(n540 ,n2443);
    not g2565(n539 ,n2467);
    not g2566(n538 ,n2484);
    not g2567(n537 ,n2476);
    not g2568(n536 ,n2489);
    not g2569(n535 ,n2466);
    not g2570(n534 ,n2459);
    not g2571(n533 ,n2486);
    not g2572(n532 ,n2454);
    not g2573(n531 ,n2436);
    not g2574(n530 ,n2464);
    not g2575(n529 ,n2465);
    not g2576(n528 ,n2478);
    not g2577(n527 ,n2491);
    or g2578(n2428 ,n1022 ,n1021);
    nor g2579(n1022 ,n1019 ,n1020);
    or g2580(n1021 ,n2412 ,n2398);
    not g2581(n1020 ,n2414);
    not g2582(n1019 ,n2413);
    or g2583(n2427 ,n2407 ,n1025);
    nor g2584(n1025 ,n1023 ,n1024);
    not g2585(n1024 ,n2409);
    not g2586(n1023 ,n2408);
    nor g2587(n2421 ,n2417 ,n2525);
    nor g2588(n2419 ,n2526 ,n2527);
    nor g2589(n2422 ,n2503 ,n2523);
    nor g2590(n2527 ,n2502 ,n2524);
    nor g2591(n2417 ,n5[2] ,n2521);
    nor g2592(n2526 ,n5[0] ,n2522);
    nor g2593(n2525 ,n2516 ,n2520);
    nor g2594(n2524 ,n2509 ,n2514);
    nor g2595(n2418 ,n2519 ,n2514);
    or g2596(n2420 ,n2516 ,n2515);
    or g2597(n2523 ,n2505 ,n2519);
    or g2598(n2522 ,n2510 ,n2516);
    not g2599(n2521 ,n2520);
    nor g2600(n2520 ,n2518 ,n2517);
    nor g2601(n2519 ,n2501 ,n2507);
    nor g2602(n2518 ,n2502 ,n2512);
    nor g2603(n2416 ,n2506 ,n2508);
    nor g2604(n2517 ,n5[0] ,n2504);
    nor g2605(n2415 ,n5[0] ,n2508);
    nor g2606(n2516 ,n5[2] ,n2513);
    nor g2607(n2515 ,n2511 ,n2506);
    or g2608(n2514 ,n5[2] ,n2505);
    or g2609(n2513 ,n2500 ,n2501);
    nor g2610(n2512 ,n2499 ,n5[1]);
    not g2611(n2511 ,n2510);
    nor g2612(n2510 ,n2503 ,n5[1]);
    nor g2613(n2509 ,n2501 ,n2423);
    or g2614(n2508 ,n5[2] ,n5[1]);
    not g2615(n2507 ,n2506);
    nor g2616(n2506 ,n2423 ,n5[0]);
    not g2617(n2504 ,n2505);
    nor g2618(n2505 ,n2424 ,n5[1]);
    not g2619(n2503 ,n5[2]);
    not g2620(n2502 ,n5[0]);
    not g2621(n2501 ,n5[1]);
    not g2622(n2500 ,n2424);
    not g2623(n2499 ,n2423);
    buf g2624(n1823 ,n1768);
    buf g2625(n2365 ,n2375);
    not g2626(n1189 ,n2408);
    buf g2627(n2297 ,n2398);
endmodule
