module top(n0, n1, n2);
    input n0, n1;
    output n2;
    wire n0, n1;
    wire n2;
    wire [31:0] n3;
    wire [31:0] n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798;
    buf g0(n4[31], 1'b0);
    buf g1(n4[30], 1'b0);
    buf g2(n4[29], 1'b0);
    buf g3(n4[28], 1'b0);
    buf g4(n4[27], 1'b0);
    buf g5(n4[26], 1'b0);
    buf g6(n4[25], 1'b0);
    buf g7(n4[24], 1'b0);
    buf g8(n4[23], 1'b0);
    buf g9(n4[22], 1'b0);
    buf g10(n4[21], 1'b0);
    buf g11(n4[20], 1'b0);
    buf g12(n4[19], 1'b0);
    buf g13(n4[18], 1'b0);
    buf g14(n4[17], 1'b0);
    buf g15(n4[16], 1'b0);
    buf g16(n4[15], 1'b0);
    buf g17(n4[14], 1'b0);
    buf g18(n4[13], 1'b0);
    buf g19(n4[12], 1'b0);
    buf g20(n4[11], 1'b0);
    buf g21(n4[10], 1'b0);
    buf g22(n4[9], 1'b0);
    buf g23(n4[8], 1'b0);
    buf g24(n4[7], 1'b0);
    buf g25(n4[6], 1'b0);
    buf g26(n4[5], 1'b0);
    buf g27(n4[4], 1'b0);
    buf g28(n4[3], 1'b0);
    buf g29(n4[2], 1'b0);
    buf g30(n4[1], 1'b0);
    buf g31(n4[0], 1'b0);
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n599), .Q(n3[0]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n631), .Q(n3[1]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n630), .Q(n3[2]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n629), .Q(n3[3]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n628), .Q(n3[4]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n627), .Q(n3[5]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n633), .Q(n3[6]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n635), .Q(n3[7]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n622), .Q(n3[8]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n626), .Q(n3[9]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n625), .Q(n3[10]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n634), .Q(n3[11]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n623), .Q(n3[12]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n624), .Q(n3[13]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n632), .Q(n3[14]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n621), .Q(n3[15]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n620), .Q(n3[16]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n619), .Q(n3[17]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n618), .Q(n3[18]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n608), .Q(n3[19]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n616), .Q(n3[20]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n615), .Q(n3[21]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n614), .Q(n3[22]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n613), .Q(n3[23]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n612), .Q(n3[24]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n611), .Q(n3[25]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n610), .Q(n3[26]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n607), .Q(n3[27]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n609), .Q(n3[28]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n617), .Q(n3[29]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n606), .Q(n3[30]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n605), .Q(n3[31]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n638), .Q(n2));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n559), .Q(n774));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n693), .Q(n4[0]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n707), .Q(n4[1]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n706), .Q(n4[2]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n705), .Q(n4[3]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n704), .Q(n4[4]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n703), .Q(n4[5]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n702), .Q(n4[6]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n701), .Q(n4[7]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n700), .Q(n4[8]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n699), .Q(n4[9]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n698), .Q(n4[10]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n697), .Q(n4[11]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n694), .Q(n4[12]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n696), .Q(n4[13]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n695), .Q(n4[14]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n708), .Q(n4[15]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n677), .Q(n4[16]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n691), .Q(n4[17]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n690), .Q(n4[18]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n689), .Q(n4[19]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n688), .Q(n4[20]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n687), .Q(n4[21]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n686), .Q(n4[22]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n685), .Q(n4[23]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n684), .Q(n4[24]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n683), .Q(n4[25]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n682), .Q(n4[26]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n681), .Q(n4[27]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n680), .Q(n4[28]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n678), .Q(n4[29]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n679), .Q(n4[30]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n692), .Q(n4[31]));
    or g98(n708 ,n557 ,n676);
    or g99(n707 ,n596 ,n661);
    or g100(n706 ,n595 ,n675);
    or g101(n705 ,n593 ,n674);
    or g102(n704 ,n592 ,n673);
    or g103(n703 ,n591 ,n672);
    or g104(n702 ,n590 ,n671);
    or g105(n701 ,n589 ,n670);
    or g106(n700 ,n588 ,n668);
    or g107(n699 ,n586 ,n667);
    or g108(n698 ,n585 ,n666);
    or g109(n697 ,n583 ,n665);
    or g110(n696 ,n580 ,n663);
    or g111(n695 ,n579 ,n662);
    or g112(n694 ,n582 ,n664);
    or g113(n693 ,n564 ,n649);
    or g114(n692 ,n565 ,n660);
    or g115(n691 ,n573 ,n659);
    or g116(n690 ,n572 ,n658);
    or g117(n689 ,n570 ,n657);
    or g118(n688 ,n571 ,n656);
    or g119(n687 ,n597 ,n655);
    or g120(n686 ,n584 ,n654);
    or g121(n685 ,n568 ,n653);
    or g122(n684 ,n566 ,n651);
    or g123(n683 ,n594 ,n650);
    or g124(n682 ,n569 ,n652);
    or g125(n681 ,n598 ,n648);
    or g126(n680 ,n567 ,n647);
    or g127(n679 ,n587 ,n669);
    or g128(n678 ,n581 ,n646);
    or g129(n677 ,n574 ,n645);
    nor g130(n676 ,n489 ,n644);
    nor g131(n675 ,n515 ,n644);
    nor g132(n674 ,n475 ,n644);
    nor g133(n673 ,n495 ,n644);
    nor g134(n672 ,n492 ,n644);
    nor g135(n671 ,n487 ,n644);
    nor g136(n670 ,n525 ,n644);
    nor g137(n669 ,n535 ,n644);
    nor g138(n668 ,n484 ,n644);
    nor g139(n667 ,n473 ,n644);
    nor g140(n666 ,n500 ,n644);
    nor g141(n665 ,n503 ,n644);
    nor g142(n664 ,n513 ,n644);
    nor g143(n663 ,n504 ,n644);
    nor g144(n662 ,n501 ,n644);
    nor g145(n661 ,n528 ,n644);
    nor g146(n660 ,n507 ,n644);
    nor g147(n659 ,n482 ,n644);
    nor g148(n658 ,n472 ,n644);
    nor g149(n657 ,n511 ,n644);
    nor g150(n656 ,n505 ,n644);
    nor g151(n655 ,n467 ,n644);
    nor g152(n654 ,n486 ,n644);
    nor g153(n653 ,n485 ,n644);
    nor g154(n652 ,n496 ,n644);
    nor g155(n651 ,n517 ,n644);
    nor g156(n650 ,n532 ,n644);
    nor g157(n649 ,n514 ,n644);
    nor g158(n648 ,n510 ,n644);
    nor g159(n647 ,n529 ,n644);
    nor g160(n646 ,n477 ,n644);
    nor g161(n645 ,n478 ,n644);
    nor g162(n644 ,n578 ,n643);
    nor g163(n643 ,n636 ,n642);
    or g164(n642 ,n602 ,n641);
    or g165(n641 ,n554 ,n640);
    or g166(n640 ,n547 ,n639);
    or g167(n639 ,n561 ,n637);
    or g168(n638 ,n603 ,n604);
    or g169(n637 ,n556 ,n600);
    or g170(n636 ,n558 ,n601);
    nor g171(n635 ,n498 ,n577);
    nor g172(n634 ,n530 ,n577);
    nor g173(n633 ,n499 ,n577);
    nor g174(n632 ,n506 ,n577);
    nor g175(n631 ,n493 ,n577);
    nor g176(n630 ,n508 ,n577);
    nor g177(n629 ,n480 ,n577);
    nor g178(n628 ,n476 ,n577);
    nor g179(n627 ,n502 ,n577);
    nor g180(n626 ,n491 ,n577);
    nor g181(n625 ,n526 ,n577);
    nor g182(n624 ,n470 ,n577);
    nor g183(n623 ,n469 ,n577);
    nor g184(n622 ,n488 ,n577);
    nor g185(n621 ,n479 ,n577);
    nor g186(n620 ,n536 ,n577);
    nor g187(n619 ,n497 ,n577);
    nor g188(n618 ,n531 ,n577);
    nor g189(n617 ,n474 ,n577);
    nor g190(n616 ,n524 ,n577);
    nor g191(n615 ,n509 ,n577);
    nor g192(n614 ,n518 ,n577);
    nor g193(n613 ,n483 ,n577);
    nor g194(n612 ,n490 ,n577);
    nor g195(n611 ,n471 ,n577);
    nor g196(n610 ,n481 ,n577);
    nor g197(n609 ,n494 ,n577);
    nor g198(n608 ,n527 ,n577);
    nor g199(n607 ,n468 ,n577);
    nor g200(n606 ,n512 ,n577);
    nor g201(n605 ,n533 ,n577);
    nor g202(n604 ,n451 ,n577);
    nor g203(n603 ,n519 ,n576);
    or g204(n602 ,n562 ,n563);
    or g205(n601 ,n543 ,n575);
    or g206(n600 ,n4[25] ,n560);
    nor g207(n599 ,n3[0] ,n577);
    nor g208(n598 ,n463 ,n555);
    nor g209(n597 ,n465 ,n555);
    nor g210(n596 ,n442 ,n555);
    nor g211(n595 ,n520 ,n555);
    nor g212(n594 ,n466 ,n555);
    nor g213(n593 ,n439 ,n555);
    nor g214(n592 ,n450 ,n555);
    nor g215(n591 ,n456 ,n555);
    nor g216(n590 ,n460 ,n555);
    nor g217(n589 ,n457 ,n555);
    nor g218(n588 ,n452 ,n555);
    nor g219(n587 ,n455 ,n555);
    nor g220(n586 ,n523 ,n555);
    nor g221(n585 ,n454 ,n555);
    nor g222(n584 ,n449 ,n555);
    nor g223(n583 ,n440 ,n555);
    nor g224(n582 ,n521 ,n555);
    nor g225(n581 ,n441 ,n555);
    nor g226(n580 ,n458 ,n555);
    nor g227(n579 ,n444 ,n555);
    nor g228(n578 ,n464 ,n554);
    not g229(n577 ,n576);
    or g230(n575 ,n4[26] ,n552);
    nor g231(n574 ,n445 ,n555);
    nor g232(n573 ,n522 ,n555);
    nor g233(n572 ,n448 ,n555);
    nor g234(n571 ,n443 ,n555);
    nor g235(n570 ,n462 ,n555);
    nor g236(n569 ,n459 ,n555);
    nor g237(n568 ,n447 ,n555);
    nor g238(n567 ,n461 ,n555);
    nor g239(n566 ,n453 ,n555);
    nor g240(n565 ,n464 ,n555);
    nor g241(n564 ,n516 ,n555);
    or g242(n563 ,n548 ,n540);
    or g243(n562 ,n550 ,n553);
    or g244(n561 ,n551 ,n539);
    or g245(n560 ,n541 ,n542);
    nor g246(n559 ,n546 ,n544);
    or g247(n558 ,n537 ,n538);
    nor g248(n557 ,n446 ,n555);
    or g249(n556 ,n4[24] ,n549);
    nor g250(n576 ,n545 ,n544);
    not g251(n554 ,n555);
    or g252(n553 ,n4[21] ,n4[20]);
    nor g253(n552 ,n439 ,n520);
    or g254(n551 ,n4[9] ,n4[8]);
    or g255(n550 ,n4[29] ,n4[28]);
    nor g256(n549 ,n439 ,n442);
    or g257(n548 ,n4[23] ,n4[22]);
    or g258(n547 ,n4[7] ,n4[6]);
    nor g259(n555 ,n534 ,n1);
    not g260(n546 ,n545);
    or g261(n543 ,n4[30] ,n4[27]);
    or g262(n542 ,n4[13] ,n4[12]);
    or g263(n541 ,n4[19] ,n4[18]);
    or g264(n540 ,n4[11] ,n4[10]);
    or g265(n539 ,n4[5] ,n4[4]);
    or g266(n538 ,n4[15] ,n4[14]);
    or g267(n537 ,n4[17] ,n4[16]);
    nor g268(n545 ,n773 ,n739);
    or g269(n544 ,n1 ,n6);
    not g270(n536 ,n723);
    not g271(n535 ,n771);
    not g272(n534 ,n774);
    not g273(n533 ,n738);
    not g274(n532 ,n766);
    not g275(n531 ,n725);
    not g276(n530 ,n718);
    not g277(n529 ,n769);
    not g278(n528 ,n742);
    not g279(n527 ,n726);
    not g280(n526 ,n717);
    not g281(n525 ,n748);
    not g282(n524 ,n727);
    not g283(n523 ,n4[9]);
    not g284(n522 ,n4[17]);
    not g285(n521 ,n4[12]);
    not g286(n520 ,n4[2]);
    not g287(n519 ,n2);
    not g288(n518 ,n729);
    not g289(n517 ,n765);
    not g290(n516 ,n4[0]);
    not g291(n515 ,n743);
    not g292(n514 ,n741);
    not g293(n513 ,n753);
    not g294(n512 ,n737);
    not g295(n511 ,n760);
    not g296(n510 ,n768);
    not g297(n509 ,n728);
    not g298(n508 ,n709);
    not g299(n507 ,n772);
    not g300(n506 ,n721);
    not g301(n505 ,n761);
    not g302(n504 ,n754);
    not g303(n503 ,n752);
    not g304(n502 ,n712);
    not g305(n501 ,n755);
    not g306(n500 ,n751);
    not g307(n499 ,n713);
    not g308(n498 ,n714);
    not g309(n497 ,n724);
    not g310(n496 ,n767);
    not g311(n495 ,n745);
    not g312(n494 ,n735);
    not g313(n493 ,n740);
    not g314(n492 ,n746);
    not g315(n491 ,n716);
    not g316(n490 ,n731);
    not g317(n489 ,n756);
    not g318(n488 ,n715);
    not g319(n487 ,n747);
    not g320(n486 ,n763);
    not g321(n485 ,n764);
    not g322(n484 ,n749);
    not g323(n483 ,n730);
    not g324(n482 ,n758);
    not g325(n481 ,n733);
    not g326(n480 ,n710);
    not g327(n479 ,n722);
    not g328(n478 ,n757);
    not g329(n477 ,n770);
    not g330(n476 ,n711);
    not g331(n475 ,n744);
    not g332(n474 ,n736);
    not g333(n473 ,n750);
    not g334(n472 ,n759);
    not g335(n471 ,n732);
    not g336(n470 ,n720);
    not g337(n469 ,n719);
    not g338(n468 ,n734);
    not g339(n467 ,n762);
    not g340(n466 ,n4[25]);
    not g341(n465 ,n4[21]);
    not g342(n464 ,n4[31]);
    not g343(n463 ,n4[27]);
    not g344(n462 ,n4[19]);
    not g345(n461 ,n4[28]);
    not g346(n460 ,n4[6]);
    not g347(n459 ,n4[26]);
    not g348(n458 ,n4[13]);
    not g349(n457 ,n4[7]);
    not g350(n456 ,n4[5]);
    not g351(n455 ,n4[30]);
    not g352(n454 ,n4[10]);
    not g353(n453 ,n4[24]);
    not g354(n452 ,n4[8]);
    not g355(n451 ,n773);
    not g356(n450 ,n4[4]);
    not g357(n449 ,n4[22]);
    not g358(n448 ,n4[18]);
    not g359(n447 ,n4[23]);
    not g360(n446 ,n4[15]);
    not g361(n445 ,n4[16]);
    not g362(n444 ,n4[14]);
    not g363(n443 ,n4[20]);
    not g364(n442 ,n4[1]);
    not g365(n441 ,n4[29]);
    not g366(n440 ,n4[11]);
    not g367(n439 ,n4[3]);
    xor g368(n738 ,n3[31] ,n114);
    nor g369(n737 ,n113 ,n114);
    nor g370(n114 ,n37 ,n112);
    nor g371(n113 ,n3[30] ,n111);
    xor g372(n736 ,n3[29] ,n109);
    not g373(n112 ,n111);
    nor g374(n111 ,n24 ,n110);
    nor g375(n735 ,n108 ,n109);
    not g376(n110 ,n109);
    nor g377(n109 ,n35 ,n107);
    nor g378(n108 ,n3[28] ,n106);
    xor g379(n734 ,n3[27] ,n104);
    not g380(n107 ,n106);
    nor g381(n106 ,n10 ,n105);
    nor g382(n733 ,n103 ,n104);
    xor g383(n732 ,n3[25] ,n102);
    not g384(n105 ,n104);
    nor g385(n104 ,n22 ,n101);
    nor g386(n103 ,n3[26] ,n100);
    nor g387(n731 ,n99 ,n102);
    nor g388(n102 ,n20 ,n98);
    not g389(n101 ,n100);
    nor g390(n100 ,n43 ,n98);
    nor g391(n99 ,n3[24] ,n97);
    xor g392(n730 ,n3[23] ,n95);
    not g393(n98 ,n97);
    nor g394(n97 ,n9 ,n96);
    nor g395(n729 ,n94 ,n95);
    xor g396(n728 ,n3[21] ,n93);
    xor g397(n726 ,n3[19] ,n92);
    not g398(n96 ,n95);
    nor g399(n95 ,n36 ,n91);
    nor g400(n94 ,n3[22] ,n90);
    nor g401(n727 ,n89 ,n93);
    nor g402(n725 ,n88 ,n92);
    xor g403(n724 ,n3[17] ,n87);
    nor g404(n93 ,n31 ,n84);
    nor g405(n92 ,n19 ,n86);
    not g406(n91 ,n90);
    nor g407(n90 ,n46 ,n84);
    nor g408(n89 ,n3[20] ,n83);
    nor g409(n88 ,n3[18] ,n85);
    nor g410(n723 ,n82 ,n87);
    nor g411(n87 ,n15 ,n81);
    not g412(n86 ,n85);
    nor g413(n85 ,n44 ,n81);
    not g414(n84 ,n83);
    nor g415(n83 ,n54 ,n81);
    nor g416(n82 ,n3[16] ,n80);
    xor g417(n722 ,n3[15] ,n78);
    not g418(n81 ,n80);
    nor g419(n80 ,n30 ,n79);
    nor g420(n721 ,n77 ,n78);
    xor g421(n720 ,n3[13] ,n76);
    xor g422(n718 ,n3[11] ,n75);
    or g423(n79 ,n13 ,n74);
    nor g424(n78 ,n30 ,n74);
    nor g425(n77 ,n3[14] ,n73);
    nor g426(n719 ,n71 ,n76);
    nor g427(n717 ,n72 ,n75);
    xor g428(n716 ,n3[9] ,n70);
    nor g429(n76 ,n18 ,n69);
    nor g430(n75 ,n16 ,n67);
    not g431(n74 ,n73);
    nor g432(n73 ,n45 ,n69);
    nor g433(n72 ,n3[10] ,n66);
    nor g434(n71 ,n3[12] ,n68);
    nor g435(n715 ,n65 ,n70);
    nor g436(n70 ,n25 ,n64);
    not g437(n69 ,n68);
    nor g438(n68 ,n55 ,n64);
    not g439(n67 ,n66);
    nor g440(n66 ,n42 ,n64);
    nor g441(n65 ,n3[8] ,n63);
    xor g442(n714 ,n3[7] ,n62);
    not g443(n64 ,n63);
    nor g444(n63 ,n27 ,n61);
    nor g445(n713 ,n60 ,n62);
    xor g446(n712 ,n3[5] ,n59);
    nor g447(n62 ,n27 ,n58);
    or g448(n61 ,n23 ,n58);
    nor g449(n60 ,n3[6] ,n57);
    nor g450(n711 ,n56 ,n59);
    nor g451(n59 ,n12 ,n53);
    not g452(n58 ,n57);
    nor g453(n57 ,n41 ,n53);
    nor g454(n56 ,n3[4] ,n52);
    xor g455(n710 ,n3[3] ,n50);
    or g456(n55 ,n16 ,n48);
    or g457(n54 ,n19 ,n51);
    not g458(n53 ,n52);
    nor g459(n52 ,n7 ,n49);
    nor g460(n709 ,n47 ,n50);
    or g461(n51 ,n14 ,n44);
    nor g462(n50 ,n32 ,n40);
    or g463(n49 ,n32 ,n40);
    or g464(n48 ,n11 ,n42);
    nor g465(n47 ,n3[2] ,n39);
    nor g466(n740 ,n39 ,n38);
    or g467(n46 ,n26 ,n31);
    or g468(n45 ,n8 ,n18);
    or g469(n44 ,n33 ,n15);
    or g470(n43 ,n17 ,n20);
    or g471(n42 ,n28 ,n25);
    or g472(n41 ,n29 ,n12);
    not g473(n40 ,n39);
    nor g474(n39 ,n21 ,n34);
    nor g475(n38 ,n3[1] ,n3[0]);
    not g476(n37 ,n3[30]);
    not g477(n36 ,n3[22]);
    not g478(n35 ,n3[28]);
    not g479(n34 ,n3[0]);
    not g480(n33 ,n3[17]);
    not g481(n32 ,n3[2]);
    not g482(n31 ,n3[20]);
    not g483(n30 ,n3[14]);
    not g484(n29 ,n3[5]);
    not g485(n28 ,n3[9]);
    not g486(n27 ,n3[6]);
    not g487(n26 ,n3[21]);
    not g488(n25 ,n3[8]);
    not g489(n24 ,n3[29]);
    not g490(n23 ,n3[7]);
    not g491(n22 ,n3[26]);
    not g492(n21 ,n3[1]);
    not g493(n20 ,n3[24]);
    not g494(n19 ,n3[18]);
    not g495(n18 ,n3[12]);
    not g496(n17 ,n3[25]);
    not g497(n16 ,n3[10]);
    not g498(n15 ,n3[16]);
    not g499(n14 ,n3[19]);
    not g500(n13 ,n3[15]);
    not g501(n12 ,n3[4]);
    not g502(n11 ,n3[11]);
    not g503(n10 ,n3[27]);
    not g504(n9 ,n3[23]);
    not g505(n8 ,n3[13]);
    not g506(n7 ,n3[3]);
    xor g507(n772 ,n221 ,n4[31]);
    nor g508(n771 ,n220 ,n221);
    nor g509(n221 ,n144 ,n219);
    nor g510(n220 ,n4[30] ,n218);
    xor g511(n770 ,n216 ,n4[29]);
    not g512(n219 ,n218);
    nor g513(n218 ,n132 ,n217);
    nor g514(n769 ,n215 ,n216);
    not g515(n217 ,n216);
    nor g516(n216 ,n142 ,n214);
    nor g517(n215 ,n4[28] ,n213);
    xor g518(n768 ,n211 ,n4[27]);
    not g519(n214 ,n213);
    nor g520(n213 ,n118 ,n212);
    nor g521(n767 ,n210 ,n211);
    xor g522(n766 ,n209 ,n4[25]);
    not g523(n212 ,n211);
    nor g524(n211 ,n130 ,n208);
    nor g525(n210 ,n4[26] ,n207);
    nor g526(n765 ,n206 ,n209);
    nor g527(n209 ,n128 ,n205);
    not g528(n208 ,n207);
    nor g529(n207 ,n150 ,n205);
    nor g530(n206 ,n4[24] ,n204);
    xor g531(n764 ,n202 ,n4[23]);
    not g532(n205 ,n204);
    nor g533(n204 ,n117 ,n203);
    nor g534(n763 ,n201 ,n202);
    xor g535(n762 ,n200 ,n4[21]);
    xor g536(n760 ,n199 ,n4[19]);
    not g537(n203 ,n202);
    nor g538(n202 ,n143 ,n198);
    nor g539(n201 ,n4[22] ,n197);
    nor g540(n761 ,n196 ,n200);
    nor g541(n759 ,n195 ,n199);
    xor g542(n758 ,n194 ,n4[17]);
    nor g543(n200 ,n138 ,n191);
    nor g544(n199 ,n127 ,n193);
    not g545(n198 ,n197);
    nor g546(n197 ,n153 ,n191);
    nor g547(n196 ,n4[20] ,n190);
    nor g548(n195 ,n4[18] ,n192);
    nor g549(n757 ,n189 ,n194);
    nor g550(n194 ,n123 ,n188);
    not g551(n193 ,n192);
    nor g552(n192 ,n151 ,n188);
    not g553(n191 ,n190);
    nor g554(n190 ,n161 ,n188);
    nor g555(n189 ,n4[16] ,n187);
    xor g556(n756 ,n185 ,n4[15]);
    not g557(n188 ,n187);
    nor g558(n187 ,n137 ,n186);
    nor g559(n755 ,n184 ,n185);
    xor g560(n754 ,n183 ,n4[13]);
    xor g561(n752 ,n182 ,n4[11]);
    or g562(n186 ,n121 ,n181);
    nor g563(n185 ,n137 ,n181);
    nor g564(n184 ,n4[14] ,n180);
    nor g565(n753 ,n178 ,n183);
    nor g566(n751 ,n179 ,n182);
    xor g567(n750 ,n177 ,n4[9]);
    nor g568(n183 ,n126 ,n176);
    nor g569(n182 ,n124 ,n174);
    not g570(n181 ,n180);
    nor g571(n180 ,n152 ,n176);
    nor g572(n179 ,n4[10] ,n173);
    nor g573(n178 ,n4[12] ,n175);
    nor g574(n749 ,n172 ,n177);
    nor g575(n177 ,n133 ,n171);
    not g576(n176 ,n175);
    nor g577(n175 ,n162 ,n171);
    not g578(n174 ,n173);
    nor g579(n173 ,n149 ,n171);
    nor g580(n172 ,n4[8] ,n170);
    xor g581(n748 ,n169 ,n4[7]);
    not g582(n171 ,n170);
    nor g583(n170 ,n135 ,n168);
    nor g584(n747 ,n167 ,n169);
    xor g585(n746 ,n166 ,n4[5]);
    nor g586(n169 ,n135 ,n165);
    or g587(n168 ,n131 ,n165);
    nor g588(n167 ,n4[6] ,n164);
    nor g589(n745 ,n163 ,n166);
    nor g590(n166 ,n120 ,n160);
    not g591(n165 ,n164);
    nor g592(n164 ,n148 ,n160);
    nor g593(n163 ,n4[4] ,n159);
    xor g594(n744 ,n157 ,n4[3]);
    or g595(n162 ,n124 ,n155);
    or g596(n161 ,n127 ,n158);
    not g597(n160 ,n159);
    nor g598(n159 ,n115 ,n156);
    nor g599(n743 ,n154 ,n157);
    or g600(n158 ,n122 ,n151);
    nor g601(n157 ,n139 ,n147);
    or g602(n156 ,n139 ,n147);
    or g603(n155 ,n119 ,n149);
    nor g604(n154 ,n4[2] ,n146);
    nor g605(n742 ,n146 ,n145);
    or g606(n153 ,n141 ,n138);
    or g607(n152 ,n116 ,n126);
    or g608(n151 ,n140 ,n123);
    or g609(n150 ,n125 ,n128);
    or g610(n149 ,n134 ,n133);
    or g611(n148 ,n136 ,n120);
    not g612(n147 ,n146);
    nor g613(n146 ,n129 ,n741);
    nor g614(n145 ,n4[1] ,n4[0]);
    not g615(n144 ,n4[30]);
    not g616(n143 ,n4[22]);
    not g617(n142 ,n4[28]);
    not g618(n141 ,n4[21]);
    not g619(n140 ,n4[17]);
    not g620(n139 ,n4[2]);
    not g621(n138 ,n4[20]);
    not g622(n137 ,n4[14]);
    not g623(n136 ,n4[5]);
    not g624(n741 ,n4[0]);
    not g625(n135 ,n4[6]);
    not g626(n134 ,n4[9]);
    not g627(n133 ,n4[8]);
    not g628(n132 ,n4[29]);
    not g629(n131 ,n4[7]);
    not g630(n130 ,n4[26]);
    not g631(n129 ,n4[1]);
    not g632(n128 ,n4[24]);
    not g633(n127 ,n4[18]);
    not g634(n126 ,n4[12]);
    not g635(n125 ,n4[25]);
    not g636(n124 ,n4[10]);
    not g637(n123 ,n4[16]);
    not g638(n122 ,n4[19]);
    not g639(n121 ,n4[15]);
    not g640(n120 ,n4[4]);
    not g641(n119 ,n4[11]);
    not g642(n118 ,n4[27]);
    not g643(n117 ,n4[23]);
    not g644(n116 ,n4[13]);
    not g645(n115 ,n4[3]);
    or g646(n739 ,n3[31] ,n251);
    nor g647(n251 ,n247 ,n250);
    or g648(n250 ,n249 ,n248);
    or g649(n249 ,n236 ,n244);
    or g650(n248 ,n246 ,n245);
    or g651(n247 ,n241 ,n239);
    or g652(n246 ,n242 ,n240);
    or g653(n245 ,n238 ,n237);
    or g654(n244 ,n3[4] ,n243);
    nor g655(n243 ,n222 ,n229);
    or g656(n242 ,n235 ,n233);
    or g657(n241 ,n228 ,n234);
    or g658(n240 ,n231 ,n223);
    or g659(n239 ,n226 ,n230);
    or g660(n238 ,n227 ,n232);
    or g661(n237 ,n225 ,n224);
    or g662(n236 ,n3[6] ,n3[5]);
    or g663(n235 ,n3[30] ,n3[29]);
    or g664(n234 ,n3[12] ,n3[11]);
    or g665(n233 ,n3[28] ,n3[27]);
    or g666(n232 ,n3[20] ,n3[19]);
    or g667(n231 ,n3[26] ,n3[25]);
    or g668(n230 ,n3[8] ,n3[7]);
    nor g669(n229 ,n3[2] ,n3[1]);
    or g670(n228 ,n3[14] ,n3[13]);
    or g671(n227 ,n3[22] ,n3[21]);
    or g672(n226 ,n3[10] ,n3[9]);
    or g673(n225 ,n3[18] ,n3[17]);
    or g674(n224 ,n3[16] ,n3[15]);
    or g675(n223 ,n3[24] ,n3[23]);
    not g676(n222 ,n3[3]);
    or g677(n773 ,n343 ,n438);
    nor g678(n438 ,n383 ,n437);
    nor g679(n437 ,n386 ,n436);
    nor g680(n436 ,n408 ,n435);
    nor g681(n435 ,n388 ,n434);
    nor g682(n434 ,n379 ,n433);
    nor g683(n433 ,n403 ,n432);
    nor g684(n432 ,n395 ,n431);
    nor g685(n431 ,n390 ,n430);
    nor g686(n430 ,n385 ,n429);
    nor g687(n429 ,n381 ,n428);
    nor g688(n428 ,n401 ,n427);
    nor g689(n427 ,n405 ,n426);
    nor g690(n426 ,n400 ,n425);
    nor g691(n425 ,n397 ,n424);
    nor g692(n424 ,n378 ,n423);
    nor g693(n423 ,n389 ,n422);
    nor g694(n422 ,n387 ,n421);
    nor g695(n421 ,n384 ,n420);
    nor g696(n420 ,n382 ,n419);
    nor g697(n419 ,n380 ,n418);
    nor g698(n418 ,n393 ,n417);
    nor g699(n417 ,n407 ,n416);
    nor g700(n416 ,n406 ,n415);
    nor g701(n415 ,n404 ,n414);
    nor g702(n414 ,n402 ,n413);
    nor g703(n413 ,n399 ,n412);
    nor g704(n412 ,n398 ,n411);
    nor g705(n411 ,n396 ,n410);
    nor g706(n410 ,n394 ,n409);
    nor g707(n409 ,n392 ,n391);
    or g708(n408 ,n356 ,n348);
    or g709(n407 ,n374 ,n372);
    or g710(n406 ,n369 ,n368);
    or g711(n405 ,n363 ,n347);
    or g712(n404 ,n364 ,n362);
    or g713(n403 ,n360 ,n354);
    or g714(n402 ,n359 ,n357);
    or g715(n401 ,n373 ,n370);
    or g716(n400 ,n353 ,n352);
    or g717(n399 ,n365 ,n361);
    or g718(n398 ,n350 ,n349);
    or g719(n397 ,n330 ,n324);
    or g720(n396 ,n375 ,n331);
    or g721(n395 ,n345 ,n341);
    or g722(n394 ,n371 ,n344);
    or g723(n393 ,n315 ,n377);
    nor g724(n392 ,n346 ,n339);
    or g725(n391 ,n337 ,n342);
    or g726(n390 ,n335 ,n332);
    or g727(n389 ,n336 ,n334);
    or g728(n388 ,n333 ,n355);
    or g729(n387 ,n351 ,n329);
    or g730(n386 ,n328 ,n367);
    or g731(n385 ,n326 ,n325);
    or g732(n384 ,n327 ,n358);
    or g733(n383 ,n321 ,n366);
    or g734(n382 ,n323 ,n322);
    or g735(n381 ,n319 ,n316);
    or g736(n380 ,n320 ,n318);
    or g737(n379 ,n317 ,n376);
    or g738(n378 ,n340 ,n338);
    nor g739(n377 ,n253 ,n4[10]);
    nor g740(n376 ,n272 ,n4[26]);
    nor g741(n375 ,n313 ,n3[4]);
    nor g742(n374 ,n274 ,n3[10]);
    nor g743(n373 ,n267 ,n4[21]);
    nor g744(n372 ,n309 ,n3[9]);
    nor g745(n371 ,n258 ,n4[3]);
    nor g746(n370 ,n301 ,n4[20]);
    nor g747(n369 ,n286 ,n4[9]);
    nor g748(n368 ,n294 ,n4[8]);
    nor g749(n367 ,n280 ,n3[29]);
    nor g750(n366 ,n276 ,n4[30]);
    nor g751(n365 ,n308 ,n3[6]);
    nor g752(n364 ,n292 ,n3[8]);
    nor g753(n363 ,n269 ,n3[20]);
    nor g754(n362 ,n252 ,n3[7]);
    nor g755(n361 ,n300 ,n3[5]);
    nor g756(n360 ,n299 ,n3[26]);
    nor g757(n359 ,n289 ,n4[7]);
    nor g758(n358 ,n288 ,n3[13]);
    nor g759(n357 ,n296 ,n4[6]);
    nor g760(n356 ,n306 ,n4[29]);
    nor g761(n355 ,n259 ,n3[27]);
    nor g762(n354 ,n278 ,n3[25]);
    nor g763(n353 ,n298 ,n4[19]);
    nor g764(n352 ,n262 ,n4[18]);
    nor g765(n351 ,n271 ,n4[15]);
    nor g766(n350 ,n282 ,n4[5]);
    nor g767(n349 ,n302 ,n4[4]);
    nor g768(n348 ,n279 ,n4[28]);
    nor g769(n347 ,n275 ,n3[19]);
    nor g770(n346 ,n307 ,n4[1]);
    nor g771(n345 ,n257 ,n4[25]);
    nor g772(n344 ,n255 ,n4[2]);
    nor g773(n343 ,n295 ,n4[31]);
    nor g774(n342 ,n283 ,n3[1]);
    nor g775(n341 ,n293 ,n4[24]);
    nor g776(n340 ,n263 ,n4[17]);
    nor g777(n339 ,n314 ,n4[0]);
    nor g778(n338 ,n303 ,n4[16]);
    nor g779(n337 ,n273 ,n3[2]);
    nor g780(n336 ,n261 ,n3[16]);
    nor g781(n335 ,n304 ,n3[24]);
    nor g782(n334 ,n260 ,n3[15]);
    nor g783(n333 ,n281 ,n3[28]);
    nor g784(n332 ,n291 ,n3[23]);
    nor g785(n331 ,n305 ,n3[3]);
    nor g786(n330 ,n277 ,n3[18]);
    nor g787(n329 ,n290 ,n4[14]);
    nor g788(n328 ,n311 ,n3[30]);
    nor g789(n327 ,n254 ,n3[14]);
    nor g790(n326 ,n270 ,n4[23]);
    nor g791(n325 ,n268 ,n4[22]);
    nor g792(n324 ,n297 ,n3[17]);
    nor g793(n323 ,n256 ,n4[13]);
    nor g794(n322 ,n310 ,n4[12]);
    nor g795(n321 ,n266 ,n3[31]);
    nor g796(n320 ,n285 ,n3[12]);
    nor g797(n319 ,n264 ,n3[22]);
    nor g798(n318 ,n284 ,n3[11]);
    nor g799(n317 ,n287 ,n4[27]);
    nor g800(n316 ,n265 ,n3[21]);
    nor g801(n315 ,n312 ,n4[11]);
    not g802(n314 ,n3[0]);
    not g803(n313 ,n4[4]);
    not g804(n312 ,n3[11]);
    not g805(n311 ,n4[30]);
    not g806(n310 ,n3[12]);
    not g807(n309 ,n4[9]);
    not g808(n308 ,n4[6]);
    not g809(n307 ,n3[1]);
    not g810(n306 ,n3[29]);
    not g811(n305 ,n4[3]);
    not g812(n304 ,n4[24]);
    not g813(n303 ,n3[16]);
    not g814(n302 ,n3[4]);
    not g815(n301 ,n3[20]);
    not g816(n300 ,n4[5]);
    not g817(n299 ,n4[26]);
    not g818(n298 ,n3[19]);
    not g819(n297 ,n4[17]);
    not g820(n296 ,n3[6]);
    not g821(n295 ,n3[31]);
    not g822(n294 ,n3[8]);
    not g823(n293 ,n3[24]);
    not g824(n292 ,n4[8]);
    not g825(n291 ,n4[23]);
    not g826(n290 ,n3[14]);
    not g827(n289 ,n3[7]);
    not g828(n288 ,n4[13]);
    not g829(n287 ,n3[27]);
    not g830(n286 ,n3[9]);
    not g831(n285 ,n4[12]);
    not g832(n284 ,n4[11]);
    not g833(n283 ,n4[1]);
    not g834(n282 ,n3[5]);
    not g835(n281 ,n4[28]);
    not g836(n280 ,n4[29]);
    not g837(n279 ,n3[28]);
    not g838(n278 ,n4[25]);
    not g839(n277 ,n4[18]);
    not g840(n276 ,n3[30]);
    not g841(n275 ,n4[19]);
    not g842(n274 ,n4[10]);
    not g843(n273 ,n4[2]);
    not g844(n272 ,n3[26]);
    not g845(n271 ,n3[15]);
    not g846(n270 ,n3[23]);
    not g847(n269 ,n4[20]);
    not g848(n268 ,n3[22]);
    not g849(n267 ,n3[21]);
    not g850(n266 ,n4[31]);
    not g851(n265 ,n4[21]);
    not g852(n264 ,n4[22]);
    not g853(n263 ,n3[17]);
    not g854(n262 ,n3[18]);
    not g855(n261 ,n4[16]);
    not g856(n260 ,n4[15]);
    not g857(n259 ,n4[27]);
    not g858(n258 ,n3[3]);
    not g859(n257 ,n3[25]);
    not g860(n256 ,n3[13]);
    not g861(n255 ,n3[2]);
    not g862(n254 ,n4[14]);
    not g863(n253 ,n3[10]);
    not g864(n252 ,n4[7]);
    dff g865(.RN(n775), .SN(1'b1), .CK(n0), .D(n798), .Q(n6));
    nor g866(n798 ,n797 ,n796);
    or g867(n797 ,n792 ,n795);
    or g868(n796 ,n793 ,n794);
    or g869(n795 ,n790 ,n789);
    or g870(n794 ,n791 ,n786);
    or g871(n793 ,n785 ,n784);
    or g872(n792 ,n788 ,n787);
    dff g873(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[4]), .Q(n5[4]));
    dff g874(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[1]), .Q(n5[1]));
    dff g875(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[2]), .Q(n5[2]));
    dff g876(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[3]), .Q(n5[3]));
    dff g877(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[0]), .Q(n5[0]));
    dff g878(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[5]), .Q(n5[5]));
    dff g879(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[7]), .Q(n5[7]));
    dff g880(.RN(n775), .SN(1'b1), .CK(n0), .D(n3[6]), .Q(n5[6]));
    or g881(n791 ,n3[5] ,n3[3]);
    or g882(n790 ,n779 ,n778);
    or g883(n789 ,n776 ,n777);
    or g884(n788 ,n780 ,n783);
    or g885(n787 ,n782 ,n781);
    or g886(n786 ,n3[7] ,n3[1]);
    or g887(n785 ,n5[0] ,n5[2]);
    or g888(n784 ,n5[4] ,n5[6]);
    not g889(n783 ,n5[3]);
    not g890(n782 ,n5[5]);
    not g891(n781 ,n5[7]);
    not g892(n780 ,n5[1]);
    not g893(n779 ,n3[6]);
    not g894(n778 ,n3[4]);
    not g895(n777 ,n3[0]);
    not g896(n776 ,n3[2]);
    not g897(n775 ,n1);
endmodule
