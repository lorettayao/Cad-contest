
module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   CRC_OUT_1_14, CRC_OUT_1_31, CRC_OUT_2_19, CRC_OUT_2_2, CRC_OUT_3_24,
         CRC_OUT_3_7, CRC_OUT_4_12, CRC_OUT_4_29, CRC_OUT_5_0, CRC_OUT_5_17,
         CRC_OUT_6_22, CRC_OUT_6_5, CRC_OUT_7_10, CRC_OUT_7_27, CRC_OUT_8_25,
         CRC_OUT_8_7, CRC_OUT_9_1, CRC_OUT_9_19, WX485, WX484, WX487, WX486,
         WX489, WX488, WX491, WX490, WX493, WX492, WX495, WX494, WX497, WX496,
         WX499, WX498, WX501, WX500, WX503, WX502, WX505, WX504, WX507, WX506,
         WX509, WX508, WX511, WX510, WX513, WX512, WX515, WX514, WX517, WX516,
         WX518, WX521, WX520, WX523, WX522, WX525, WX524, WX527, WX526, WX529,
         WX528, WX531, WX530, WX533, WX532, WX535, WX534, WX537, WX536, WX539,
         WX538, WX541, WX540, WX543, WX542, WX545, WX544, WX547, WX546, WX645,
         WX644, WX647, WX646, WX649, WX648, WX650, WX653, WX652, WX655, WX654,
         WX657, WX656, WX659, WX658, WX661, WX660, WX663, WX662, WX665, WX664,
         WX667, WX666, WX669, WX668, WX671, WX670, WX673, WX672, WX675, WX674,
         WX677, WX676, WX679, WX678, WX681, WX680, WX683, WX682, WX685, WX684,
         WX686, WX689, WX688, WX691, WX690, WX693, WX692, WX695, WX694, WX697,
         WX696, WX699, WX698, WX701, WX700, WX703, WX702, WX705, WX704, WX707,
         WX706, WX709, WX708, WX711, WX710, WX713, WX712, WX715, WX714, WX717,
         WX716, WX719, WX718, WX721, WX720, WX722, WX725, WX724, WX727, WX726,
         WX729, WX728, WX731, WX730, WX733, WX732, WX735, WX734, WX737, WX736,
         WX739, WX738, WX741, WX740, WX743, WX742, WX745, WX744, WX747, WX746,
         WX749, WX748, WX751, WX750, WX753, WX752, WX755, WX754, WX757, WX756,
         WX758, WX761, WX760, WX763, WX762, WX765, WX764, WX767, WX766, WX769,
         WX768, WX771, WX770, WX773, WX772, WX775, WX774, WX777, WX776, WX779,
         WX778, WX781, WX780, WX783, WX782, WX785, WX784, WX787, WX786, WX789,
         WX788, WX791, WX790, WX793, WX792, WX794, WX797, WX796, WX799, WX798,
         WX801, WX800, WX803, WX802, WX805, WX804, WX807, WX806, WX809, WX808,
         WX811, WX810, WX813, WX812, WX815, WX814, WX817, WX816, WX819, WX818,
         WX821, WX820, WX823, WX822, WX825, WX824, WX827, WX826, WX829, WX828,
         WX830, WX833, WX832, WX835, WX834, WX837, WX836, WX839, WX838, WX841,
         WX840, WX843, WX842, WX845, WX844, WX847, WX846, WX849, WX848, WX851,
         WX850, WX853, WX852, WX855, WX854, WX857, WX856, WX859, WX858, WX861,
         WX860, WX863, WX862, WX865, WX864, WX866, WX869, WX868, WX871, WX870,
         WX873, WX872, WX875, WX874, WX877, WX876, WX879, WX878, WX881, WX880,
         WX883, WX882, WX885, WX884, WX887, WX886, WX889, WX888, WX891, WX890,
         WX893, WX892, WX895, WX894, WX897, WX896, WX899, WX898, WX1264,
         WX1266, WX1268, WX1270, WX1272, WX1274, WX1276, WX1278, WX1280,
         WX1282, WX1284, WX1286, WX1288, WX1290, WX1292, WX1294, WX1296,
         WX1298, WX1300, WX1302, WX1304, WX1306, WX1308, WX1310, WX1312,
         WX1314, WX1316, WX1318, WX1320, WX1322, WX1324, WX1326, WX1778,
         WX1777, WX1779, WX1781, WX1783, WX1785, WX1787, WX1789, WX1791,
         WX1793, WX1795, WX1797, WX1799, WX1801, WX1803, WX1805, WX1807,
         WX1809, WX1811, WX1813, WX1815, WX1817, WX1819, WX1821, WX1823,
         WX1825, WX1827, WX1829, WX1831, WX1833, WX1835, WX1837, WX1839,
         WX1937, WX1939, WX1941, WX1943, WX1945, WX1947, WX1949, WX1951,
         WX1953, WX1955, WX1957, WX1959, WX1961, WX1963, WX1965, WX1967,
         WX1970, WX1969, WX1972, WX1971, WX1974, WX1973, WX1976, WX1975,
         WX1978, WX1977, WX1980, WX1979, WX1982, WX1981, WX1984, WX1983,
         WX1986, WX1985, WX1988, WX1987, WX1990, WX1989, WX1991, WX1994,
         WX1993, WX1996, WX1995, WX1998, WX1997, WX2000, WX1999, WX2002,
         WX2001, WX2004, WX2003, WX2006, WX2005, WX2008, WX2007, WX2010,
         WX2009, WX2012, WX2011, WX2014, WX2013, WX2016, WX2015, WX2018,
         WX2017, WX2020, WX2019, WX2022, WX2021, WX2024, WX2023, WX2026,
         WX2025, WX2027, WX2030, WX2029, WX2032, WX2031, WX2034, WX2033,
         WX2036, WX2035, WX2038, WX2037, WX2040, WX2039, WX2042, WX2041,
         WX2044, WX2043, WX2046, WX2045, WX2048, WX2047, WX2050, WX2049,
         WX2052, WX2051, WX2054, WX2053, WX2056, WX2055, WX2058, WX2057,
         WX2060, WX2059, WX2062, WX2061, WX2063, WX2066, WX2065, WX2068,
         WX2067, WX2070, WX2069, WX2072, WX2071, WX2074, WX2073, WX2076,
         WX2075, WX2078, WX2077, WX2080, WX2079, WX2082, WX2081, WX2084,
         WX2083, WX2086, WX2085, WX2088, WX2087, WX2090, WX2089, WX2092,
         WX2091, WX2094, WX2093, WX2096, WX2095, WX2098, WX2097, WX2099,
         WX2102, WX2101, WX2104, WX2103, WX2106, WX2105, WX2108, WX2107,
         WX2110, WX2109, WX2112, WX2111, WX2114, WX2113, WX2116, WX2115,
         WX2118, WX2117, WX2120, WX2119, WX2122, WX2121, WX2124, WX2123,
         WX2126, WX2125, WX2128, WX2127, WX2130, WX2129, WX2132, WX2131,
         WX2134, WX2133, WX2135, WX2138, WX2137, WX2140, WX2139, WX2142,
         WX2141, WX2144, WX2143, WX2146, WX2145, WX2148, WX2147, WX2150,
         WX2149, WX2152, WX2151, WX2154, WX2153, WX2156, WX2155, WX2158,
         WX2157, WX2160, WX2159, WX2162, WX2161, WX2164, WX2163, WX2166,
         WX2165, WX2168, WX2167, WX2170, WX2169, WX2171, WX2174, WX2173,
         WX2176, WX2175, WX2178, WX2177, WX2180, WX2179, WX2182, WX2181,
         WX2184, WX2183, WX2186, WX2185, WX2188, WX2187, WX2190, WX2189,
         WX2192, WX2191, WX2557, WX2559, WX2561, WX2563, WX2565, WX2567,
         WX2569, WX2571, WX2573, WX2575, WX2577, WX2579, WX2581, WX2583,
         WX2585, WX2587, WX2589, WX2591, WX2593, WX2595, WX2597, WX2599,
         WX2601, WX2603, WX2605, WX2607, WX2609, WX2611, WX2613, WX2615,
         WX2617, WX2619, WX3071, WX3070, WX3072, WX3074, WX3076, WX3078,
         WX3080, WX3082, WX3084, WX3086, WX3088, WX3090, WX3092, WX3094,
         WX3096, WX3098, WX3100, WX3102, WX3104, WX3106, WX3108, WX3110,
         WX3112, WX3114, WX3116, WX3118, WX3120, WX3122, WX3124, WX3126,
         WX3128, WX3130, WX3132, WX3230, WX3232, WX3234, WX3236, WX3238,
         WX3240, WX3242, WX3244, WX3246, WX3248, WX3250, WX3252, WX3254,
         WX3256, WX3258, WX3260, WX3263, WX3262, WX3265, WX3264, WX3267,
         WX3266, WX3269, WX3268, WX3271, WX3270, WX3273, WX3272, WX3275,
         WX3274, WX3277, WX3276, WX3279, WX3278, WX3281, WX3280, WX3283,
         WX3282, WX3285, WX3284, WX3287, WX3286, WX3289, WX3288, WX3291,
         WX3290, WX3293, WX3292, WX3295, WX3294, WX3296, WX3299, WX3298,
         WX3301, WX3300, WX3303, WX3302, WX3305, WX3304, WX3307, WX3306,
         WX3309, WX3308, WX3311, WX3310, WX3313, WX3312, WX3315, WX3314,
         WX3317, WX3316, WX3319, WX3318, WX3321, WX3320, WX3323, WX3322,
         WX3325, WX3324, WX3327, WX3326, WX3329, WX3328, WX3331, WX3330,
         WX3332, WX3335, WX3334, WX3337, WX3336, WX3339, WX3338, WX3341,
         WX3340, WX3343, WX3342, WX3345, WX3344, WX3347, WX3346, WX3349,
         WX3348, WX3351, WX3350, WX3353, WX3352, WX3355, WX3354, WX3357,
         WX3356, WX3359, WX3358, WX3361, WX3360, WX3363, WX3362, WX3365,
         WX3364, WX3367, WX3366, WX3368, WX3371, WX3370, WX3373, WX3372,
         WX3375, WX3374, WX3377, WX3376, WX3379, WX3378, WX3381, WX3380,
         WX3383, WX3382, WX3385, WX3384, WX3387, WX3386, WX3389, WX3388,
         WX3391, WX3390, WX3393, WX3392, WX3395, WX3394, WX3397, WX3396,
         WX3399, WX3398, WX3401, WX3400, WX3403, WX3402, WX3404, WX3407,
         WX3406, WX3409, WX3408, WX3411, WX3410, WX3413, WX3412, WX3415,
         WX3414, WX3417, WX3416, WX3419, WX3418, WX3421, WX3420, WX3423,
         WX3422, WX3425, WX3424, WX3427, WX3426, WX3429, WX3428, WX3431,
         WX3430, WX3433, WX3432, WX3435, WX3434, WX3437, WX3436, WX3438,
         WX3441, WX3440, WX3443, WX3442, WX3445, WX3444, WX3447, WX3446,
         WX3449, WX3448, WX3451, WX3450, WX3453, WX3452, WX3455, WX3454,
         WX3457, WX3456, WX3459, WX3458, WX3461, WX3460, WX3463, WX3462,
         WX3465, WX3464, WX3467, WX3466, WX3469, WX3468, WX3471, WX3470,
         WX3472, WX3475, WX3474, WX3477, WX3476, WX3479, WX3478, WX3481,
         WX3480, WX3483, WX3482, WX3485, WX3484, WX3850, WX3852, WX3854,
         WX3856, WX3858, WX3860, WX3862, WX3864, WX3866, WX3868, WX3870,
         WX3872, WX3874, WX3876, WX3878, WX3880, WX3882, WX3884, WX3886,
         WX3888, WX3890, WX3892, WX3894, WX3896, WX3898, WX3900, WX3902,
         WX3904, WX3906, WX3908, WX3910, WX3912, WX4364, WX4363, WX4365,
         WX4367, WX4369, WX4371, WX4373, WX4375, WX4377, WX4379, WX4381,
         WX4383, WX4385, WX4387, WX4389, WX4391, WX4393, WX4395, WX4397,
         WX4399, WX4401, WX4403, WX4405, WX4407, WX4409, WX4411, WX4413,
         WX4415, WX4417, WX4419, WX4421, WX4423, WX4425, WX4523, WX4525,
         WX4527, WX4529, WX4531, WX4533, WX4535, WX4537, WX4539, WX4541,
         WX4543, WX4545, WX4547, WX4549, WX4551, WX4553, WX4556, WX4555,
         WX4558, WX4557, WX4560, WX4559, WX4562, WX4561, WX4564, WX4563,
         WX4566, WX4565, WX4568, WX4567, WX4570, WX4569, WX4572, WX4571,
         WX4574, WX4573, WX4576, WX4575, WX4578, WX4577, WX4580, WX4579,
         WX4582, WX4581, WX4584, WX4583, WX4585, WX4588, WX4587, WX4590,
         WX4589, WX4592, WX4591, WX4594, WX4593, WX4596, WX4595, WX4598,
         WX4597, WX4600, WX4599, WX4602, WX4601, WX4604, WX4603, WX4606,
         WX4605, WX4608, WX4607, WX4610, WX4609, WX4612, WX4611, WX4614,
         WX4613, WX4616, WX4615, WX4618, WX4617, WX4619, WX4622, WX4621,
         WX4624, WX4623, WX4626, WX4625, WX4628, WX4627, WX4630, WX4629,
         WX4632, WX4631, WX4634, WX4633, WX4636, WX4635, WX4638, WX4637,
         WX4640, WX4639, WX4642, WX4641, WX4644, WX4643, WX4646, WX4645,
         WX4648, WX4647, WX4650, WX4649, WX4652, WX4651, WX4653, WX4656,
         WX4655, WX4658, WX4657, WX4660, WX4659, WX4662, WX4661, WX4664,
         WX4663, WX4666, WX4665, WX4668, WX4667, WX4670, WX4669, WX4672,
         WX4671, WX4674, WX4673, WX4676, WX4675, WX4678, WX4677, WX4680,
         WX4679, WX4682, WX4681, WX4684, WX4683, WX4686, WX4685, WX4687,
         WX4690, WX4689, WX4692, WX4691, WX4694, WX4693, WX4696, WX4695,
         WX4698, WX4697, WX4700, WX4699, WX4702, WX4701, WX4704, WX4703,
         WX4706, WX4705, WX4708, WX4707, WX4710, WX4709, WX4712, WX4711,
         WX4714, WX4713, WX4716, WX4715, WX4718, WX4717, WX4720, WX4719,
         WX4721, WX4724, WX4723, WX4726, WX4725, WX4728, WX4727, WX4730,
         WX4729, WX4732, WX4731, WX4734, WX4733, WX4736, WX4735, WX4738,
         WX4737, WX4740, WX4739, WX4742, WX4741, WX4744, WX4743, WX4746,
         WX4745, WX4748, WX4747, WX4750, WX4749, WX4752, WX4751, WX4754,
         WX4753, WX4755, WX4758, WX4757, WX4760, WX4759, WX4762, WX4761,
         WX4764, WX4763, WX4766, WX4765, WX4768, WX4767, WX4770, WX4769,
         WX4772, WX4771, WX4774, WX4773, WX4776, WX4775, WX4778, WX4777,
         WX5143, WX5145, WX5147, WX5149, WX5151, WX5153, WX5155, WX5157,
         WX5159, WX5161, WX5163, WX5165, WX5167, WX5169, WX5171, WX5173,
         WX5175, WX5177, WX5179, WX5181, WX5183, WX5185, WX5187, WX5189,
         WX5191, WX5193, WX5195, WX5197, WX5199, WX5201, WX5203, WX5205,
         WX5657, WX5656, WX5658, WX5660, WX5662, WX5664, WX5666, WX5668,
         WX5670, WX5672, WX5674, WX5676, WX5678, WX5680, WX5682, WX5684,
         WX5686, WX5688, WX5690, WX5692, WX5694, WX5696, WX5698, WX5700,
         WX5702, WX5704, WX5706, WX5708, WX5710, WX5712, WX5714, WX5716,
         WX5718, WX5816, WX5818, WX5820, WX5822, WX5824, WX5826, WX5828,
         WX5830, WX5832, WX5834, WX5836, WX5838, WX5840, WX5842, WX5844,
         WX5846, WX5849, WX5848, WX5851, WX5850, WX5853, WX5852, WX5855,
         WX5854, WX5857, WX5856, WX5859, WX5858, WX5861, WX5860, WX5863,
         WX5862, WX5865, WX5864, WX5867, WX5866, WX5868, WX5871, WX5870,
         WX5873, WX5872, WX5875, WX5874, WX5877, WX5876, WX5879, WX5878,
         WX5881, WX5880, WX5883, WX5882, WX5885, WX5884, WX5887, WX5886,
         WX5889, WX5888, WX5891, WX5890, WX5893, WX5892, WX5895, WX5894,
         WX5897, WX5896, WX5899, WX5898, WX5901, WX5900, WX5902, WX5905,
         WX5904, WX5907, WX5906, WX5909, WX5908, WX5911, WX5910, WX5913,
         WX5912, WX5915, WX5914, WX5917, WX5916, WX5919, WX5918, WX5921,
         WX5920, WX5923, WX5922, WX5925, WX5924, WX5927, WX5926, WX5929,
         WX5928, WX5931, WX5930, WX5933, WX5932, WX5935, WX5934, WX5936,
         WX5939, WX5938, WX5941, WX5940, WX5943, WX5942, WX5945, WX5944,
         WX5947, WX5946, WX5949, WX5948, WX5951, WX5950, WX5953, WX5952,
         WX5955, WX5954, WX5957, WX5956, WX5959, WX5958, WX5961, WX5960,
         WX5963, WX5962, WX5965, WX5964, WX5967, WX5966, WX5969, WX5968,
         WX5970, WX5973, WX5972, WX5975, WX5974, WX5977, WX5976, WX5979,
         WX5978, WX5981, WX5980, WX5983, WX5982, WX5985, WX5984, WX5987,
         WX5986, WX5989, WX5988, WX5991, WX5990, WX5993, WX5992, WX5995,
         WX5994, WX5997, WX5996, WX5999, WX5998, WX6001, WX6000, WX6003,
         WX6002, WX6004, WX6007, WX6006, WX6009, WX6008, WX6011, WX6010,
         WX6013, WX6012, WX6015, WX6014, WX6017, WX6016, WX6019, WX6018,
         WX6021, WX6020, WX6023, WX6022, WX6025, WX6024, WX6027, WX6026,
         WX6029, WX6028, WX6031, WX6030, WX6033, WX6032, WX6035, WX6034,
         WX6037, WX6036, WX6038, WX6041, WX6040, WX6043, WX6042, WX6045,
         WX6044, WX6047, WX6046, WX6049, WX6048, WX6051, WX6050, WX6053,
         WX6052, WX6055, WX6054, WX6057, WX6056, WX6059, WX6058, WX6061,
         WX6060, WX6063, WX6062, WX6065, WX6064, WX6067, WX6066, WX6069,
         WX6068, WX6071, WX6070, WX6436, WX6438, WX6440, WX6442, WX6444,
         WX6446, WX6448, WX6450, WX6452, WX6454, WX6456, WX6458, WX6460,
         WX6462, WX6464, WX6466, WX6468, WX6470, WX6472, WX6474, WX6476,
         WX6478, WX6480, WX6482, WX6484, WX6486, WX6488, WX6490, WX6492,
         WX6494, WX6496, WX6498, WX6950, WX6949, WX6951, WX6953, WX6955,
         WX6957, WX6959, WX6961, WX6963, WX6965, WX6967, WX6969, WX6971,
         WX6973, WX6975, WX6977, WX6979, WX6981, WX6983, WX6985, WX6987,
         WX6989, WX6991, WX6993, WX6995, WX6997, WX6999, WX7001, WX7003,
         WX7005, WX7007, WX7009, WX7011, WX7109, WX7111, WX7113, WX7115,
         WX7117, WX7119, WX7121, WX7123, WX7125, WX7127, WX7129, WX7131,
         WX7133, WX7135, WX7137, WX7139, WX7142, WX7141, WX7144, WX7143,
         WX7146, WX7145, WX7148, WX7147, WX7150, WX7149, WX7151, WX7154,
         WX7153, WX7156, WX7155, WX7158, WX7157, WX7160, WX7159, WX7162,
         WX7161, WX7164, WX7163, WX7166, WX7165, WX7168, WX7167, WX7170,
         WX7169, WX7172, WX7171, WX7174, WX7173, WX7176, WX7175, WX7178,
         WX7177, WX7180, WX7179, WX7182, WX7181, WX7184, WX7183, WX7185,
         WX7188, WX7187, WX7190, WX7189, WX7192, WX7191, WX7194, WX7193,
         WX7196, WX7195, WX7198, WX7197, WX7200, WX7199, WX7202, WX7201,
         WX7204, WX7203, WX7206, WX7205, WX7208, WX7207, WX7210, WX7209,
         WX7212, WX7211, WX7214, WX7213, WX7216, WX7215, WX7218, WX7217,
         WX7219, WX7222, WX7221, WX7224, WX7223, WX7226, WX7225, WX7228,
         WX7227, WX7230, WX7229, WX7232, WX7231, WX7234, WX7233, WX7236,
         WX7235, WX7238, WX7237, WX7240, WX7239, WX7242, WX7241, WX7244,
         WX7243, WX7246, WX7245, WX7248, WX7247, WX7250, WX7249, WX7252,
         WX7251, WX7253, WX7256, WX7255, WX7258, WX7257, WX7260, WX7259,
         WX7262, WX7261, WX7264, WX7263, WX7266, WX7265, WX7268, WX7267,
         WX7270, WX7269, WX7272, WX7271, WX7274, WX7273, WX7276, WX7275,
         WX7278, WX7277, WX7280, WX7279, WX7282, WX7281, WX7284, WX7283,
         WX7286, WX7285, WX7287, WX7290, WX7289, WX7292, WX7291, WX7294,
         WX7293, WX7296, WX7295, WX7298, WX7297, WX7300, WX7299, WX7302,
         WX7301, WX7304, WX7303, WX7306, WX7305, WX7308, WX7307, WX7310,
         WX7309, WX7312, WX7311, WX7314, WX7313, WX7316, WX7315, WX7318,
         WX7317, WX7320, WX7319, WX7321, WX7324, WX7323, WX7326, WX7325,
         WX7328, WX7327, WX7330, WX7329, WX7332, WX7331, WX7334, WX7333,
         WX7336, WX7335, WX7338, WX7337, WX7340, WX7339, WX7342, WX7341,
         WX7344, WX7343, WX7346, WX7345, WX7348, WX7347, WX7350, WX7349,
         WX7352, WX7351, WX7354, WX7353, WX7355, WX7358, WX7357, WX7360,
         WX7359, WX7362, WX7361, WX7364, WX7363, WX7729, WX7731, WX7733,
         WX7735, WX7737, WX7739, WX7741, WX7743, WX7745, WX7747, WX7749,
         WX7751, WX7753, WX7755, WX7757, WX7759, WX7761, WX7763, WX7765,
         WX7767, WX7769, WX7771, WX7773, WX7775, WX7777, WX7779, WX7781,
         WX7783, WX7785, WX7787, WX7789, WX7791, WX8243, WX8242, WX8244,
         WX8246, WX8248, WX8250, WX8252, WX8254, WX8256, WX8258, WX8260,
         WX8262, WX8264, WX8266, WX8268, WX8270, WX8272, WX8274, WX8276,
         WX8278, WX8280, WX8282, WX8284, WX8286, WX8288, WX8290, WX8292,
         WX8294, WX8296, WX8298, WX8300, WX8302, WX8304, WX8402, WX8404,
         WX8406, WX8408, WX8410, WX8412, WX8414, WX8416, WX8418, WX8420,
         WX8422, WX8424, WX8426, WX8428, WX8430, WX8432, WX8434, WX8437,
         WX8436, WX8439, WX8438, WX8441, WX8440, WX8443, WX8442, WX8445,
         WX8444, WX8447, WX8446, WX8449, WX8448, WX8451, WX8450, WX8453,
         WX8452, WX8455, WX8454, WX8457, WX8456, WX8459, WX8458, WX8461,
         WX8460, WX8463, WX8462, WX8465, WX8464, WX8467, WX8466, WX8468,
         WX8471, WX8470, WX8473, WX8472, WX8475, WX8474, WX8477, WX8476,
         WX8479, WX8478, WX8481, WX8480, WX8483, WX8482, WX8485, WX8484,
         WX8487, WX8486, WX8489, WX8488, WX8491, WX8490, WX8493, WX8492,
         WX8495, WX8494, WX8497, WX8496, WX8499, WX8498, WX8501, WX8500,
         WX8502, WX8505, WX8504, WX8507, WX8506, WX8509, WX8508, WX8511,
         WX8510, WX8513, WX8512, WX8515, WX8514, WX8517, WX8516, WX8519,
         WX8518, WX8521, WX8520, WX8523, WX8522, WX8525, WX8524, WX8527,
         WX8526, WX8529, WX8528, WX8531, WX8530, WX8533, WX8532, WX8535,
         WX8534, WX8536, WX8539, WX8538, WX8541, WX8540, WX8543, WX8542,
         WX8545, WX8544, WX8547, WX8546, WX8549, WX8548, WX8551, WX8550,
         WX8553, WX8552, WX8555, WX8554, WX8557, WX8556, WX8559, WX8558,
         WX8561, WX8560, WX8563, WX8562, WX8565, WX8564, WX8567, WX8566,
         WX8569, WX8568, WX8570, WX8573, WX8572, WX8575, WX8574, WX8577,
         WX8576, WX8579, WX8578, WX8581, WX8580, WX8583, WX8582, WX8585,
         WX8584, WX8587, WX8586, WX8589, WX8588, WX8591, WX8590, WX8593,
         WX8592, WX8595, WX8594, WX8597, WX8596, WX8599, WX8598, WX8601,
         WX8600, WX8603, WX8602, WX8604, WX8607, WX8606, WX8609, WX8608,
         WX8611, WX8610, WX8613, WX8612, WX8615, WX8614, WX8617, WX8616,
         WX8619, WX8618, WX8621, WX8620, WX8623, WX8622, WX8625, WX8624,
         WX8627, WX8626, WX8629, WX8628, WX8631, WX8630, WX8633, WX8632,
         WX8635, WX8634, WX8637, WX8636, WX8638, WX8641, WX8640, WX8643,
         WX8642, WX8645, WX8644, WX8647, WX8646, WX8649, WX8648, WX8651,
         WX8650, WX8653, WX8652, WX8655, WX8654, WX8657, WX8656, WX9022,
         WX9024, WX9026, WX9028, WX9030, WX9032, WX9034, WX9036, WX9038,
         WX9040, WX9042, WX9044, WX9046, WX9048, WX9050, WX9052, WX9054,
         WX9056, WX9058, WX9060, WX9062, WX9064, WX9066, WX9068, WX9070,
         WX9072, WX9074, WX9076, WX9078, WX9080, WX9082, WX9084, WX9536,
         WX9535, WX9537, WX9539, WX9541, WX9543, WX9545, WX9547, WX9549,
         WX9551, WX9553, WX9555, WX9557, WX9559, WX9561, WX9563, WX9565,
         WX9567, WX9569, WX9571, WX9573, WX9575, WX9577, WX9579, WX9581,
         WX9583, WX9585, WX9587, WX9589, WX9591, WX9593, WX9595, WX9597,
         WX9695, WX9697, WX9699, WX9701, WX9703, WX9705, WX9707, WX9709,
         WX9711, WX9713, WX9715, WX9717, WX9719, WX9721, WX9723, WX9725,
         WX9728, WX9727, WX9730, WX9729, WX9732, WX9731, WX9734, WX9733,
         WX9736, WX9735, WX9738, WX9737, WX9740, WX9739, WX9742, WX9741,
         WX9744, WX9743, WX9746, WX9745, WX9748, WX9747, WX9750, WX9749,
         WX9751, WX9754, WX9753, WX9756, WX9755, WX9758, WX9757, WX9760,
         WX9759, WX9762, WX9761, WX9764, WX9763, WX9766, WX9765, WX9768,
         WX9767, WX9770, WX9769, WX9772, WX9771, WX9774, WX9773, WX9776,
         WX9775, WX9778, WX9777, WX9780, WX9779, WX9782, WX9781, WX9784,
         WX9783, WX9785, WX9788, WX9787, WX9790, WX9789, WX9792, WX9791,
         WX9794, WX9793, WX9796, WX9795, WX9798, WX9797, WX9800, WX9799,
         WX9802, WX9801, WX9804, WX9803, WX9806, WX9805, WX9808, WX9807,
         WX9810, WX9809, WX9812, WX9811, WX9814, WX9813, WX9816, WX9815,
         WX9818, WX9817, WX9819, WX9822, WX9821, WX9824, WX9823, WX9826,
         WX9825, WX9828, WX9827, WX9830, WX9829, WX9832, WX9831, WX9834,
         WX9833, WX9836, WX9835, WX9838, WX9837, WX9840, WX9839, WX9842,
         WX9841, WX9844, WX9843, WX9846, WX9845, WX9848, WX9847, WX9850,
         WX9849, WX9852, WX9851, WX9853, WX9856, WX9855, WX9858, WX9857,
         WX9860, WX9859, WX9862, WX9861, WX9864, WX9863, WX9866, WX9865,
         WX9868, WX9867, WX9870, WX9869, WX9872, WX9871, WX9874, WX9873,
         WX9876, WX9875, WX9878, WX9877, WX9880, WX9879, WX9882, WX9881,
         WX9884, WX9883, WX9886, WX9885, WX9887, WX9890, WX9889, WX9892,
         WX9891, WX9894, WX9893, WX9896, WX9895, WX9898, WX9897, WX9900,
         WX9899, WX9902, WX9901, WX9904, WX9903, WX9906, WX9905, WX9908,
         WX9907, WX9910, WX9909, WX9912, WX9911, WX9914, WX9913, WX9916,
         WX9915, WX9918, WX9917, WX9920, WX9919, WX9921, WX9924, WX9923,
         WX9926, WX9925, WX9928, WX9927, WX9930, WX9929, WX9932, WX9931,
         WX9934, WX9933, WX9936, WX9935, WX9938, WX9937, WX9940, WX9939,
         WX9942, WX9941, WX9944, WX9943, WX9946, WX9945, WX9948, WX9947,
         WX9950, WX9949, WX10315, WX10317, WX10319, WX10321, WX10323, WX10325,
         WX10327, WX10329, WX10331, WX10333, WX10335, WX10337, WX10339,
         WX10341, WX10343, WX10345, WX10347, WX10349, WX10351, WX10353,
         WX10355, WX10357, WX10359, WX10361, WX10363, WX10365, WX10367,
         WX10369, WX10371, WX10373, WX10375, WX10377, WX10829, WX10828,
         WX10830, WX10832, WX10834, WX10836, WX10838, WX10840, WX10842,
         WX10844, WX10846, WX10848, WX10850, WX10852, WX10854, WX10856,
         WX10858, WX10860, WX10862, WX10864, WX10866, WX10868, WX10870,
         WX10872, WX10874, WX10876, WX10878, WX10880, WX10882, WX10884,
         WX10886, WX10888, WX10890, WX10988, WX10990, WX10992, WX10994,
         WX10996, WX10998, WX11000, WX11002, WX11004, WX11006, WX11008,
         WX11010, WX11012, WX11014, WX11016, WX11018, WX11021, WX11020,
         WX11023, WX11022, WX11025, WX11024, WX11027, WX11026, WX11029,
         WX11028, WX11031, WX11030, WX11033, WX11032, WX11034, WX11037,
         WX11036, WX11039, WX11038, WX11041, WX11040, WX11043, WX11042,
         WX11045, WX11044, WX11047, WX11046, WX11049, WX11048, WX11051,
         WX11050, WX11053, WX11052, WX11055, WX11054, WX11057, WX11056,
         WX11059, WX11058, WX11061, WX11060, WX11063, WX11062, WX11065,
         WX11064, WX11067, WX11066, WX11068, WX11071, WX11070, WX11073,
         WX11072, WX11075, WX11074, WX11077, WX11076, WX11079, WX11078,
         WX11081, WX11080, WX11083, WX11082, WX11085, WX11084, WX11087,
         WX11086, WX11089, WX11088, WX11091, WX11090, WX11093, WX11092,
         WX11095, WX11094, WX11097, WX11096, WX11099, WX11098, WX11101,
         WX11100, WX11102, WX11105, WX11104, WX11107, WX11106, WX11109,
         WX11108, WX11111, WX11110, WX11113, WX11112, WX11115, WX11114,
         WX11117, WX11116, WX11119, WX11118, WX11121, WX11120, WX11123,
         WX11122, WX11125, WX11124, WX11127, WX11126, WX11129, WX11128,
         WX11131, WX11130, WX11133, WX11132, WX11135, WX11134, WX11136,
         WX11139, WX11138, WX11141, WX11140, WX11143, WX11142, WX11145,
         WX11144, WX11147, WX11146, WX11149, WX11148, WX11151, WX11150,
         WX11153, WX11152, WX11155, WX11155_Tj_Payload, WX11154, WX11157, WX11156, WX11159,
         WX11158, WX11161, WX11160, WX11163, WX11162, WX11165, WX11164,
         WX11167, WX11166, WX11169, WX11168, WX11170, WX11173, WX11172,
         WX11175, WX11174, WX11177, WX11176, WX11179, WX11178, WX11181,
         WX11180, WX11183, WX11182, WX11185, WX11184, WX11187, WX11186,
         WX11189, WX11188, WX11191, WX11190, WX11193, WX11192, WX11195,
         WX11194, WX11197, WX11196, WX11199, WX11198, WX11201, WX11200,
         WX11203, WX11202, WX11204, WX11207, WX11206, WX11209, WX11208,
         WX11211, WX11210, WX11213, WX11212, WX11215, WX11214, WX11217,
         WX11216, WX11219, WX11218, WX11221, WX11220, WX11223, WX11222,
         WX11225, WX11224, WX11227, WX11226, WX11229, WX11228, WX11231,
         WX11230, WX11233, WX11232, WX11235, WX11234, WX11237, WX11236,
         WX11238, WX11241, WX11240, WX11243, WX11242, WX11608, WX11610,
         WX11612, WX11614, WX11616, WX11618, WX11620, WX11622, WX11624,
         WX11626, WX11628, WX11630, WX11632, WX11634, WX11636, WX11638,
         WX11640, WX11642, WX11644, WX11646, WX11648, WX11650, WX11652,
         WX11654, WX11656, WX11658, WX11660, WX11662, WX11664, WX11666,
         WX11668, WX11670, DFF_160_n1, DFF_161_n1, DFF_162_n1, DFF_163_n1,
         DFF_164_n1, DFF_165_n1, DFF_166_n1, DFF_167_n1, DFF_168_n1,
         DFF_169_n1, DFF_170_n1, DFF_171_n1, DFF_172_n1, DFF_173_n1,
         DFF_174_n1, DFF_175_n1, DFF_176_n1, DFF_177_n1, DFF_178_n1,
         DFF_179_n1, DFF_180_n1, DFF_181_n1, DFF_182_n1, DFF_183_n1,
         DFF_184_n1, DFF_185_n1, DFF_186_n1, DFF_187_n1, DFF_188_n1,
         DFF_189_n1, DFF_190_n1, DFF_191_n1, DFF_352_n1, DFF_353_n1,
         DFF_354_n1, DFF_355_n1, DFF_356_n1, DFF_357_n1, DFF_358_n1,
         DFF_359_n1, DFF_360_n1, DFF_361_n1, DFF_362_n1, DFF_363_n1,
         DFF_364_n1, DFF_365_n1, DFF_366_n1, DFF_367_n1, DFF_368_n1,
         DFF_369_n1, DFF_370_n1, DFF_371_n1, DFF_372_n1, DFF_373_n1,
         DFF_374_n1, DFF_375_n1, DFF_376_n1, DFF_377_n1, DFF_378_n1,
         DFF_379_n1, DFF_380_n1, DFF_381_n1, DFF_382_n1, DFF_383_n1,
         DFF_544_n1, DFF_545_n1, DFF_546_n1, DFF_547_n1, DFF_548_n1,
         DFF_549_n1, DFF_550_n1, DFF_551_n1, DFF_552_n1, DFF_553_n1,
         DFF_554_n1, DFF_555_n1, DFF_556_n1, DFF_557_n1, DFF_558_n1,
         DFF_559_n1, DFF_560_n1, DFF_561_n1, DFF_562_n1, DFF_563_n1,
         DFF_564_n1, DFF_565_n1, DFF_566_n1, DFF_567_n1, DFF_568_n1,
         DFF_569_n1, DFF_570_n1, DFF_571_n1, DFF_572_n1, DFF_573_n1,
         DFF_574_n1, DFF_575_n1, DFF_736_n1, DFF_737_n1, DFF_738_n1,
         DFF_739_n1, DFF_740_n1, DFF_741_n1, DFF_742_n1, DFF_743_n1,
         DFF_744_n1, DFF_745_n1, DFF_746_n1, DFF_747_n1, DFF_748_n1,
         DFF_749_n1, DFF_750_n1, DFF_751_n1, DFF_752_n1, DFF_753_n1,
         DFF_754_n1, DFF_755_n1, DFF_756_n1, DFF_757_n1, DFF_758_n1,
         DFF_759_n1, DFF_760_n1, DFF_761_n1, DFF_762_n1, DFF_763_n1,
         DFF_764_n1, DFF_765_n1, DFF_766_n1, DFF_767_n1, DFF_928_n1,
         DFF_929_n1, DFF_930_n1, DFF_931_n1, DFF_932_n1, DFF_933_n1,
         DFF_934_n1, DFF_935_n1, DFF_936_n1, DFF_937_n1, DFF_938_n1,
         DFF_939_n1, DFF_940_n1, DFF_941_n1, DFF_942_n1, DFF_943_n1,
         DFF_944_n1, DFF_945_n1, DFF_946_n1, DFF_947_n1, DFF_948_n1,
         DFF_949_n1, DFF_950_n1, DFF_951_n1, DFF_952_n1, DFF_953_n1,
         DFF_954_n1, DFF_955_n1, DFF_956_n1, DFF_957_n1, DFF_958_n1,
         DFF_959_n1, DFF_1120_n1, DFF_1121_n1, DFF_1122_n1, DFF_1123_n1,
         DFF_1124_n1, DFF_1125_n1, DFF_1126_n1, DFF_1127_n1, DFF_1128_n1,
         DFF_1129_n1, DFF_1130_n1, DFF_1131_n1, DFF_1132_n1, DFF_1133_n1,
         DFF_1134_n1, DFF_1135_n1, DFF_1136_n1, DFF_1137_n1, DFF_1138_n1,
         DFF_1139_n1, DFF_1140_n1, DFF_1141_n1, DFF_1142_n1, DFF_1143_n1,
         DFF_1144_n1, DFF_1145_n1, DFF_1146_n1, DFF_1147_n1, DFF_1148_n1,
         DFF_1149_n1, DFF_1150_n1, DFF_1151_n1, DFF_1312_n1, DFF_1313_n1,
         DFF_1314_n1, DFF_1315_n1, DFF_1316_n1, DFF_1317_n1, DFF_1318_n1,
         DFF_1319_n1, DFF_1320_n1, DFF_1321_n1, DFF_1322_n1, DFF_1323_n1,
         DFF_1324_n1, DFF_1325_n1, DFF_1326_n1, DFF_1327_n1, DFF_1328_n1,
         DFF_1329_n1, DFF_1330_n1, DFF_1331_n1, DFF_1332_n1, DFF_1333_n1,
         DFF_1334_n1, DFF_1335_n1, DFF_1336_n1, DFF_1337_n1, DFF_1338_n1,
         DFF_1339_n1, DFF_1340_n1, DFF_1341_n1, DFF_1342_n1, DFF_1343_n1,
         DFF_1504_n1, DFF_1505_n1, DFF_1506_n1, DFF_1507_n1, DFF_1508_n1,
         DFF_1509_n1, DFF_1510_n1, DFF_1511_n1, DFF_1512_n1, DFF_1513_n1,
         DFF_1514_n1, DFF_1515_n1, DFF_1516_n1, DFF_1517_n1, DFF_1518_n1,
         DFF_1519_n1, DFF_1520_n1, DFF_1521_n1, DFF_1522_n1, DFF_1523_n1,
         DFF_1524_n1, DFF_1525_n1, DFF_1526_n1, DFF_1527_n1, DFF_1528_n1,
         DFF_1529_n1, DFF_1530_n1, DFF_1531_n1, DFF_1532_n1, DFF_1533_n1,
         DFF_1534_n1, DFF_1535_n1, DFF_1696_n1, DFF_1697_n1, DFF_1698_n1,
         DFF_1699_n1, DFF_1700_n1, DFF_1701_n1, DFF_1702_n1, DFF_1703_n1,
         DFF_1704_n1, DFF_1705_n1, DFF_1706_n1, DFF_1707_n1, DFF_1708_n1,
         DFF_1709_n1, DFF_1710_n1, DFF_1711_n1, DFF_1712_n1, DFF_1713_n1,
         DFF_1714_n1, DFF_1715_n1, DFF_1716_n1, DFF_1717_n1, DFF_1718_n1,
         DFF_1719_n1, DFF_1720_n1, DFF_1721_n1, DFF_1722_n1, DFF_1723_n1,
         DFF_1724_n1, DFF_1725_n1, DFF_1726_n1, DFF_1727_n1, n1729, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2284, n2285, n2287, n2288, n2290, n2291,
         n2293, n2294, n2296, n2297, n2299, n2300, n2302, n2303, n2305, n2306,
         n2308, n2309, n2311, n2312, n2314, n2315, n2317, n2318, n2320, n2321,
         n2323, n2324, n2326, n2327, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2412, n2413, n2415, n2416,
         n2418, n2419, n2421, n2422, n2424, n2425, n2427, n2428, n2430, n2431,
         n2433, n2434, n2436, n2437, n2439, n2440, n2442, n2443, n2445, n2446,
         n2448, n2449, n2451, n2452, n2454, n2455, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2636, n2637, n2639, n2640, n2642, n2643,
         n2645, n2646, n2648, n2649, n2651, n2652, n2654, n2655, n2657, n2658,
         n2660, n2661, n2663, n2664, n2666, n2667, n2669, n2670, n2672, n2673,
         n2675, n2676, n2678, n2679, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2764, n2765, n2767, n2768,
         n2770, n2771, n2773, n2774, n2776, n2777, n2779, n2780, n2782, n2783,
         n2785, n2786, n2788, n2789, n2791, n2792, n2794, n2795, n2797, n2798,
         n2800, n2801, n2803, n2804, n2806, n2807, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2892, n2893,
         n2895, n2896, n2898, n2899, n2901, n2902, n2904, n2905, n2907, n2908,
         n2910, n2911, n2913, n2914, n2916, n2917, n2919, n2920, n2922, n2923,
         n2925, n2926, n2928, n2929, n2931, n2932, n2934, n2935, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3020,
         n3023, n3026, n3029, n3032, n3035, n3038, n3041, n3044, n3047, n3050,
         n3053, n3056, n3059, n3062, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3147, n3149, n3151, n3153, n3155,
         n3157, n3159, n3161, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3199, n3201, n3203,
         n3205, n3207, n3209, n3211, n3213, n3215, n3217, n3219, n3221, n3223,
         n3225, n3227, n3229, n3231, n3233, n3235, n3237, n3239, n3241, n3243,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3282, n3284, n3286, n3288, n3290,
         n3292, n3294, n3296, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3332, n3334, n3336, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8293, n8294, n8295, n8304, n8305, n8306, n8307,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8470, n8479,
         n8480, n8481, n8482, n8483, n8484, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8523, n8524, n8525,
         n8526, n8527, n8528, n8537, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8653, n8654, n8655, n8656, n8657, n8658, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8699, n8700, n8701, n8702;
  assign test_so99 = CRC_OUT_1_14;
  assign test_so100 = CRC_OUT_1_31;
  assign test_so88 = CRC_OUT_2_19;
  assign test_so87 = CRC_OUT_2_2;
  assign test_so77 = CRC_OUT_3_24;
  assign test_so76 = CRC_OUT_3_7;
  assign test_so65 = CRC_OUT_4_12;
  assign test_so66 = CRC_OUT_4_29;
  assign test_so53 = CRC_OUT_5_0;
  assign test_so54 = CRC_OUT_5_17;
  assign test_so43 = CRC_OUT_6_22;
  assign test_so42 = CRC_OUT_6_5;
  assign test_so31 = CRC_OUT_7_10;
  assign test_so32 = CRC_OUT_7_27;
  assign test_so21 = CRC_OUT_8_25;
  assign test_so20 = CRC_OUT_8_7;
  assign test_so9 = CRC_OUT_9_1;
  assign test_so10 = CRC_OUT_9_19;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(test_se), .CLK(CK), .Q(
        WX485), .QN() );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(test_se), .CLK(CK), .Q(WX487), .QN() );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(test_se), .CLK(CK), .Q(WX489), .QN() );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(test_se), .CLK(CK), .Q(WX491), .QN() );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(test_se), .CLK(CK), .Q(WX493), .QN() );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(test_se), .CLK(CK), .Q(WX495), .QN() );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(test_se), .CLK(CK), .Q(WX497), .QN() );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(test_se), .CLK(CK), .Q(WX499), .QN() );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(test_se), .CLK(CK), .Q(WX501), .QN() );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(test_se), .CLK(CK), .Q(WX503), .QN() );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(test_se), .CLK(CK), .Q(
        WX505), .QN() );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(test_se), .CLK(CK), .Q(
        WX507), .QN() );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(test_se), .CLK(CK), .Q(
        WX509), .QN() );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(test_se), .CLK(CK), .Q(
        WX511), .QN() );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(test_se), .CLK(CK), .Q(
        WX513), .QN() );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(test_se), .CLK(CK), .Q(
        WX515), .QN() );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(test_se), .CLK(CK), .Q(
        WX517), .QN() );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(test_se), .CLK(CK), .Q(
        test_so1), .QN() );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(test_se), .CLK(CK), .Q(
        WX521), .QN() );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(test_se), .CLK(CK), .Q(
        WX523), .QN() );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(test_se), .CLK(CK), .Q(
        WX525), .QN() );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(test_se), .CLK(CK), .Q(
        WX527), .QN() );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(test_se), .CLK(CK), .Q(
        WX529), .QN() );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(test_se), .CLK(CK), .Q(
        WX531), .QN() );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(test_se), .CLK(CK), .Q(
        WX533), .QN() );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(test_se), .CLK(CK), .Q(
        WX535), .QN() );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(test_se), .CLK(CK), .Q(
        WX537), .QN() );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(test_se), .CLK(CK), .Q(
        WX539), .QN() );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(test_se), .CLK(CK), .Q(
        WX541), .QN() );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(test_se), .CLK(CK), .Q(
        WX543), .QN() );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(test_se), .CLK(CK), .Q(
        WX545), .QN() );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(test_se), .CLK(CK), .Q(
        WX547), .QN() );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(test_se), .CLK(CK), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(test_se), .CLK(CK), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(test_se), .CLK(CK), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(test_se), .CLK(CK), .Q(
        test_so2), .QN(n3523) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(test_se), .CLK(CK), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(test_se), .CLK(CK), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(test_se), .CLK(CK), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(test_se), .CLK(CK), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(test_se), .CLK(CK), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(test_se), .CLK(CK), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(test_se), .CLK(CK), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(test_se), .CLK(CK), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(test_se), .CLK(CK), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(test_se), .CLK(CK), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(test_se), .CLK(CK), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(test_se), .CLK(CK), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(test_se), .CLK(CK), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(test_se), .CLK(CK), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(test_se), .CLK(CK), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(test_se), .CLK(CK), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(test_se), .CLK(CK), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(test_se), .CLK(CK), .Q(
        test_so3), .QN(n3487) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(test_se), .CLK(CK), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(test_se), .CLK(CK), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(test_se), .CLK(CK), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(test_se), .CLK(CK), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(test_se), .CLK(CK), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(test_se), .CLK(CK), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(test_se), .CLK(CK), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(test_se), .CLK(CK), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(test_se), .CLK(CK), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(test_se), .CLK(CK), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(test_se), .CLK(CK), .Q(
        WX709), .QN() );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(test_se), .CLK(CK), .Q(
        WX711), .QN() );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(test_se), .CLK(CK), .Q(
        WX713), .QN() );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(test_se), .CLK(CK), .Q(
        WX715), .QN() );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(test_se), .CLK(CK), .Q(
        WX717), .QN() );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(test_se), .CLK(CK), .Q(
        WX719), .QN() );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(test_se), .CLK(CK), .Q(
        WX721), .QN() );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(test_se), .CLK(CK), .Q(
        test_so4), .QN() );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(test_se), .CLK(CK), .Q(
        WX725), .QN() );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(test_se), .CLK(CK), .Q(
        WX727), .QN() );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(test_se), .CLK(CK), .Q(
        WX729), .QN() );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(test_se), .CLK(CK), .Q(
        WX731), .QN() );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(test_se), .CLK(CK), .Q(
        WX733), .QN() );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(test_se), .CLK(CK), .Q(
        WX735), .QN() );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(test_se), .CLK(CK), .Q(
        WX737), .QN() );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(test_se), .CLK(CK), .Q(
        WX739), .QN() );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(test_se), .CLK(CK), .Q(
        WX741), .QN() );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(test_se), .CLK(CK), .Q(
        WX743), .QN() );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(test_se), .CLK(CK), .Q(
        WX745), .QN() );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(test_se), .CLK(CK), .Q(
        WX747), .QN() );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(test_se), .CLK(CK), .Q(
        WX749), .QN() );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(test_se), .CLK(CK), .Q(
        WX751), .QN() );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(test_se), .CLK(CK), .Q(
        WX753), .QN() );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(test_se), .CLK(CK), .Q(
        WX755), .QN() );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(test_se), .CLK(CK), .Q(
        WX757), .QN() );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(test_se), .CLK(CK), .Q(
        test_so5), .QN() );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(test_se), .CLK(CK), .Q(
        WX761), .QN() );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(test_se), .CLK(CK), .Q(
        WX763), .QN() );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(test_se), .CLK(CK), .Q(
        WX765), .QN() );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(test_se), .CLK(CK), .Q(
        WX767), .QN() );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(test_se), .CLK(CK), .Q(
        WX769), .QN() );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(test_se), .CLK(CK), .Q(
        WX771), .QN() );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(test_se), .CLK(CK), .Q(
        WX773), .QN() );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(test_se), .CLK(CK), .Q(
        WX775), .QN() );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(test_se), .CLK(CK), .Q(
        WX777), .QN() );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(test_se), .CLK(CK), .Q(
        WX779), .QN() );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(test_se), .CLK(CK), .Q(
        WX781), .QN() );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(test_se), .CLK(CK), .Q(
        WX783), .QN() );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(test_se), .CLK(CK), .Q(
        WX785), .QN() );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(test_se), .CLK(CK), .Q(
        WX787), .QN() );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(test_se), .CLK(CK), .Q(
        WX789), .QN() );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(test_se), .CLK(CK), .Q(
        WX791), .QN() );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(test_se), .CLK(CK), .Q(
        WX793), .QN() );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(test_se), .CLK(CK), .Q(
        test_so6), .QN() );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(test_se), .CLK(CK), .Q(
        WX797), .QN() );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(test_se), .CLK(CK), .Q(
        WX799), .QN() );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(test_se), .CLK(CK), .Q(
        WX801), .QN() );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(test_se), .CLK(CK), .Q(
        WX803), .QN() );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(test_se), .CLK(CK), .Q(
        WX805), .QN() );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(test_se), .CLK(CK), .Q(
        WX807), .QN() );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(test_se), .CLK(CK), .Q(
        WX809), .QN() );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(test_se), .CLK(CK), .Q(
        WX811), .QN() );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(test_se), .CLK(CK), .Q(
        WX813), .QN() );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(test_se), .CLK(CK), .Q(
        WX815), .QN() );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(test_se), .CLK(CK), .Q(
        WX817), .QN() );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(test_se), .CLK(CK), .Q(
        WX819), .QN() );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(test_se), .CLK(CK), .Q(
        WX821), .QN() );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(test_se), .CLK(CK), .Q(
        WX823), .QN() );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(test_se), .CLK(CK), .Q(
        WX825), .QN() );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(test_se), .CLK(CK), .Q(
        WX827), .QN() );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(test_se), .CLK(CK), .Q(
        WX829), .QN() );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(test_se), .CLK(CK), .Q(
        test_so7), .QN() );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(test_se), .CLK(CK), .Q(
        WX833), .QN() );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(test_se), .CLK(CK), .Q(
        WX835), .QN() );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(test_se), .CLK(CK), .Q(
        WX837), .QN() );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(test_se), .CLK(CK), .Q(
        WX839), .QN() );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(test_se), .CLK(CK), .Q(
        WX841), .QN() );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(test_se), .CLK(CK), .Q(
        WX843), .QN() );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(test_se), .CLK(CK), .Q(
        WX845), .QN() );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(test_se), .CLK(CK), .Q(
        WX847), .QN() );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(test_se), .CLK(CK), .Q(
        WX849), .QN() );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(test_se), .CLK(CK), .Q(
        WX851), .QN() );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(test_se), .CLK(CK), .Q(
        WX853), .QN() );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(test_se), .CLK(CK), .Q(
        WX855), .QN() );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(test_se), .CLK(CK), .Q(
        WX857), .QN() );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(test_se), .CLK(CK), .Q(
        WX859), .QN() );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(test_se), .CLK(CK), .Q(
        WX861), .QN() );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(test_se), .CLK(CK), .Q(
        WX863), .QN() );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(test_se), .CLK(CK), .Q(
        WX865), .QN() );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(test_se), .CLK(CK), .Q(
        test_so8), .QN() );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(test_se), .CLK(CK), .Q(
        WX869), .QN() );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(test_se), .CLK(CK), .Q(
        WX871), .QN() );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(test_se), .CLK(CK), .Q(
        WX873), .QN() );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(test_se), .CLK(CK), .Q(
        WX875), .QN() );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(test_se), .CLK(CK), .Q(
        WX877), .QN() );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(test_se), .CLK(CK), .Q(
        WX879), .QN() );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(test_se), .CLK(CK), .Q(
        WX881), .QN() );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(test_se), .CLK(CK), .Q(
        WX883), .QN() );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(test_se), .CLK(CK), .Q(
        WX885), .QN() );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(test_se), .CLK(CK), .Q(
        WX887), .QN() );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(test_se), .CLK(CK), .Q(
        WX889), .QN() );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(test_se), .CLK(CK), .Q(
        WX891), .QN() );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(test_se), .CLK(CK), .Q(
        WX893), .QN() );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(test_se), .CLK(CK), .Q(
        WX895), .QN() );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(test_se), .CLK(CK), .Q(
        WX897), .QN() );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(test_se), .CLK(CK), .Q(
        WX899), .QN() );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_1), .QN(DFF_161_n1) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_19), .QN(DFF_179_n1) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(WX1777), .SI(CRC_OUT_9_31), .SE(test_se), .CLK(CK), 
        .Q(WX1778), .QN() );
  SDFFX1 DFF_193_Q_reg ( .D(WX1779), .SI(WX1778), .SE(test_se), .CLK(CK), .Q(
        n8702), .QN(n4033) );
  SDFFX1 DFF_194_Q_reg ( .D(WX1781), .SI(n8702), .SE(test_se), .CLK(CK), .Q(
        n8701), .QN(n4032) );
  SDFFX1 DFF_195_Q_reg ( .D(WX1783), .SI(n8701), .SE(test_se), .CLK(CK), .Q(
        n8700), .QN(n4031) );
  SDFFX1 DFF_196_Q_reg ( .D(WX1785), .SI(n8700), .SE(test_se), .CLK(CK), .Q(
        n8699), .QN(n4030) );
  SDFFX1 DFF_197_Q_reg ( .D(WX1787), .SI(n8699), .SE(test_se), .CLK(CK), .Q(
        test_so11), .QN(n4029) );
  SDFFX1 DFF_198_Q_reg ( .D(WX1789), .SI(test_si12), .SE(test_se), .CLK(CK), 
        .Q(n8696), .QN(n4028) );
  SDFFX1 DFF_199_Q_reg ( .D(WX1791), .SI(n8696), .SE(test_se), .CLK(CK), .Q(
        n8695), .QN(n4027) );
  SDFFX1 DFF_200_Q_reg ( .D(WX1793), .SI(n8695), .SE(test_se), .CLK(CK), .Q(
        n8694), .QN(n4026) );
  SDFFX1 DFF_201_Q_reg ( .D(WX1795), .SI(n8694), .SE(test_se), .CLK(CK), .Q(
        n8693), .QN(n4025) );
  SDFFX1 DFF_202_Q_reg ( .D(WX1797), .SI(n8693), .SE(test_se), .CLK(CK), .Q(
        n8692), .QN(n4024) );
  SDFFX1 DFF_203_Q_reg ( .D(WX1799), .SI(n8692), .SE(test_se), .CLK(CK), .Q(
        n8691), .QN(n4023) );
  SDFFX1 DFF_204_Q_reg ( .D(WX1801), .SI(n8691), .SE(test_se), .CLK(CK), .Q(
        n8690), .QN(n4022) );
  SDFFX1 DFF_205_Q_reg ( .D(WX1803), .SI(n8690), .SE(test_se), .CLK(CK), .Q(
        n8689), .QN(n4021) );
  SDFFX1 DFF_206_Q_reg ( .D(WX1805), .SI(n8689), .SE(test_se), .CLK(CK), .Q(
        n8688), .QN(n4020) );
  SDFFX1 DFF_207_Q_reg ( .D(WX1807), .SI(n8688), .SE(test_se), .CLK(CK), .Q(
        n8687), .QN(n4019) );
  SDFFX1 DFF_208_Q_reg ( .D(WX1809), .SI(n8687), .SE(test_se), .CLK(CK), .Q(
        n8686), .QN(n4018) );
  SDFFX1 DFF_209_Q_reg ( .D(WX1811), .SI(n8686), .SE(test_se), .CLK(CK), .Q(
        n8685), .QN(n4017) );
  SDFFX1 DFF_210_Q_reg ( .D(WX1813), .SI(n8685), .SE(test_se), .CLK(CK), .Q(
        n8684), .QN(n4016) );
  SDFFX1 DFF_211_Q_reg ( .D(WX1815), .SI(n8684), .SE(test_se), .CLK(CK), .Q(
        n8683), .QN(n4015) );
  SDFFX1 DFF_212_Q_reg ( .D(WX1817), .SI(n8683), .SE(test_se), .CLK(CK), .Q(
        n8682), .QN(n4014) );
  SDFFX1 DFF_213_Q_reg ( .D(WX1819), .SI(n8682), .SE(test_se), .CLK(CK), .Q(
        n8681), .QN(n4013) );
  SDFFX1 DFF_214_Q_reg ( .D(WX1821), .SI(n8681), .SE(test_se), .CLK(CK), .Q(
        n8680), .QN(n4012) );
  SDFFX1 DFF_215_Q_reg ( .D(WX1823), .SI(n8680), .SE(test_se), .CLK(CK), .Q(
        test_so12), .QN(n4011) );
  SDFFX1 DFF_216_Q_reg ( .D(WX1825), .SI(test_si13), .SE(test_se), .CLK(CK), 
        .Q(n8677), .QN(n4010) );
  SDFFX1 DFF_217_Q_reg ( .D(WX1827), .SI(n8677), .SE(test_se), .CLK(CK), .Q(
        n8676), .QN(n4009) );
  SDFFX1 DFF_218_Q_reg ( .D(WX1829), .SI(n8676), .SE(test_se), .CLK(CK), .Q(
        n8675), .QN(n4008) );
  SDFFX1 DFF_219_Q_reg ( .D(WX1831), .SI(n8675), .SE(test_se), .CLK(CK), .Q(
        n8674), .QN(n4007) );
  SDFFX1 DFF_220_Q_reg ( .D(WX1833), .SI(n8674), .SE(test_se), .CLK(CK), .Q(
        n8673), .QN(n4006) );
  SDFFX1 DFF_221_Q_reg ( .D(WX1835), .SI(n8673), .SE(test_se), .CLK(CK), .Q(
        n8672), .QN(n4005) );
  SDFFX1 DFF_222_Q_reg ( .D(WX1837), .SI(n8672), .SE(test_se), .CLK(CK), .Q(
        n8671), .QN(n4004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(test_se), .CLK(CK), .Q(
        n8670), .QN(n4003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(test_se), .CLK(CK), .Q(
        n8669), .QN(n3345) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(test_se), .CLK(CK), .Q(
        n8668), .QN(n3465) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(test_se), .CLK(CK), .Q(
        n8667), .QN(n3464) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(test_se), .CLK(CK), .Q(
        n8666), .QN(n3463) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(test_se), .CLK(CK), .Q(
        n8665), .QN(n3462) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(test_se), .CLK(CK), .Q(
        n8664), .QN(n3461) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(test_se), .CLK(CK), .Q(
        n8663), .QN(n3460) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(test_se), .CLK(CK), .Q(
        n8662), .QN(n3459) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(test_se), .CLK(CK), .Q(
        n8661), .QN(n3458) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(test_se), .CLK(CK), .Q(
        test_so13), .QN(n3457) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(test_se), .CLK(CK), 
        .Q(n8658), .QN(n3456) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(test_se), .CLK(CK), .Q(
        n8657), .QN(n3455) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(test_se), .CLK(CK), .Q(
        n8656), .QN(n3454) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(test_se), .CLK(CK), .Q(
        n8655), .QN(n3453) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(test_se), .CLK(CK), .Q(
        n8654), .QN(n3452) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(test_se), .CLK(CK), .Q(
        n8653), .QN(n3451) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(test_se), .CLK(CK), .Q(
        WX1970), .QN() );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(test_se), .CLK(CK), .Q(
        WX1972), .QN() );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(test_se), .CLK(CK), .Q(
        WX1974), .QN() );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(test_se), .CLK(CK), .Q(
        WX1976), .QN() );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(test_se), .CLK(CK), .Q(
        WX1978), .QN() );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(test_se), .CLK(CK), .Q(
        WX1980), .QN() );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(test_se), .CLK(CK), .Q(
        WX1982), .QN() );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(test_se), .CLK(CK), .Q(
        WX1984), .QN() );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(test_se), .CLK(CK), .Q(
        WX1986), .QN() );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(test_se), .CLK(CK), .Q(
        WX1988), .QN() );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(test_se), .CLK(CK), .Q(
        WX1990), .QN() );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(test_se), .CLK(CK), .Q(
        test_so14), .QN() );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(test_se), .CLK(CK), 
        .Q(WX1994), .QN() );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(test_se), .CLK(CK), .Q(
        WX1996), .QN() );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(test_se), .CLK(CK), .Q(
        WX1998), .QN() );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(test_se), .CLK(CK), .Q(
        WX2000), .QN() );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(test_se), .CLK(CK), .Q(
        WX2002), .QN() );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(test_se), .CLK(CK), .Q(
        WX2004), .QN() );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(test_se), .CLK(CK), .Q(
        WX2006), .QN() );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(test_se), .CLK(CK), .Q(
        WX2008), .QN() );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(test_se), .CLK(CK), .Q(
        WX2010), .QN() );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(test_se), .CLK(CK), .Q(
        WX2012), .QN() );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(test_se), .CLK(CK), .Q(
        WX2014), .QN() );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(test_se), .CLK(CK), .Q(
        WX2016), .QN() );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(test_se), .CLK(CK), .Q(
        WX2018), .QN() );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(test_se), .CLK(CK), .Q(
        WX2020), .QN() );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(test_se), .CLK(CK), .Q(
        WX2022), .QN() );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(test_se), .CLK(CK), .Q(
        WX2024), .QN() );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(test_se), .CLK(CK), .Q(
        WX2026), .QN() );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(test_se), .CLK(CK), .Q(
        test_so15), .QN() );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(test_se), .CLK(CK), 
        .Q(WX2030), .QN() );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(test_se), .CLK(CK), .Q(
        WX2032), .QN() );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(test_se), .CLK(CK), .Q(
        WX2034), .QN(n3785) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(test_se), .CLK(CK), .Q(
        WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(test_se), .CLK(CK), .Q(
        WX2038), .QN(n3781) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(test_se), .CLK(CK), .Q(
        WX2040), .QN(n3779) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(test_se), .CLK(CK), .Q(
        WX2042), .QN(n3777) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(test_se), .CLK(CK), .Q(
        WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(test_se), .CLK(CK), .Q(
        WX2046), .QN(n3773) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(test_se), .CLK(CK), .Q(
        WX2048), .QN(n3771) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(test_se), .CLK(CK), .Q(
        WX2050), .QN(n3769) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(test_se), .CLK(CK), .Q(
        WX2052), .QN(n3767) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(test_se), .CLK(CK), .Q(
        WX2054), .QN(n3765) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(test_se), .CLK(CK), .Q(
        WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(test_se), .CLK(CK), .Q(
        WX2058), .QN(n3761) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(test_se), .CLK(CK), .Q(
        WX2060), .QN(n3759) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(test_se), .CLK(CK), .Q(
        WX2062), .QN(n3757) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(test_se), .CLK(CK), .Q(
        test_so16), .QN(n3755) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(test_se), .CLK(CK), 
        .Q(WX2066), .QN() );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(test_se), .CLK(CK), .Q(
        WX2068), .QN() );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(test_se), .CLK(CK), .Q(
        WX2070), .QN() );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(test_se), .CLK(CK), .Q(
        WX2072), .QN() );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(test_se), .CLK(CK), .Q(
        WX2074), .QN() );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(test_se), .CLK(CK), .Q(
        WX2076), .QN() );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(test_se), .CLK(CK), .Q(
        WX2078), .QN() );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(test_se), .CLK(CK), .Q(
        WX2080), .QN() );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(test_se), .CLK(CK), .Q(
        WX2082), .QN() );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(test_se), .CLK(CK), .Q(
        WX2084), .QN() );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(test_se), .CLK(CK), .Q(
        WX2086), .QN() );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(test_se), .CLK(CK), .Q(
        WX2088), .QN() );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(test_se), .CLK(CK), .Q(
        WX2090), .QN() );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(test_se), .CLK(CK), .Q(
        WX2092), .QN() );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(test_se), .CLK(CK), .Q(
        WX2094), .QN() );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(test_se), .CLK(CK), .Q(
        WX2096), .QN() );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(test_se), .CLK(CK), .Q(
        WX2098), .QN() );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(test_se), .CLK(CK), .Q(
        test_so17), .QN() );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(test_se), .CLK(CK), 
        .Q(WX2102), .QN() );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(test_se), .CLK(CK), .Q(
        WX2104), .QN() );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(test_se), .CLK(CK), .Q(
        WX2106), .QN() );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(test_se), .CLK(CK), .Q(
        WX2108), .QN() );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(test_se), .CLK(CK), .Q(
        WX2110), .QN() );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(test_se), .CLK(CK), .Q(
        WX2112), .QN() );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(test_se), .CLK(CK), .Q(
        WX2114), .QN() );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(test_se), .CLK(CK), .Q(
        WX2116), .QN() );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(test_se), .CLK(CK), .Q(
        WX2118), .QN() );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(test_se), .CLK(CK), .Q(
        WX2120), .QN() );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(test_se), .CLK(CK), .Q(
        WX2122), .QN() );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(test_se), .CLK(CK), .Q(
        WX2124), .QN() );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(test_se), .CLK(CK), .Q(
        WX2126), .QN() );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(test_se), .CLK(CK), .Q(
        WX2128), .QN() );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(test_se), .CLK(CK), .Q(
        WX2130), .QN() );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(test_se), .CLK(CK), .Q(
        WX2132), .QN() );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(test_se), .CLK(CK), .Q(
        WX2134), .QN() );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(test_se), .CLK(CK), .Q(
        test_so18), .QN() );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(test_se), .CLK(CK), 
        .Q(WX2138), .QN() );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(test_se), .CLK(CK), .Q(
        WX2140), .QN() );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(test_se), .CLK(CK), .Q(
        WX2142), .QN() );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(test_se), .CLK(CK), .Q(
        WX2144), .QN() );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(test_se), .CLK(CK), .Q(
        WX2146), .QN() );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(test_se), .CLK(CK), .Q(
        WX2148), .QN() );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(test_se), .CLK(CK), .Q(
        WX2150), .QN() );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(test_se), .CLK(CK), .Q(
        WX2152), .QN() );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(test_se), .CLK(CK), .Q(
        WX2154), .QN() );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(test_se), .CLK(CK), .Q(
        WX2156), .QN() );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(test_se), .CLK(CK), .Q(
        WX2158), .QN() );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(test_se), .CLK(CK), .Q(
        WX2160), .QN() );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(test_se), .CLK(CK), .Q(
        WX2162), .QN() );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(test_se), .CLK(CK), .Q(
        WX2164), .QN() );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(test_se), .CLK(CK), .Q(
        WX2166), .QN() );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(test_se), .CLK(CK), .Q(
        WX2168), .QN() );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(test_se), .CLK(CK), .Q(
        WX2170), .QN() );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(test_se), .CLK(CK), .Q(
        test_so19), .QN() );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(test_se), .CLK(CK), 
        .Q(WX2174), .QN() );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(test_se), .CLK(CK), .Q(
        WX2176), .QN() );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(test_se), .CLK(CK), .Q(
        WX2178), .QN() );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(test_se), .CLK(CK), .Q(
        WX2180), .QN() );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(test_se), .CLK(CK), .Q(
        WX2182), .QN() );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(test_se), .CLK(CK), .Q(
        WX2184), .QN() );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(test_se), .CLK(CK), .Q(
        WX2186), .QN() );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(test_se), .CLK(CK), .Q(
        WX2188), .QN() );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(test_se), .CLK(CK), .Q(
        WX2190), .QN() );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(test_se), .CLK(CK), .Q(
        WX2192), .QN() );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_7), .QN(DFF_359_n1) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_25), .QN(DFF_377_n1) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(WX3070), .SI(CRC_OUT_8_31), .SE(test_se), .CLK(CK), 
        .Q(WX3071), .QN() );
  SDFFX1 DFF_385_Q_reg ( .D(WX3072), .SI(WX3071), .SE(test_se), .CLK(CK), .Q(
        n8644), .QN(n4002) );
  SDFFX1 DFF_386_Q_reg ( .D(WX3074), .SI(n8644), .SE(test_se), .CLK(CK), .Q(
        n8643), .QN(n4001) );
  SDFFX1 DFF_387_Q_reg ( .D(WX3076), .SI(n8643), .SE(test_se), .CLK(CK), .Q(
        n8642), .QN(n4000) );
  SDFFX1 DFF_388_Q_reg ( .D(WX3078), .SI(n8642), .SE(test_se), .CLK(CK), .Q(
        n8641), .QN(n3999) );
  SDFFX1 DFF_389_Q_reg ( .D(WX3080), .SI(n8641), .SE(test_se), .CLK(CK), .Q(
        n8640), .QN(n3998) );
  SDFFX1 DFF_390_Q_reg ( .D(WX3082), .SI(n8640), .SE(test_se), .CLK(CK), .Q(
        n8639), .QN(n3997) );
  SDFFX1 DFF_391_Q_reg ( .D(WX3084), .SI(n8639), .SE(test_se), .CLK(CK), .Q(
        n8638), .QN(n3996) );
  SDFFX1 DFF_392_Q_reg ( .D(WX3086), .SI(n8638), .SE(test_se), .CLK(CK), .Q(
        n8637), .QN(n3995) );
  SDFFX1 DFF_393_Q_reg ( .D(WX3088), .SI(n8637), .SE(test_se), .CLK(CK), .Q(
        n8636), .QN(n3994) );
  SDFFX1 DFF_394_Q_reg ( .D(WX3090), .SI(n8636), .SE(test_se), .CLK(CK), .Q(
        n8635), .QN(n3993) );
  SDFFX1 DFF_395_Q_reg ( .D(WX3092), .SI(n8635), .SE(test_se), .CLK(CK), .Q(
        test_so22), .QN(n3992) );
  SDFFX1 DFF_396_Q_reg ( .D(WX3094), .SI(test_si23), .SE(test_se), .CLK(CK), 
        .Q(n8632), .QN(n3991) );
  SDFFX1 DFF_397_Q_reg ( .D(WX3096), .SI(n8632), .SE(test_se), .CLK(CK), .Q(
        n8631), .QN(n3990) );
  SDFFX1 DFF_398_Q_reg ( .D(WX3098), .SI(n8631), .SE(test_se), .CLK(CK), .Q(
        n8630), .QN(n3989) );
  SDFFX1 DFF_399_Q_reg ( .D(WX3100), .SI(n8630), .SE(test_se), .CLK(CK), .Q(
        n8629), .QN(n3988) );
  SDFFX1 DFF_400_Q_reg ( .D(WX3102), .SI(n8629), .SE(test_se), .CLK(CK), .Q(
        n8628), .QN(n3987) );
  SDFFX1 DFF_401_Q_reg ( .D(WX3104), .SI(n8628), .SE(test_se), .CLK(CK), .Q(
        n8627), .QN(n3986) );
  SDFFX1 DFF_402_Q_reg ( .D(WX3106), .SI(n8627), .SE(test_se), .CLK(CK), .Q(
        n8626), .QN(n3985) );
  SDFFX1 DFF_403_Q_reg ( .D(WX3108), .SI(n8626), .SE(test_se), .CLK(CK), .Q(
        n8625), .QN(n3984) );
  SDFFX1 DFF_404_Q_reg ( .D(WX3110), .SI(n8625), .SE(test_se), .CLK(CK), .Q(
        n8624), .QN(n3983) );
  SDFFX1 DFF_405_Q_reg ( .D(WX3112), .SI(n8624), .SE(test_se), .CLK(CK), .Q(
        n8623), .QN(n3982) );
  SDFFX1 DFF_406_Q_reg ( .D(WX3114), .SI(n8623), .SE(test_se), .CLK(CK), .Q(
        n8622), .QN(n3981) );
  SDFFX1 DFF_407_Q_reg ( .D(WX3116), .SI(n8622), .SE(test_se), .CLK(CK), .Q(
        n8621), .QN(n3980) );
  SDFFX1 DFF_408_Q_reg ( .D(WX3118), .SI(n8621), .SE(test_se), .CLK(CK), .Q(
        n8620), .QN(n3979) );
  SDFFX1 DFF_409_Q_reg ( .D(WX3120), .SI(n8620), .SE(test_se), .CLK(CK), .Q(
        n8619), .QN(n3978) );
  SDFFX1 DFF_410_Q_reg ( .D(WX3122), .SI(n8619), .SE(test_se), .CLK(CK), .Q(
        n8618), .QN(n3977) );
  SDFFX1 DFF_411_Q_reg ( .D(WX3124), .SI(n8618), .SE(test_se), .CLK(CK), .Q(
        n8617), .QN(n3976) );
  SDFFX1 DFF_412_Q_reg ( .D(WX3126), .SI(n8617), .SE(test_se), .CLK(CK), .Q(
        n8616), .QN(n3975) );
  SDFFX1 DFF_413_Q_reg ( .D(WX3128), .SI(n8616), .SE(test_se), .CLK(CK), .Q(
        test_so23), .QN(n3974) );
  SDFFX1 DFF_414_Q_reg ( .D(WX3130), .SI(test_si24), .SE(test_se), .CLK(CK), 
        .Q(n8613), .QN(n3973) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(test_se), .CLK(CK), .Q(
        n8612), .QN(n3972) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(test_se), .CLK(CK), .Q(
        n8611), .QN(n3344) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(test_se), .CLK(CK), .Q(
        n8610), .QN(n3450) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(test_se), .CLK(CK), .Q(
        n8609), .QN(n3449) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(test_se), .CLK(CK), .Q(
        n8608), .QN(n3448) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(test_se), .CLK(CK), .Q(
        n8607), .QN(n3447) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(test_se), .CLK(CK), .Q(
        n8606), .QN(n3446) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(test_se), .CLK(CK), .Q(
        n8605), .QN(n3445) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(test_se), .CLK(CK), .Q(
        n8604), .QN(n3444) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(test_se), .CLK(CK), .Q(
        n8603), .QN(n3443) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(test_se), .CLK(CK), .Q(
        n8602), .QN(n3442) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(test_se), .CLK(CK), .Q(
        n8601), .QN(n3441) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(test_se), .CLK(CK), .Q(
        n8600), .QN(n3440) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(test_se), .CLK(CK), .Q(
        n8599), .QN(n3439) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(test_se), .CLK(CK), .Q(
        n8598), .QN(n3438) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(test_se), .CLK(CK), .Q(
        n8597), .QN(n3437) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(test_se), .CLK(CK), .Q(
        test_so24), .QN(n3436) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(test_se), .CLK(CK), 
        .Q(WX3263), .QN() );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(test_se), .CLK(CK), .Q(
        WX3265), .QN() );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(test_se), .CLK(CK), .Q(
        WX3267), .QN() );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(test_se), .CLK(CK), .Q(
        WX3269), .QN() );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(test_se), .CLK(CK), .Q(
        WX3271), .QN() );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(test_se), .CLK(CK), .Q(
        WX3273), .QN() );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(test_se), .CLK(CK), .Q(
        WX3275), .QN() );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(test_se), .CLK(CK), .Q(
        WX3277), .QN() );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(test_se), .CLK(CK), .Q(
        WX3279), .QN() );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(test_se), .CLK(CK), .Q(
        WX3281), .QN() );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(test_se), .CLK(CK), .Q(
        WX3283), .QN() );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(test_se), .CLK(CK), .Q(
        WX3285), .QN() );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(test_se), .CLK(CK), .Q(
        WX3287), .QN() );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(test_se), .CLK(CK), .Q(
        WX3289), .QN() );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(test_se), .CLK(CK), .Q(
        WX3291), .QN() );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(test_se), .CLK(CK), .Q(
        WX3293), .QN() );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(test_se), .CLK(CK), .Q(
        WX3295), .QN() );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(test_se), .CLK(CK), .Q(
        test_so25), .QN() );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(test_se), .CLK(CK), 
        .Q(WX3299), .QN() );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(test_se), .CLK(CK), .Q(
        WX3301), .QN() );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(test_se), .CLK(CK), .Q(
        WX3303), .QN() );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(test_se), .CLK(CK), .Q(
        WX3305), .QN() );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(test_se), .CLK(CK), .Q(
        WX3307), .QN() );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(test_se), .CLK(CK), .Q(
        WX3309), .QN() );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(test_se), .CLK(CK), .Q(
        WX3311), .QN() );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(test_se), .CLK(CK), .Q(
        WX3313), .QN() );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(test_se), .CLK(CK), .Q(
        WX3315), .QN() );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(test_se), .CLK(CK), .Q(
        WX3317), .QN() );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(test_se), .CLK(CK), .Q(
        WX3319), .QN() );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(test_se), .CLK(CK), .Q(
        WX3321), .QN() );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(test_se), .CLK(CK), .Q(
        WX3323), .QN() );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(test_se), .CLK(CK), .Q(
        WX3325), .QN() );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(test_se), .CLK(CK), .Q(
        WX3327), .QN(n3753) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(test_se), .CLK(CK), .Q(
        WX3329), .QN(n3751) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(test_se), .CLK(CK), .Q(
        WX3331), .QN(n3749) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(test_se), .CLK(CK), .Q(
        test_so26), .QN(n3747) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(test_se), .CLK(CK), 
        .Q(WX3335), .QN(n3745) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(test_se), .CLK(CK), .Q(
        WX3337), .QN(n3743) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(test_se), .CLK(CK), .Q(
        WX3339), .QN(n3741) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(test_se), .CLK(CK), .Q(
        WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(test_se), .CLK(CK), .Q(
        WX3343), .QN(n3737) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(test_se), .CLK(CK), .Q(
        WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(test_se), .CLK(CK), .Q(
        WX3347), .QN(n3733) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(test_se), .CLK(CK), .Q(
        WX3349), .QN(n3731) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(test_se), .CLK(CK), .Q(
        WX3351), .QN(n3729) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(test_se), .CLK(CK), .Q(
        WX3353), .QN(n3727) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(test_se), .CLK(CK), .Q(
        WX3355), .QN(n3725) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(test_se), .CLK(CK), .Q(
        WX3357), .QN(n3723) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(test_se), .CLK(CK), .Q(
        WX3359), .QN() );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(test_se), .CLK(CK), .Q(
        WX3361), .QN() );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(test_se), .CLK(CK), .Q(
        WX3363), .QN() );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(test_se), .CLK(CK), .Q(
        WX3365), .QN() );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(test_se), .CLK(CK), .Q(
        WX3367), .QN() );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(test_se), .CLK(CK), .Q(
        test_so27), .QN() );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(test_se), .CLK(CK), 
        .Q(WX3371), .QN() );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(test_se), .CLK(CK), .Q(
        WX3373), .QN() );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(test_se), .CLK(CK), .Q(
        WX3375), .QN() );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(test_se), .CLK(CK), .Q(
        WX3377), .QN() );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(test_se), .CLK(CK), .Q(
        WX3379), .QN() );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(test_se), .CLK(CK), .Q(
        WX3381), .QN() );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(test_se), .CLK(CK), .Q(
        WX3383), .QN() );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(test_se), .CLK(CK), .Q(
        WX3385), .QN() );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(test_se), .CLK(CK), .Q(
        WX3387), .QN() );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(test_se), .CLK(CK), .Q(
        WX3389), .QN() );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(test_se), .CLK(CK), .Q(
        WX3391), .QN() );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(test_se), .CLK(CK), .Q(
        WX3393), .QN() );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(test_se), .CLK(CK), .Q(
        WX3395), .QN() );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(test_se), .CLK(CK), .Q(
        WX3397), .QN() );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(test_se), .CLK(CK), .Q(
        WX3399), .QN() );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(test_se), .CLK(CK), .Q(
        WX3401), .QN() );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(test_se), .CLK(CK), .Q(
        WX3403), .QN() );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(test_se), .CLK(CK), .Q(
        test_so28), .QN() );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(test_se), .CLK(CK), 
        .Q(WX3407), .QN() );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(test_se), .CLK(CK), .Q(
        WX3409), .QN() );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(test_se), .CLK(CK), .Q(
        WX3411), .QN() );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(test_se), .CLK(CK), .Q(
        WX3413), .QN() );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(test_se), .CLK(CK), .Q(
        WX3415), .QN() );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(test_se), .CLK(CK), .Q(
        WX3417), .QN() );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(test_se), .CLK(CK), .Q(
        WX3419), .QN() );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(test_se), .CLK(CK), .Q(
        WX3421), .QN() );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(test_se), .CLK(CK), .Q(
        WX3423), .QN() );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(test_se), .CLK(CK), .Q(
        WX3425), .QN() );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(test_se), .CLK(CK), .Q(
        WX3427), .QN() );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(test_se), .CLK(CK), .Q(
        WX3429), .QN() );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(test_se), .CLK(CK), .Q(
        WX3431), .QN() );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(test_se), .CLK(CK), .Q(
        WX3433), .QN() );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(test_se), .CLK(CK), .Q(
        WX3435), .QN() );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(test_se), .CLK(CK), .Q(
        WX3437), .QN() );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(test_se), .CLK(CK), .Q(
        test_so29), .QN() );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(test_se), .CLK(CK), 
        .Q(WX3441), .QN() );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(test_se), .CLK(CK), .Q(
        WX3443), .QN() );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(test_se), .CLK(CK), .Q(
        WX3445), .QN() );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(test_se), .CLK(CK), .Q(
        WX3447), .QN() );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(test_se), .CLK(CK), .Q(
        WX3449), .QN() );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(test_se), .CLK(CK), .Q(
        WX3451), .QN() );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(test_se), .CLK(CK), .Q(
        WX3453), .QN() );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(test_se), .CLK(CK), .Q(
        WX3455), .QN() );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(test_se), .CLK(CK), .Q(
        WX3457), .QN() );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(test_se), .CLK(CK), .Q(
        WX3459), .QN() );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(test_se), .CLK(CK), .Q(
        WX3461), .QN() );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(test_se), .CLK(CK), .Q(
        WX3463), .QN() );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(test_se), .CLK(CK), .Q(
        WX3465), .QN() );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(test_se), .CLK(CK), .Q(
        WX3467), .QN() );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(test_se), .CLK(CK), .Q(
        WX3469), .QN() );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(test_se), .CLK(CK), .Q(
        WX3471), .QN() );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(test_se), .CLK(CK), .Q(
        test_so30), .QN() );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(test_se), .CLK(CK), 
        .Q(WX3475), .QN() );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(test_se), .CLK(CK), .Q(
        WX3477), .QN() );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(test_se), .CLK(CK), .Q(
        WX3479), .QN() );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(test_se), .CLK(CK), .Q(
        WX3481), .QN() );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(test_se), .CLK(CK), .Q(
        WX3483), .QN() );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(test_se), .CLK(CK), .Q(
        WX3485), .QN() );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_10), .QN(DFF_554_n1) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_27), .QN(DFF_571_n1) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(WX4363), .SI(CRC_OUT_7_31), .SE(test_se), .CLK(CK), 
        .Q(WX4364), .QN() );
  SDFFX1 DFF_577_Q_reg ( .D(WX4365), .SI(WX4364), .SE(test_se), .CLK(CK), .Q(
        n8586), .QN(n3971) );
  SDFFX1 DFF_578_Q_reg ( .D(WX4367), .SI(n8586), .SE(test_se), .CLK(CK), .Q(
        n8585), .QN(n3970) );
  SDFFX1 DFF_579_Q_reg ( .D(WX4369), .SI(n8585), .SE(test_se), .CLK(CK), .Q(
        n8584), .QN(n3969) );
  SDFFX1 DFF_580_Q_reg ( .D(WX4371), .SI(n8584), .SE(test_se), .CLK(CK), .Q(
        n8583), .QN(n3968) );
  SDFFX1 DFF_581_Q_reg ( .D(WX4373), .SI(n8583), .SE(test_se), .CLK(CK), .Q(
        n8582), .QN(n3967) );
  SDFFX1 DFF_582_Q_reg ( .D(WX4375), .SI(n8582), .SE(test_se), .CLK(CK), .Q(
        n8581), .QN(n3966) );
  SDFFX1 DFF_583_Q_reg ( .D(WX4377), .SI(n8581), .SE(test_se), .CLK(CK), .Q(
        n8580), .QN(n3965) );
  SDFFX1 DFF_584_Q_reg ( .D(WX4379), .SI(n8580), .SE(test_se), .CLK(CK), .Q(
        n8579), .QN(n3964) );
  SDFFX1 DFF_585_Q_reg ( .D(WX4381), .SI(n8579), .SE(test_se), .CLK(CK), .Q(
        n8578), .QN(n3963) );
  SDFFX1 DFF_586_Q_reg ( .D(WX4383), .SI(n8578), .SE(test_se), .CLK(CK), .Q(
        n8577), .QN(n3962) );
  SDFFX1 DFF_587_Q_reg ( .D(WX4385), .SI(n8577), .SE(test_se), .CLK(CK), .Q(
        n8576), .QN(n3961) );
  SDFFX1 DFF_588_Q_reg ( .D(WX4387), .SI(n8576), .SE(test_se), .CLK(CK), .Q(
        test_so33), .QN(n3960) );
  SDFFX1 DFF_589_Q_reg ( .D(WX4389), .SI(test_si34), .SE(test_se), .CLK(CK), 
        .Q(n8573), .QN(n3959) );
  SDFFX1 DFF_590_Q_reg ( .D(WX4391), .SI(n8573), .SE(test_se), .CLK(CK), .Q(
        n8572), .QN(n3958) );
  SDFFX1 DFF_591_Q_reg ( .D(WX4393), .SI(n8572), .SE(test_se), .CLK(CK), .Q(
        n8571), .QN(n3957) );
  SDFFX1 DFF_592_Q_reg ( .D(WX4395), .SI(n8571), .SE(test_se), .CLK(CK), .Q(
        n8570), .QN(n3956) );
  SDFFX1 DFF_593_Q_reg ( .D(WX4397), .SI(n8570), .SE(test_se), .CLK(CK), .Q(
        n8569), .QN(n3955) );
  SDFFX1 DFF_594_Q_reg ( .D(WX4399), .SI(n8569), .SE(test_se), .CLK(CK), .Q(
        n8568), .QN(n3954) );
  SDFFX1 DFF_595_Q_reg ( .D(WX4401), .SI(n8568), .SE(test_se), .CLK(CK), .Q(
        n8567), .QN(n3953) );
  SDFFX1 DFF_596_Q_reg ( .D(WX4403), .SI(n8567), .SE(test_se), .CLK(CK), .Q(
        n8566), .QN(n3952) );
  SDFFX1 DFF_597_Q_reg ( .D(WX4405), .SI(n8566), .SE(test_se), .CLK(CK), .Q(
        n8565), .QN(n3951) );
  SDFFX1 DFF_598_Q_reg ( .D(WX4407), .SI(n8565), .SE(test_se), .CLK(CK), .Q(
        n8564), .QN(n3950) );
  SDFFX1 DFF_599_Q_reg ( .D(WX4409), .SI(n8564), .SE(test_se), .CLK(CK), .Q(
        n8563), .QN(n3949) );
  SDFFX1 DFF_600_Q_reg ( .D(WX4411), .SI(n8563), .SE(test_se), .CLK(CK), .Q(
        n8562), .QN(n3948) );
  SDFFX1 DFF_601_Q_reg ( .D(WX4413), .SI(n8562), .SE(test_se), .CLK(CK), .Q(
        n8561), .QN(n3947) );
  SDFFX1 DFF_602_Q_reg ( .D(WX4415), .SI(n8561), .SE(test_se), .CLK(CK), .Q(
        n8560), .QN(n3946) );
  SDFFX1 DFF_603_Q_reg ( .D(WX4417), .SI(n8560), .SE(test_se), .CLK(CK), .Q(
        n8559), .QN(n3945) );
  SDFFX1 DFF_604_Q_reg ( .D(WX4419), .SI(n8559), .SE(test_se), .CLK(CK), .Q(
        n8558), .QN(n3944) );
  SDFFX1 DFF_605_Q_reg ( .D(WX4421), .SI(n8558), .SE(test_se), .CLK(CK), .Q(
        test_so34), .QN(n3943) );
  SDFFX1 DFF_606_Q_reg ( .D(WX4423), .SI(test_si35), .SE(test_se), .CLK(CK), 
        .Q(n8555), .QN(n3942) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(test_se), .CLK(CK), .Q(
        n8554), .QN(n3941) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(test_se), .CLK(CK), .Q(
        n8553), .QN(n3343) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(test_se), .CLK(CK), .Q(
        n8552), .QN(n3435) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(test_se), .CLK(CK), .Q(
        n8551), .QN(n3434) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(test_se), .CLK(CK), .Q(
        n8550), .QN(n3433) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(test_se), .CLK(CK), .Q(
        n8549), .QN(n3432) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(test_se), .CLK(CK), .Q(
        n8548), .QN(n3431) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(test_se), .CLK(CK), .Q(
        n8547), .QN(n3430) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(test_se), .CLK(CK), .Q(
        n8546), .QN(n3429) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(test_se), .CLK(CK), .Q(
        n8545), .QN(n3428) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(test_se), .CLK(CK), .Q(
        n8544), .QN(n3427) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(test_se), .CLK(CK), .Q(
        n8543), .QN(n3426) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(test_se), .CLK(CK), .Q(
        n8542), .QN(n3425) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(test_se), .CLK(CK), .Q(
        n8541), .QN(n3424) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(test_se), .CLK(CK), .Q(
        n8540), .QN(n3423) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(test_se), .CLK(CK), .Q(
        test_so35), .QN(n3422) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(test_se), .CLK(CK), 
        .Q(n8537), .QN(n3421) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(test_se), .CLK(CK), .Q(
        WX4556), .QN() );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(test_se), .CLK(CK), .Q(
        WX4558), .QN() );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(test_se), .CLK(CK), .Q(
        WX4560), .QN() );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(test_se), .CLK(CK), .Q(
        WX4562), .QN() );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(test_se), .CLK(CK), .Q(
        WX4564), .QN() );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(test_se), .CLK(CK), .Q(
        WX4566), .QN() );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(test_se), .CLK(CK), .Q(
        WX4568), .QN() );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(test_se), .CLK(CK), .Q(
        WX4570), .QN() );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(test_se), .CLK(CK), .Q(
        WX4572), .QN() );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(test_se), .CLK(CK), .Q(
        WX4574), .QN() );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(test_se), .CLK(CK), .Q(
        WX4576), .QN() );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(test_se), .CLK(CK), .Q(
        WX4578), .QN() );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(test_se), .CLK(CK), .Q(
        WX4580), .QN() );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(test_se), .CLK(CK), .Q(
        WX4582), .QN() );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(test_se), .CLK(CK), .Q(
        WX4584), .QN() );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(test_se), .CLK(CK), .Q(
        test_so36), .QN() );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(test_se), .CLK(CK), 
        .Q(WX4588), .QN() );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(test_se), .CLK(CK), .Q(
        WX4590), .QN() );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(test_se), .CLK(CK), .Q(
        WX4592), .QN() );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(test_se), .CLK(CK), .Q(
        WX4594), .QN() );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(test_se), .CLK(CK), .Q(
        WX4596), .QN() );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(test_se), .CLK(CK), .Q(
        WX4598), .QN() );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(test_se), .CLK(CK), .Q(
        WX4600), .QN() );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(test_se), .CLK(CK), .Q(
        WX4602), .QN() );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(test_se), .CLK(CK), .Q(
        WX4604), .QN() );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(test_se), .CLK(CK), .Q(
        WX4606), .QN() );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(test_se), .CLK(CK), .Q(
        WX4608), .QN() );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(test_se), .CLK(CK), .Q(
        WX4610), .QN() );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(test_se), .CLK(CK), .Q(
        WX4612), .QN() );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(test_se), .CLK(CK), .Q(
        WX4614), .QN() );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(test_se), .CLK(CK), .Q(
        WX4616), .QN() );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(test_se), .CLK(CK), .Q(
        WX4618), .QN() );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(test_se), .CLK(CK), .Q(
        test_so37), .QN(n3721) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(test_se), .CLK(CK), 
        .Q(WX4622), .QN(n3719) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(test_se), .CLK(CK), .Q(
        WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(test_se), .CLK(CK), .Q(
        WX4626), .QN(n3715) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(test_se), .CLK(CK), .Q(
        WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(test_se), .CLK(CK), .Q(
        WX4630), .QN(n3711) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(test_se), .CLK(CK), .Q(
        WX4632), .QN(n3709) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(test_se), .CLK(CK), .Q(
        WX4634), .QN(n3707) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(test_se), .CLK(CK), .Q(
        WX4636), .QN(n3705) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(test_se), .CLK(CK), .Q(
        WX4638), .QN(n3703) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(test_se), .CLK(CK), .Q(
        WX4640), .QN(n3701) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(test_se), .CLK(CK), .Q(
        WX4642), .QN(n3699) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(test_se), .CLK(CK), .Q(
        WX4644), .QN(n3697) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(test_se), .CLK(CK), .Q(
        WX4646), .QN(n3695) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(test_se), .CLK(CK), .Q(
        WX4648), .QN(n3693) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(test_se), .CLK(CK), .Q(
        WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(test_se), .CLK(CK), .Q(
        WX4652), .QN() );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(test_se), .CLK(CK), .Q(
        test_so38), .QN() );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(test_se), .CLK(CK), 
        .Q(WX4656), .QN() );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(test_se), .CLK(CK), .Q(
        WX4658), .QN() );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(test_se), .CLK(CK), .Q(
        WX4660), .QN() );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(test_se), .CLK(CK), .Q(
        WX4662), .QN() );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(test_se), .CLK(CK), .Q(
        WX4664), .QN() );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(test_se), .CLK(CK), .Q(
        WX4666), .QN() );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(test_se), .CLK(CK), .Q(
        WX4668), .QN() );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(test_se), .CLK(CK), .Q(
        WX4670), .QN() );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(test_se), .CLK(CK), .Q(
        WX4672), .QN() );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(test_se), .CLK(CK), .Q(
        WX4674), .QN() );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(test_se), .CLK(CK), .Q(
        WX4676), .QN() );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(test_se), .CLK(CK), .Q(
        WX4678), .QN() );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(test_se), .CLK(CK), .Q(
        WX4680), .QN() );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(test_se), .CLK(CK), .Q(
        WX4682), .QN() );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(test_se), .CLK(CK), .Q(
        WX4684), .QN() );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(test_se), .CLK(CK), .Q(
        WX4686), .QN() );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(test_se), .CLK(CK), .Q(
        test_so39), .QN() );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(test_se), .CLK(CK), 
        .Q(WX4690), .QN() );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(test_se), .CLK(CK), .Q(
        WX4692), .QN() );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(test_se), .CLK(CK), .Q(
        WX4694), .QN() );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(test_se), .CLK(CK), .Q(
        WX4696), .QN() );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(test_se), .CLK(CK), .Q(
        WX4698), .QN() );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(test_se), .CLK(CK), .Q(
        WX4700), .QN() );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(test_se), .CLK(CK), .Q(
        WX4702), .QN() );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(test_se), .CLK(CK), .Q(
        WX4704), .QN() );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(test_se), .CLK(CK), .Q(
        WX4706), .QN() );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(test_se), .CLK(CK), .Q(
        WX4708), .QN() );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(test_se), .CLK(CK), .Q(
        WX4710), .QN() );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(test_se), .CLK(CK), .Q(
        WX4712), .QN() );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(test_se), .CLK(CK), .Q(
        WX4714), .QN() );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(test_se), .CLK(CK), .Q(
        WX4716), .QN() );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(test_se), .CLK(CK), .Q(
        WX4718), .QN() );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(test_se), .CLK(CK), .Q(
        WX4720), .QN() );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(test_se), .CLK(CK), .Q(
        test_so40), .QN() );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(test_se), .CLK(CK), 
        .Q(WX4724), .QN() );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(test_se), .CLK(CK), .Q(
        WX4726), .QN() );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(test_se), .CLK(CK), .Q(
        WX4728), .QN() );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(test_se), .CLK(CK), .Q(
        WX4730), .QN() );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(test_se), .CLK(CK), .Q(
        WX4732), .QN() );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(test_se), .CLK(CK), .Q(
        WX4734), .QN() );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(test_se), .CLK(CK), .Q(
        WX4736), .QN() );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(test_se), .CLK(CK), .Q(
        WX4738), .QN() );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(test_se), .CLK(CK), .Q(
        WX4740), .QN() );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(test_se), .CLK(CK), .Q(
        WX4742), .QN() );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(test_se), .CLK(CK), .Q(
        WX4744), .QN() );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(test_se), .CLK(CK), .Q(
        WX4746), .QN() );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(test_se), .CLK(CK), .Q(
        WX4748), .QN() );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(test_se), .CLK(CK), .Q(
        WX4750), .QN() );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(test_se), .CLK(CK), .Q(
        WX4752), .QN() );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(test_se), .CLK(CK), .Q(
        WX4754), .QN() );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(test_se), .CLK(CK), .Q(
        test_so41), .QN() );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(test_se), .CLK(CK), 
        .Q(WX4758), .QN() );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(test_se), .CLK(CK), .Q(
        WX4760), .QN() );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(test_se), .CLK(CK), .Q(
        WX4762), .QN() );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(test_se), .CLK(CK), .Q(
        WX4764), .QN() );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(test_se), .CLK(CK), .Q(
        WX4766), .QN() );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(test_se), .CLK(CK), .Q(
        WX4768), .QN() );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(test_se), .CLK(CK), .Q(
        WX4770), .QN() );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(test_se), .CLK(CK), .Q(
        WX4772), .QN() );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(test_se), .CLK(CK), .Q(
        WX4774), .QN() );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(test_se), .CLK(CK), .Q(
        WX4776), .QN() );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(test_se), .CLK(CK), .Q(
        WX4778), .QN() );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_5), .QN(DFF_741_n1) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_22), .QN(DFF_758_n1) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(WX5656), .SI(CRC_OUT_6_31), .SE(test_se), .CLK(CK), 
        .Q(WX5657), .QN() );
  SDFFX1 DFF_769_Q_reg ( .D(WX5658), .SI(WX5657), .SE(test_se), .CLK(CK), .Q(
        n8528), .QN(n3940) );
  SDFFX1 DFF_770_Q_reg ( .D(WX5660), .SI(n8528), .SE(test_se), .CLK(CK), .Q(
        n8527), .QN(n3939) );
  SDFFX1 DFF_771_Q_reg ( .D(WX5662), .SI(n8527), .SE(test_se), .CLK(CK), .Q(
        n8526), .QN(n3938) );
  SDFFX1 DFF_772_Q_reg ( .D(WX5664), .SI(n8526), .SE(test_se), .CLK(CK), .Q(
        n8525), .QN(n3937) );
  SDFFX1 DFF_773_Q_reg ( .D(WX5666), .SI(n8525), .SE(test_se), .CLK(CK), .Q(
        n8524), .QN(n3936) );
  SDFFX1 DFF_774_Q_reg ( .D(WX5668), .SI(n8524), .SE(test_se), .CLK(CK), .Q(
        n8523), .QN(n3935) );
  SDFFX1 DFF_775_Q_reg ( .D(WX5670), .SI(n8523), .SE(test_se), .CLK(CK), .Q(
        test_so44), .QN(n3934) );
  SDFFX1 DFF_776_Q_reg ( .D(WX5672), .SI(test_si45), .SE(test_se), .CLK(CK), 
        .Q(n8520), .QN(n3933) );
  SDFFX1 DFF_777_Q_reg ( .D(WX5674), .SI(n8520), .SE(test_se), .CLK(CK), .Q(
        n8519), .QN(n3932) );
  SDFFX1 DFF_778_Q_reg ( .D(WX5676), .SI(n8519), .SE(test_se), .CLK(CK), .Q(
        n8518), .QN(n3931) );
  SDFFX1 DFF_779_Q_reg ( .D(WX5678), .SI(n8518), .SE(test_se), .CLK(CK), .Q(
        n8517), .QN(n3930) );
  SDFFX1 DFF_780_Q_reg ( .D(WX5680), .SI(n8517), .SE(test_se), .CLK(CK), .Q(
        n8516), .QN(n3929) );
  SDFFX1 DFF_781_Q_reg ( .D(WX5682), .SI(n8516), .SE(test_se), .CLK(CK), .Q(
        n8515), .QN(n3928) );
  SDFFX1 DFF_782_Q_reg ( .D(WX5684), .SI(n8515), .SE(test_se), .CLK(CK), .Q(
        n8514), .QN(n3927) );
  SDFFX1 DFF_783_Q_reg ( .D(WX5686), .SI(n8514), .SE(test_se), .CLK(CK), .Q(
        n8513), .QN(n3926) );
  SDFFX1 DFF_784_Q_reg ( .D(WX5688), .SI(n8513), .SE(test_se), .CLK(CK), .Q(
        n8512), .QN(n3925) );
  SDFFX1 DFF_785_Q_reg ( .D(WX5690), .SI(n8512), .SE(test_se), .CLK(CK), .Q(
        n8511), .QN(n3924) );
  SDFFX1 DFF_786_Q_reg ( .D(WX5692), .SI(n8511), .SE(test_se), .CLK(CK), .Q(
        n8510), .QN(n3923) );
  SDFFX1 DFF_787_Q_reg ( .D(WX5694), .SI(n8510), .SE(test_se), .CLK(CK), .Q(
        n8509), .QN(n3922) );
  SDFFX1 DFF_788_Q_reg ( .D(WX5696), .SI(n8509), .SE(test_se), .CLK(CK), .Q(
        n8508), .QN(n3921) );
  SDFFX1 DFF_789_Q_reg ( .D(WX5698), .SI(n8508), .SE(test_se), .CLK(CK), .Q(
        n8507), .QN(n3920) );
  SDFFX1 DFF_790_Q_reg ( .D(WX5700), .SI(n8507), .SE(test_se), .CLK(CK), .Q(
        n8506), .QN(n3919) );
  SDFFX1 DFF_791_Q_reg ( .D(WX5702), .SI(n8506), .SE(test_se), .CLK(CK), .Q(
        n8505), .QN(n3918) );
  SDFFX1 DFF_792_Q_reg ( .D(WX5704), .SI(n8505), .SE(test_se), .CLK(CK), .Q(
        test_so45), .QN(n3917) );
  SDFFX1 DFF_793_Q_reg ( .D(WX5706), .SI(test_si46), .SE(test_se), .CLK(CK), 
        .Q(n8502), .QN(n3916) );
  SDFFX1 DFF_794_Q_reg ( .D(WX5708), .SI(n8502), .SE(test_se), .CLK(CK), .Q(
        n8501), .QN(n3915) );
  SDFFX1 DFF_795_Q_reg ( .D(WX5710), .SI(n8501), .SE(test_se), .CLK(CK), .Q(
        n8500), .QN(n3914) );
  SDFFX1 DFF_796_Q_reg ( .D(WX5712), .SI(n8500), .SE(test_se), .CLK(CK), .Q(
        n8499), .QN(n3913) );
  SDFFX1 DFF_797_Q_reg ( .D(WX5714), .SI(n8499), .SE(test_se), .CLK(CK), .Q(
        n8498), .QN(n3912) );
  SDFFX1 DFF_798_Q_reg ( .D(WX5716), .SI(n8498), .SE(test_se), .CLK(CK), .Q(
        n8497), .QN(n3911) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(test_se), .CLK(CK), .Q(
        n8496), .QN(n3910) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(test_se), .CLK(CK), .Q(
        n8495), .QN(n3342) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(test_se), .CLK(CK), .Q(
        n8494), .QN(n3420) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(test_se), .CLK(CK), .Q(
        n8493), .QN(n3419) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(test_se), .CLK(CK), .Q(
        n8492), .QN(n3418) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(test_se), .CLK(CK), .Q(
        n8491), .QN(n3417) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(test_se), .CLK(CK), .Q(
        n8490), .QN(n3416) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(test_se), .CLK(CK), .Q(
        n8489), .QN(n3415) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(test_se), .CLK(CK), .Q(
        n8488), .QN(n3414) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(test_se), .CLK(CK), .Q(
        n8487), .QN(n3413) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(test_se), .CLK(CK), .Q(
        test_so46), .QN(n3412) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(test_se), .CLK(CK), 
        .Q(n8484), .QN(n3411) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(test_se), .CLK(CK), .Q(
        n8483), .QN(n3410) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(test_se), .CLK(CK), .Q(
        n8482), .QN(n3409) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(test_se), .CLK(CK), .Q(
        n8481), .QN(n3408) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(test_se), .CLK(CK), .Q(
        n8480), .QN(n3407) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(test_se), .CLK(CK), .Q(
        n8479), .QN(n3406) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(test_se), .CLK(CK), .Q(
        WX5849), .QN() );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(test_se), .CLK(CK), .Q(
        WX5851), .QN() );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(test_se), .CLK(CK), .Q(
        WX5853), .QN() );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(test_se), .CLK(CK), .Q(
        WX5855), .QN() );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(test_se), .CLK(CK), .Q(
        WX5857), .QN() );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(test_se), .CLK(CK), .Q(
        WX5859), .QN() );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(test_se), .CLK(CK), .Q(
        WX5861), .QN() );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(test_se), .CLK(CK), .Q(
        WX5863), .QN() );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(test_se), .CLK(CK), .Q(
        WX5865), .QN() );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(test_se), .CLK(CK), .Q(
        WX5867), .QN() );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(test_se), .CLK(CK), .Q(
        test_so47), .QN() );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(test_se), .CLK(CK), 
        .Q(WX5871), .QN() );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(test_se), .CLK(CK), .Q(
        WX5873), .QN() );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(test_se), .CLK(CK), .Q(
        WX5875), .QN() );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(test_se), .CLK(CK), .Q(
        WX5877), .QN() );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(test_se), .CLK(CK), .Q(
        WX5879), .QN() );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(test_se), .CLK(CK), .Q(
        WX5881), .QN() );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(test_se), .CLK(CK), .Q(
        WX5883), .QN() );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(test_se), .CLK(CK), .Q(
        WX5885), .QN() );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(test_se), .CLK(CK), .Q(
        WX5887), .QN() );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(test_se), .CLK(CK), .Q(
        WX5889), .QN() );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(test_se), .CLK(CK), .Q(
        WX5891), .QN() );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(test_se), .CLK(CK), .Q(
        WX5893), .QN() );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(test_se), .CLK(CK), .Q(
        WX5895), .QN() );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(test_se), .CLK(CK), .Q(
        WX5897), .QN() );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(test_se), .CLK(CK), .Q(
        WX5899), .QN() );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(test_se), .CLK(CK), .Q(
        WX5901), .QN() );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(test_se), .CLK(CK), .Q(
        test_so48), .QN() );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(test_se), .CLK(CK), 
        .Q(WX5905), .QN() );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(test_se), .CLK(CK), .Q(
        WX5907), .QN() );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(test_se), .CLK(CK), .Q(
        WX5909), .QN() );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(test_se), .CLK(CK), .Q(
        WX5911), .QN() );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(test_se), .CLK(CK), .Q(
        WX5913), .QN(n3689) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(test_se), .CLK(CK), .Q(
        WX5915), .QN(n3687) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(test_se), .CLK(CK), .Q(
        WX5917), .QN(n3685) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(test_se), .CLK(CK), .Q(
        WX5919), .QN(n3683) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(test_se), .CLK(CK), .Q(
        WX5921), .QN(n3681) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(test_se), .CLK(CK), .Q(
        WX5923), .QN(n3679) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(test_se), .CLK(CK), .Q(
        WX5925), .QN(n3677) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(test_se), .CLK(CK), .Q(
        WX5927), .QN(n3675) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(test_se), .CLK(CK), .Q(
        WX5929), .QN(n3673) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(test_se), .CLK(CK), .Q(
        WX5931), .QN(n3671) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(test_se), .CLK(CK), .Q(
        WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(test_se), .CLK(CK), .Q(
        WX5935), .QN(n3667) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(test_se), .CLK(CK), .Q(
        test_so49), .QN(n3665) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(test_se), .CLK(CK), 
        .Q(WX5939), .QN(n3663) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(test_se), .CLK(CK), .Q(
        WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(test_se), .CLK(CK), .Q(
        WX5943), .QN(n3659) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(test_se), .CLK(CK), .Q(
        WX5945), .QN() );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(test_se), .CLK(CK), .Q(
        WX5947), .QN() );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(test_se), .CLK(CK), .Q(
        WX5949), .QN() );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(test_se), .CLK(CK), .Q(
        WX5951), .QN() );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(test_se), .CLK(CK), .Q(
        WX5953), .QN() );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(test_se), .CLK(CK), .Q(
        WX5955), .QN() );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(test_se), .CLK(CK), .Q(
        WX5957), .QN() );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(test_se), .CLK(CK), .Q(
        WX5959), .QN() );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(test_se), .CLK(CK), .Q(
        WX5961), .QN() );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(test_se), .CLK(CK), .Q(
        WX5963), .QN() );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(test_se), .CLK(CK), .Q(
        WX5965), .QN() );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(test_se), .CLK(CK), .Q(
        WX5967), .QN() );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(test_se), .CLK(CK), .Q(
        WX5969), .QN() );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(test_se), .CLK(CK), .Q(
        test_so50), .QN() );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(test_se), .CLK(CK), 
        .Q(WX5973), .QN() );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(test_se), .CLK(CK), .Q(
        WX5975), .QN() );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(test_se), .CLK(CK), .Q(
        WX5977), .QN() );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(test_se), .CLK(CK), .Q(
        WX5979), .QN() );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(test_se), .CLK(CK), .Q(
        WX5981), .QN() );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(test_se), .CLK(CK), .Q(
        WX5983), .QN() );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(test_se), .CLK(CK), .Q(
        WX5985), .QN() );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(test_se), .CLK(CK), .Q(
        WX5987), .QN() );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(test_se), .CLK(CK), .Q(
        WX5989), .QN() );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(test_se), .CLK(CK), .Q(
        WX5991), .QN() );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(test_se), .CLK(CK), .Q(
        WX5993), .QN() );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(test_se), .CLK(CK), .Q(
        WX5995), .QN() );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(test_se), .CLK(CK), .Q(
        WX5997), .QN() );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(test_se), .CLK(CK), .Q(
        WX5999), .QN() );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(test_se), .CLK(CK), .Q(
        WX6001), .QN() );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(test_se), .CLK(CK), .Q(
        WX6003), .QN() );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(test_se), .CLK(CK), .Q(
        test_so51), .QN() );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(test_se), .CLK(CK), 
        .Q(WX6007), .QN() );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(test_se), .CLK(CK), .Q(
        WX6009), .QN() );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(test_se), .CLK(CK), .Q(
        WX6011), .QN() );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(test_se), .CLK(CK), .Q(
        WX6013), .QN() );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(test_se), .CLK(CK), .Q(
        WX6015), .QN() );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(test_se), .CLK(CK), .Q(
        WX6017), .QN() );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(test_se), .CLK(CK), .Q(
        WX6019), .QN() );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(test_se), .CLK(CK), .Q(
        WX6021), .QN() );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(test_se), .CLK(CK), .Q(
        WX6023), .QN() );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(test_se), .CLK(CK), .Q(
        WX6025), .QN() );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(test_se), .CLK(CK), .Q(
        WX6027), .QN() );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(test_se), .CLK(CK), .Q(
        WX6029), .QN() );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(test_se), .CLK(CK), .Q(
        WX6031), .QN() );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(test_se), .CLK(CK), .Q(
        WX6033), .QN() );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(test_se), .CLK(CK), .Q(
        WX6035), .QN() );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(test_se), .CLK(CK), .Q(
        WX6037), .QN() );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(test_se), .CLK(CK), .Q(
        test_so52), .QN() );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(test_se), .CLK(CK), 
        .Q(WX6041), .QN() );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(test_se), .CLK(CK), .Q(
        WX6043), .QN() );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(test_se), .CLK(CK), .Q(
        WX6045), .QN() );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(test_se), .CLK(CK), .Q(
        WX6047), .QN() );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(test_se), .CLK(CK), .Q(
        WX6049), .QN() );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(test_se), .CLK(CK), .Q(
        WX6051), .QN() );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(test_se), .CLK(CK), .Q(
        WX6053), .QN() );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(test_se), .CLK(CK), .Q(
        WX6055), .QN() );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(test_se), .CLK(CK), .Q(
        WX6057), .QN() );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(test_se), .CLK(CK), .Q(
        WX6059), .QN() );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(test_se), .CLK(CK), .Q(
        WX6061), .QN() );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(test_se), .CLK(CK), .Q(
        WX6063), .QN() );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(test_se), .CLK(CK), .Q(
        WX6065), .QN() );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(test_se), .CLK(CK), .Q(
        WX6067), .QN() );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(test_se), .CLK(CK), .Q(
        WX6069), .QN() );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(test_se), .CLK(CK), .Q(
        WX6071), .QN() );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_5_0), .QN(DFF_928_n1) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_17), .QN(DFF_945_n1) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(WX6949), .SI(CRC_OUT_5_31), .SE(test_se), .CLK(CK), 
        .Q(WX6950), .QN() );
  SDFFX1 DFF_961_Q_reg ( .D(WX6951), .SI(WX6950), .SE(test_se), .CLK(CK), .Q(
        n8470), .QN(n3909) );
  SDFFX1 DFF_962_Q_reg ( .D(WX6953), .SI(n8470), .SE(test_se), .CLK(CK), .Q(
        test_so55), .QN(n3908) );
  SDFFX1 DFF_963_Q_reg ( .D(WX6955), .SI(test_si56), .SE(test_se), .CLK(CK), 
        .Q(n8467), .QN(n3907) );
  SDFFX1 DFF_964_Q_reg ( .D(WX6957), .SI(n8467), .SE(test_se), .CLK(CK), .Q(
        n8466), .QN(n3906) );
  SDFFX1 DFF_965_Q_reg ( .D(WX6959), .SI(n8466), .SE(test_se), .CLK(CK), .Q(
        n8465), .QN(n3905) );
  SDFFX1 DFF_966_Q_reg ( .D(WX6961), .SI(n8465), .SE(test_se), .CLK(CK), .Q(
        n8464), .QN(n3904) );
  SDFFX1 DFF_967_Q_reg ( .D(WX6963), .SI(n8464), .SE(test_se), .CLK(CK), .Q(
        n8463), .QN(n3903) );
  SDFFX1 DFF_968_Q_reg ( .D(WX6965), .SI(n8463), .SE(test_se), .CLK(CK), .Q(
        n8462), .QN(n3902) );
  SDFFX1 DFF_969_Q_reg ( .D(WX6967), .SI(n8462), .SE(test_se), .CLK(CK), .Q(
        n8461), .QN(n3901) );
  SDFFX1 DFF_970_Q_reg ( .D(WX6969), .SI(n8461), .SE(test_se), .CLK(CK), .Q(
        n8460), .QN(n3900) );
  SDFFX1 DFF_971_Q_reg ( .D(WX6971), .SI(n8460), .SE(test_se), .CLK(CK), .Q(
        n8459), .QN(n3899) );
  SDFFX1 DFF_972_Q_reg ( .D(WX6973), .SI(n8459), .SE(test_se), .CLK(CK), .Q(
        n8458), .QN(n3898) );
  SDFFX1 DFF_973_Q_reg ( .D(WX6975), .SI(n8458), .SE(test_se), .CLK(CK), .Q(
        n8457), .QN(n3897) );
  SDFFX1 DFF_974_Q_reg ( .D(WX6977), .SI(n8457), .SE(test_se), .CLK(CK), .Q(
        n8456), .QN(n3896) );
  SDFFX1 DFF_975_Q_reg ( .D(WX6979), .SI(n8456), .SE(test_se), .CLK(CK), .Q(
        n8455), .QN(n3895) );
  SDFFX1 DFF_976_Q_reg ( .D(WX6981), .SI(n8455), .SE(test_se), .CLK(CK), .Q(
        n8454), .QN(n3894) );
  SDFFX1 DFF_977_Q_reg ( .D(WX6983), .SI(n8454), .SE(test_se), .CLK(CK), .Q(
        n8453), .QN(n3893) );
  SDFFX1 DFF_978_Q_reg ( .D(WX6985), .SI(n8453), .SE(test_se), .CLK(CK), .Q(
        n8452), .QN(n3892) );
  SDFFX1 DFF_979_Q_reg ( .D(WX6987), .SI(n8452), .SE(test_se), .CLK(CK), .Q(
        test_so56), .QN(n3891) );
  SDFFX1 DFF_980_Q_reg ( .D(WX6989), .SI(test_si57), .SE(test_se), .CLK(CK), 
        .Q(n8449), .QN(n3890) );
  SDFFX1 DFF_981_Q_reg ( .D(WX6991), .SI(n8449), .SE(test_se), .CLK(CK), .Q(
        n8448), .QN(n3889) );
  SDFFX1 DFF_982_Q_reg ( .D(WX6993), .SI(n8448), .SE(test_se), .CLK(CK), .Q(
        n8447), .QN(n3888) );
  SDFFX1 DFF_983_Q_reg ( .D(WX6995), .SI(n8447), .SE(test_se), .CLK(CK), .Q(
        n8446), .QN(n3887) );
  SDFFX1 DFF_984_Q_reg ( .D(WX6997), .SI(n8446), .SE(test_se), .CLK(CK), .Q(
        n8445), .QN(n3886) );
  SDFFX1 DFF_985_Q_reg ( .D(WX6999), .SI(n8445), .SE(test_se), .CLK(CK), .Q(
        n8444), .QN(n3885) );
  SDFFX1 DFF_986_Q_reg ( .D(WX7001), .SI(n8444), .SE(test_se), .CLK(CK), .Q(
        n8443), .QN(n3884) );
  SDFFX1 DFF_987_Q_reg ( .D(WX7003), .SI(n8443), .SE(test_se), .CLK(CK), .Q(
        n8442), .QN(n3883) );
  SDFFX1 DFF_988_Q_reg ( .D(WX7005), .SI(n8442), .SE(test_se), .CLK(CK), .Q(
        n8441), .QN(n3882) );
  SDFFX1 DFF_989_Q_reg ( .D(WX7007), .SI(n8441), .SE(test_se), .CLK(CK), .Q(
        n8440), .QN(n3881) );
  SDFFX1 DFF_990_Q_reg ( .D(WX7009), .SI(n8440), .SE(test_se), .CLK(CK), .Q(
        n8439), .QN(n3880) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(test_se), .CLK(CK), .Q(
        n8438), .QN(n3879) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(test_se), .CLK(CK), .Q(
        n8437), .QN(n3341) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(test_se), .CLK(CK), .Q(
        n8436), .QN(n3405) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(test_se), .CLK(CK), .Q(
        n8435), .QN(n3404) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(test_se), .CLK(CK), .Q(
        n8434), .QN(n3403) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(test_se), .CLK(CK), .Q(
        test_so57), .QN(n3402) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(test_se), .CLK(CK), 
        .Q(n8431), .QN(n3401) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(test_se), .CLK(CK), .Q(
        n8430), .QN(n3400) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(test_se), .CLK(CK), .Q(
        n8429), .QN(n3399) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(test_se), .CLK(CK), .Q(
        n8428), .QN(n3398) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(test_se), .CLK(CK), .Q(
        n8427), .QN(n3397) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(test_se), .CLK(CK), .Q(
        n8426), .QN(n3396) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(test_se), .CLK(CK), .Q(
        n8425), .QN(n3395) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(test_se), .CLK(CK), .Q(
        n8424), .QN(n3394) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(test_se), .CLK(CK), .Q(
        n8423), .QN(n3393) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(test_se), .CLK(CK), .Q(
        n8422), .QN(n3392) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(test_se), .CLK(CK), .Q(
        n8421), .QN(n3391) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(test_se), .CLK(CK), .Q(
        WX7142), .QN() );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(test_se), .CLK(CK), .Q(
        WX7144), .QN() );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(test_se), .CLK(CK), .Q(
        WX7146), .QN() );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(test_se), .CLK(CK), .Q(
        WX7148), .QN() );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(test_se), .CLK(CK), .Q(
        WX7150), .QN() );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(test_se), .CLK(CK), .Q(
        test_so58), .QN() );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(test_se), .CLK(CK), 
        .Q(WX7154), .QN() );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(test_se), .CLK(CK), .Q(
        WX7156), .QN() );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(test_se), .CLK(CK), .Q(
        WX7158), .QN() );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(test_se), .CLK(CK), .Q(
        WX7160), .QN() );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(test_se), .CLK(CK), .Q(
        WX7162), .QN() );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(test_se), .CLK(CK), .Q(
        WX7164), .QN() );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(test_se), .CLK(CK), .Q(
        WX7166), .QN() );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(test_se), .CLK(CK), .Q(
        WX7168), .QN() );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(test_se), .CLK(CK), .Q(
        WX7170), .QN() );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(test_se), .CLK(CK), .Q(
        WX7172), .QN() );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(test_se), .CLK(CK), .Q(
        WX7174), .QN() );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(test_se), .CLK(CK), .Q(
        WX7176), .QN() );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(test_se), .CLK(CK), .Q(
        WX7178), .QN() );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(test_se), .CLK(CK), .Q(
        WX7180), .QN() );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(test_se), .CLK(CK), .Q(
        WX7182), .QN() );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(test_se), .CLK(CK), .Q(
        WX7184), .QN() );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(test_se), .CLK(CK), .Q(
        test_so59), .QN() );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(test_se), .CLK(CK), 
        .Q(WX7188), .QN() );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(test_se), .CLK(CK), .Q(
        WX7190), .QN() );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(test_se), .CLK(CK), .Q(
        WX7192), .QN() );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(test_se), .CLK(CK), .Q(
        WX7194), .QN() );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(test_se), .CLK(CK), .Q(
        WX7196), .QN() );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(test_se), .CLK(CK), .Q(
        WX7198), .QN() );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(test_se), .CLK(CK), .Q(
        WX7200), .QN() );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(test_se), .CLK(CK), .Q(
        WX7202), .QN() );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(test_se), .CLK(CK), .Q(
        WX7204), .QN() );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(test_se), .CLK(CK), .Q(
        WX7206), .QN(n3657) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(test_se), .CLK(CK), .Q(
        WX7208), .QN(n3655) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(test_se), .CLK(CK), .Q(
        WX7210), .QN(n3653) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(test_se), .CLK(CK), .Q(
        WX7212), .QN(n3651) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(test_se), .CLK(CK), .Q(
        WX7214), .QN(n3649) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(test_se), .CLK(CK), .Q(
        WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(test_se), .CLK(CK), .Q(
        WX7218), .QN(n3645) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(test_se), .CLK(CK), .Q(
        test_so60), .QN(n3643) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(test_se), .CLK(CK), 
        .Q(WX7222), .QN(n3641) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(test_se), .CLK(CK), .Q(
        WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(test_se), .CLK(CK), .Q(
        WX7226), .QN(n3637) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(test_se), .CLK(CK), .Q(
        WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(test_se), .CLK(CK), .Q(
        WX7230), .QN(n3633) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(test_se), .CLK(CK), .Q(
        WX7232), .QN(n3631) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(test_se), .CLK(CK), .Q(
        WX7234), .QN(n3629) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(test_se), .CLK(CK), .Q(
        WX7236), .QN(n3627) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(test_se), .CLK(CK), .Q(
        WX7238), .QN() );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(test_se), .CLK(CK), .Q(
        WX7240), .QN() );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(test_se), .CLK(CK), .Q(
        WX7242), .QN() );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(test_se), .CLK(CK), .Q(
        WX7244), .QN() );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(test_se), .CLK(CK), .Q(
        WX7246), .QN() );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(test_se), .CLK(CK), .Q(
        WX7248), .QN() );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(test_se), .CLK(CK), .Q(
        WX7250), .QN() );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(test_se), .CLK(CK), .Q(
        WX7252), .QN() );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(test_se), .CLK(CK), .Q(
        test_so61), .QN() );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(test_se), .CLK(CK), 
        .Q(WX7256), .QN() );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(test_se), .CLK(CK), .Q(
        WX7258), .QN() );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(test_se), .CLK(CK), .Q(
        WX7260), .QN() );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(test_se), .CLK(CK), .Q(
        WX7262), .QN() );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(test_se), .CLK(CK), .Q(
        WX7264), .QN() );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(test_se), .CLK(CK), .Q(
        WX7266), .QN() );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(test_se), .CLK(CK), .Q(
        WX7268), .QN() );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(test_se), .CLK(CK), .Q(
        WX7270), .QN() );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(test_se), .CLK(CK), .Q(
        WX7272), .QN() );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(test_se), .CLK(CK), .Q(
        WX7274), .QN() );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(test_se), .CLK(CK), .Q(
        WX7276), .QN() );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(test_se), .CLK(CK), .Q(
        WX7278), .QN() );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(test_se), .CLK(CK), .Q(
        WX7280), .QN() );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(test_se), .CLK(CK), .Q(
        WX7282), .QN() );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(test_se), .CLK(CK), .Q(
        WX7284), .QN() );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(test_se), .CLK(CK), .Q(
        WX7286), .QN() );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(test_se), .CLK(CK), .Q(
        test_so62), .QN() );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(test_se), .CLK(CK), 
        .Q(WX7290), .QN() );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(test_se), .CLK(CK), .Q(
        WX7292), .QN() );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(test_se), .CLK(CK), .Q(
        WX7294), .QN() );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(test_se), .CLK(CK), .Q(
        WX7296), .QN() );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(test_se), .CLK(CK), .Q(
        WX7298), .QN() );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(test_se), .CLK(CK), .Q(
        WX7300), .QN() );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(test_se), .CLK(CK), .Q(
        WX7302), .QN() );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(test_se), .CLK(CK), .Q(
        WX7304), .QN() );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(test_se), .CLK(CK), .Q(
        WX7306), .QN() );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(test_se), .CLK(CK), .Q(
        WX7308), .QN() );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(test_se), .CLK(CK), .Q(
        WX7310), .QN() );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(test_se), .CLK(CK), .Q(
        WX7312), .QN() );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(test_se), .CLK(CK), .Q(
        WX7314), .QN() );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(test_se), .CLK(CK), .Q(
        WX7316), .QN() );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(test_se), .CLK(CK), .Q(
        WX7318), .QN() );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(test_se), .CLK(CK), .Q(
        WX7320), .QN() );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(test_se), .CLK(CK), .Q(
        test_so63), .QN() );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(test_se), .CLK(CK), 
        .Q(WX7324), .QN() );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(test_se), .CLK(CK), .Q(
        WX7326), .QN() );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(test_se), .CLK(CK), .Q(
        WX7328), .QN() );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(test_se), .CLK(CK), .Q(
        WX7330), .QN() );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(test_se), .CLK(CK), .Q(
        WX7332), .QN() );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(test_se), .CLK(CK), .Q(
        WX7334), .QN() );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(test_se), .CLK(CK), .Q(
        WX7336), .QN() );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(test_se), .CLK(CK), .Q(
        WX7338), .QN() );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(test_se), .CLK(CK), .Q(
        WX7340), .QN() );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(test_se), .CLK(CK), .Q(
        WX7342), .QN() );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(test_se), .CLK(CK), .Q(
        WX7344), .QN() );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(test_se), .CLK(CK), .Q(
        WX7346), .QN() );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(test_se), .CLK(CK), .Q(
        WX7348), .QN() );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(test_se), .CLK(CK), .Q(
        WX7350), .QN() );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(test_se), .CLK(CK), .Q(
        WX7352), .QN() );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(test_se), .CLK(CK), .Q(
        WX7354), .QN() );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(test_se), .CLK(CK), .Q(
        test_so64), .QN() );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(test_se), .CLK(CK), 
        .Q(WX7358), .QN() );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(test_se), .CLK(CK), .Q(
        WX7360), .QN() );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(test_se), .CLK(CK), .Q(
        WX7362), .QN() );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(test_se), .CLK(CK), .Q(
        WX7364), .QN() );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_12), .QN(DFF_1132_n1) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_29), .QN(DFF_1149_n1) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(test_se), .CLK(CK), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(WX8242), .SI(CRC_OUT_4_31), .SE(test_se), .CLK(CK), .Q(WX8243), .QN() );
  SDFFX1 DFF_1153_Q_reg ( .D(WX8244), .SI(WX8243), .SE(test_se), .CLK(CK), .Q(
        n8411), .QN(n3878) );
  SDFFX1 DFF_1154_Q_reg ( .D(WX8246), .SI(n8411), .SE(test_se), .CLK(CK), .Q(
        n8410), .QN(n3877) );
  SDFFX1 DFF_1155_Q_reg ( .D(WX8248), .SI(n8410), .SE(test_se), .CLK(CK), .Q(
        n8409), .QN(n3876) );
  SDFFX1 DFF_1156_Q_reg ( .D(WX8250), .SI(n8409), .SE(test_se), .CLK(CK), .Q(
        n8408), .QN(n3875) );
  SDFFX1 DFF_1157_Q_reg ( .D(WX8252), .SI(n8408), .SE(test_se), .CLK(CK), .Q(
        n8407), .QN(n3874) );
  SDFFX1 DFF_1158_Q_reg ( .D(WX8254), .SI(n8407), .SE(test_se), .CLK(CK), .Q(
        n8406), .QN(n3873) );
  SDFFX1 DFF_1159_Q_reg ( .D(WX8256), .SI(n8406), .SE(test_se), .CLK(CK), .Q(
        n8405), .QN(n3872) );
  SDFFX1 DFF_1160_Q_reg ( .D(WX8258), .SI(n8405), .SE(test_se), .CLK(CK), .Q(
        n8404), .QN(n3871) );
  SDFFX1 DFF_1161_Q_reg ( .D(WX8260), .SI(n8404), .SE(test_se), .CLK(CK), .Q(
        n8403), .QN(n3870) );
  SDFFX1 DFF_1162_Q_reg ( .D(WX8262), .SI(n8403), .SE(test_se), .CLK(CK), .Q(
        n8402), .QN(n3869) );
  SDFFX1 DFF_1163_Q_reg ( .D(WX8264), .SI(n8402), .SE(test_se), .CLK(CK), .Q(
        n8401), .QN(n3868) );
  SDFFX1 DFF_1164_Q_reg ( .D(WX8266), .SI(n8401), .SE(test_se), .CLK(CK), .Q(
        n8400), .QN(n3867) );
  SDFFX1 DFF_1165_Q_reg ( .D(WX8268), .SI(n8400), .SE(test_se), .CLK(CK), .Q(
        n8399), .QN(n3866) );
  SDFFX1 DFF_1166_Q_reg ( .D(WX8270), .SI(n8399), .SE(test_se), .CLK(CK), .Q(
        test_so67), .QN(n3865) );
  SDFFX1 DFF_1167_Q_reg ( .D(WX8272), .SI(test_si68), .SE(test_se), .CLK(CK), 
        .Q(n8396), .QN(n3864) );
  SDFFX1 DFF_1168_Q_reg ( .D(WX8274), .SI(n8396), .SE(test_se), .CLK(CK), .Q(
        n8395), .QN(n3863) );
  SDFFX1 DFF_1169_Q_reg ( .D(WX8276), .SI(n8395), .SE(test_se), .CLK(CK), .Q(
        n8394), .QN(n3862) );
  SDFFX1 DFF_1170_Q_reg ( .D(WX8278), .SI(n8394), .SE(test_se), .CLK(CK), .Q(
        n8393), .QN(n3861) );
  SDFFX1 DFF_1171_Q_reg ( .D(WX8280), .SI(n8393), .SE(test_se), .CLK(CK), .Q(
        n8392), .QN(n3860) );
  SDFFX1 DFF_1172_Q_reg ( .D(WX8282), .SI(n8392), .SE(test_se), .CLK(CK), .Q(
        n8391), .QN(n3859) );
  SDFFX1 DFF_1173_Q_reg ( .D(WX8284), .SI(n8391), .SE(test_se), .CLK(CK), .Q(
        n8390), .QN(n3858) );
  SDFFX1 DFF_1174_Q_reg ( .D(WX8286), .SI(n8390), .SE(test_se), .CLK(CK), .Q(
        n8389), .QN(n3857) );
  SDFFX1 DFF_1175_Q_reg ( .D(WX8288), .SI(n8389), .SE(test_se), .CLK(CK), .Q(
        n8388), .QN(n3856) );
  SDFFX1 DFF_1176_Q_reg ( .D(WX8290), .SI(n8388), .SE(test_se), .CLK(CK), .Q(
        n8387), .QN(n3855) );
  SDFFX1 DFF_1177_Q_reg ( .D(WX8292), .SI(n8387), .SE(test_se), .CLK(CK), .Q(
        n8386), .QN(n3854) );
  SDFFX1 DFF_1178_Q_reg ( .D(WX8294), .SI(n8386), .SE(test_se), .CLK(CK), .Q(
        n8385), .QN(n3853) );
  SDFFX1 DFF_1179_Q_reg ( .D(WX8296), .SI(n8385), .SE(test_se), .CLK(CK), .Q(
        n8384), .QN(n3852) );
  SDFFX1 DFF_1180_Q_reg ( .D(WX8298), .SI(n8384), .SE(test_se), .CLK(CK), .Q(
        n8383), .QN(n3851) );
  SDFFX1 DFF_1181_Q_reg ( .D(WX8300), .SI(n8383), .SE(test_se), .CLK(CK), .Q(
        n8382), .QN(n3850) );
  SDFFX1 DFF_1182_Q_reg ( .D(WX8302), .SI(n8382), .SE(test_se), .CLK(CK), .Q(
        n8381), .QN(n3849) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(test_se), .CLK(CK), .Q(
        test_so68), .QN(n3848) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(test_se), .CLK(CK), 
        .Q(n8378), .QN(n3340) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(test_se), .CLK(CK), .Q(
        n8377), .QN(n3390) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(test_se), .CLK(CK), .Q(
        n8376), .QN(n3389) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(test_se), .CLK(CK), .Q(
        n8375), .QN(n3388) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(test_se), .CLK(CK), .Q(
        n8374), .QN(n3387) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(test_se), .CLK(CK), .Q(
        n8373), .QN(n3386) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(test_se), .CLK(CK), .Q(
        n8372), .QN(n3385) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(test_se), .CLK(CK), .Q(
        n8371), .QN(n3384) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(test_se), .CLK(CK), .Q(
        n8370), .QN(n3383) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(test_se), .CLK(CK), .Q(
        n8369), .QN(n3382) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(test_se), .CLK(CK), .Q(
        n8368), .QN(n3381) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(test_se), .CLK(CK), .Q(
        n8367), .QN(n3380) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(test_se), .CLK(CK), .Q(
        n8366), .QN(n3379) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(test_se), .CLK(CK), .Q(
        n8365), .QN(n3378) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(test_se), .CLK(CK), .Q(
        n8364), .QN(n3377) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(test_se), .CLK(CK), .Q(
        n8363), .QN(n3376) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(test_se), .CLK(CK), .Q(
        test_so69), .QN() );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(test_se), .CLK(CK), 
        .Q(WX8437), .QN() );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(test_se), .CLK(CK), .Q(
        WX8439), .QN() );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(test_se), .CLK(CK), .Q(
        WX8441), .QN() );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(test_se), .CLK(CK), .Q(
        WX8443), .QN() );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(test_se), .CLK(CK), .Q(
        WX8445), .QN() );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(test_se), .CLK(CK), .Q(
        WX8447), .QN() );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(test_se), .CLK(CK), .Q(
        WX8449), .QN() );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(test_se), .CLK(CK), .Q(
        WX8451), .QN() );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(test_se), .CLK(CK), .Q(
        WX8453), .QN() );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(test_se), .CLK(CK), .Q(
        WX8455), .QN() );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(test_se), .CLK(CK), .Q(
        WX8457), .QN() );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(test_se), .CLK(CK), .Q(
        WX8459), .QN() );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(test_se), .CLK(CK), .Q(
        WX8461), .QN() );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(test_se), .CLK(CK), .Q(
        WX8463), .QN() );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(test_se), .CLK(CK), .Q(
        WX8465), .QN() );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(test_se), .CLK(CK), .Q(
        WX8467), .QN() );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(test_se), .CLK(CK), .Q(
        test_so70), .QN() );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(test_se), .CLK(CK), 
        .Q(WX8471), .QN() );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(test_se), .CLK(CK), .Q(
        WX8473), .QN() );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(test_se), .CLK(CK), .Q(
        WX8475), .QN() );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(test_se), .CLK(CK), .Q(
        WX8477), .QN() );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(test_se), .CLK(CK), .Q(
        WX8479), .QN() );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(test_se), .CLK(CK), .Q(
        WX8481), .QN() );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(test_se), .CLK(CK), .Q(
        WX8483), .QN() );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(test_se), .CLK(CK), .Q(
        WX8485), .QN() );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(test_se), .CLK(CK), .Q(
        WX8487), .QN() );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(test_se), .CLK(CK), .Q(
        WX8489), .QN() );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(test_se), .CLK(CK), .Q(
        WX8491), .QN() );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(test_se), .CLK(CK), .Q(
        WX8493), .QN() );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(test_se), .CLK(CK), .Q(
        WX8495), .QN() );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(test_se), .CLK(CK), .Q(
        WX8497), .QN() );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(test_se), .CLK(CK), .Q(
        WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(test_se), .CLK(CK), .Q(
        WX8501), .QN(n3623) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(test_se), .CLK(CK), .Q(
        test_so71), .QN(n3621) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(test_se), .CLK(CK), 
        .Q(WX8505), .QN(n3619) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(test_se), .CLK(CK), .Q(
        WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(test_se), .CLK(CK), .Q(
        WX8509), .QN(n3615) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(test_se), .CLK(CK), .Q(
        WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(test_se), .CLK(CK), .Q(
        WX8513), .QN(n3611) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(test_se), .CLK(CK), .Q(
        WX8515), .QN(n3609) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(test_se), .CLK(CK), .Q(
        WX8517), .QN(n3607) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(test_se), .CLK(CK), .Q(
        WX8519), .QN(n3605) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(test_se), .CLK(CK), .Q(
        WX8521), .QN(n3603) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(test_se), .CLK(CK), .Q(
        WX8523), .QN(n3601) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(test_se), .CLK(CK), .Q(
        WX8525), .QN(n3599) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(test_se), .CLK(CK), .Q(
        WX8527), .QN(n3597) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(test_se), .CLK(CK), .Q(
        WX8529), .QN(n3595) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(test_se), .CLK(CK), .Q(
        WX8531), .QN() );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(test_se), .CLK(CK), .Q(
        WX8533), .QN() );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(test_se), .CLK(CK), .Q(
        WX8535), .QN() );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(test_se), .CLK(CK), .Q(
        test_so72), .QN() );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(test_se), .CLK(CK), 
        .Q(WX8539), .QN() );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(test_se), .CLK(CK), .Q(
        WX8541), .QN() );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(test_se), .CLK(CK), .Q(
        WX8543), .QN() );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(test_se), .CLK(CK), .Q(
        WX8545), .QN() );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(test_se), .CLK(CK), .Q(
        WX8547), .QN() );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(test_se), .CLK(CK), .Q(
        WX8549), .QN() );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(test_se), .CLK(CK), .Q(
        WX8551), .QN() );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(test_se), .CLK(CK), .Q(
        WX8553), .QN() );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(test_se), .CLK(CK), .Q(
        WX8555), .QN() );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(test_se), .CLK(CK), .Q(
        WX8557), .QN() );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(test_se), .CLK(CK), .Q(
        WX8559), .QN() );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(test_se), .CLK(CK), .Q(
        WX8561), .QN() );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(test_se), .CLK(CK), .Q(
        WX8563), .QN() );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(test_se), .CLK(CK), .Q(
        WX8565), .QN() );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(test_se), .CLK(CK), .Q(
        WX8567), .QN() );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(test_se), .CLK(CK), .Q(
        WX8569), .QN() );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(test_se), .CLK(CK), .Q(
        test_so73), .QN() );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(test_se), .CLK(CK), 
        .Q(WX8573), .QN() );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(test_se), .CLK(CK), .Q(
        WX8575), .QN() );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(test_se), .CLK(CK), .Q(
        WX8577), .QN() );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(test_se), .CLK(CK), .Q(
        WX8579), .QN() );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(test_se), .CLK(CK), .Q(
        WX8581), .QN() );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(test_se), .CLK(CK), .Q(
        WX8583), .QN() );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(test_se), .CLK(CK), .Q(
        WX8585), .QN() );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(test_se), .CLK(CK), .Q(
        WX8587), .QN() );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(test_se), .CLK(CK), .Q(
        WX8589), .QN() );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(test_se), .CLK(CK), .Q(
        WX8591), .QN() );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(test_se), .CLK(CK), .Q(
        WX8593), .QN() );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(test_se), .CLK(CK), .Q(
        WX8595), .QN() );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(test_se), .CLK(CK), .Q(
        WX8597), .QN() );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(test_se), .CLK(CK), .Q(
        WX8599), .QN() );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(test_se), .CLK(CK), .Q(
        WX8601), .QN() );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(test_se), .CLK(CK), .Q(
        WX8603), .QN() );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(test_se), .CLK(CK), .Q(
        test_so74), .QN() );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(test_se), .CLK(CK), 
        .Q(WX8607), .QN() );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(test_se), .CLK(CK), .Q(
        WX8609), .QN() );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(test_se), .CLK(CK), .Q(
        WX8611), .QN() );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(test_se), .CLK(CK), .Q(
        WX8613), .QN() );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(test_se), .CLK(CK), .Q(
        WX8615), .QN() );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(test_se), .CLK(CK), .Q(
        WX8617), .QN() );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(test_se), .CLK(CK), .Q(
        WX8619), .QN() );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(test_se), .CLK(CK), .Q(
        WX8621), .QN() );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(test_se), .CLK(CK), .Q(
        WX8623), .QN() );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(test_se), .CLK(CK), .Q(
        WX8625), .QN() );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(test_se), .CLK(CK), .Q(
        WX8627), .QN() );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(test_se), .CLK(CK), .Q(
        WX8629), .QN() );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(test_se), .CLK(CK), .Q(
        WX8631), .QN() );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(test_se), .CLK(CK), .Q(
        WX8633), .QN() );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(test_se), .CLK(CK), .Q(
        WX8635), .QN() );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(test_se), .CLK(CK), .Q(
        WX8637), .QN() );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(test_se), .CLK(CK), .Q(
        test_so75), .QN() );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(test_se), .CLK(CK), 
        .Q(WX8641), .QN() );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(test_se), .CLK(CK), .Q(
        WX8643), .QN() );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(test_se), .CLK(CK), .Q(
        WX8645), .QN() );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(test_se), .CLK(CK), .Q(
        WX8647), .QN() );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(test_se), .CLK(CK), .Q(
        WX8649), .QN() );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(test_se), .CLK(CK), .Q(
        WX8651), .QN() );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(test_se), .CLK(CK), .Q(
        WX8653), .QN() );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(test_se), .CLK(CK), .Q(
        WX8655), .QN() );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(test_se), .CLK(CK), .Q(
        WX8657), .QN() );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(test_se), .CLK(CK), .Q(
        CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_7), .QN(DFF_1319_n1) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_24), .QN(DFF_1336_n1) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(test_se), .CLK(CK), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(WX9535), .SI(CRC_OUT_3_31), .SE(test_se), .CLK(CK), .Q(WX9536), .QN() );
  SDFFX1 DFF_1345_Q_reg ( .D(WX9537), .SI(WX9536), .SE(test_se), .CLK(CK), .Q(
        n8353), .QN(n3847) );
  SDFFX1 DFF_1346_Q_reg ( .D(WX9539), .SI(n8353), .SE(test_se), .CLK(CK), .Q(
        n8352), .QN(n3846) );
  SDFFX1 DFF_1347_Q_reg ( .D(WX9541), .SI(n8352), .SE(test_se), .CLK(CK), .Q(
        n8351), .QN(n3845) );
  SDFFX1 DFF_1348_Q_reg ( .D(WX9543), .SI(n8351), .SE(test_se), .CLK(CK), .Q(
        n8350), .QN(n3844) );
  SDFFX1 DFF_1349_Q_reg ( .D(WX9545), .SI(n8350), .SE(test_se), .CLK(CK), .Q(
        n8349), .QN(n3843) );
  SDFFX1 DFF_1350_Q_reg ( .D(WX9547), .SI(n8349), .SE(test_se), .CLK(CK), .Q(
        n8348), .QN(n3842) );
  SDFFX1 DFF_1351_Q_reg ( .D(WX9549), .SI(n8348), .SE(test_se), .CLK(CK), .Q(
        n8347), .QN(n3841) );
  SDFFX1 DFF_1352_Q_reg ( .D(WX9551), .SI(n8347), .SE(test_se), .CLK(CK), .Q(
        n8346), .QN(n3840) );
  SDFFX1 DFF_1353_Q_reg ( .D(WX9553), .SI(n8346), .SE(test_se), .CLK(CK), .Q(
        test_so78), .QN(n3839) );
  SDFFX1 DFF_1354_Q_reg ( .D(WX9555), .SI(test_si79), .SE(test_se), .CLK(CK), 
        .Q(n8343), .QN(n3838) );
  SDFFX1 DFF_1355_Q_reg ( .D(WX9557), .SI(n8343), .SE(test_se), .CLK(CK), .Q(
        n8342), .QN(n3837) );
  SDFFX1 DFF_1356_Q_reg ( .D(WX9559), .SI(n8342), .SE(test_se), .CLK(CK), .Q(
        n8341), .QN(n3836) );
  SDFFX1 DFF_1357_Q_reg ( .D(WX9561), .SI(n8341), .SE(test_se), .CLK(CK), .Q(
        n8340), .QN(n3835) );
  SDFFX1 DFF_1358_Q_reg ( .D(WX9563), .SI(n8340), .SE(test_se), .CLK(CK), .Q(
        n8339), .QN(n3834) );
  SDFFX1 DFF_1359_Q_reg ( .D(WX9565), .SI(n8339), .SE(test_se), .CLK(CK), .Q(
        n8338), .QN(n3833) );
  SDFFX1 DFF_1360_Q_reg ( .D(WX9567), .SI(n8338), .SE(test_se), .CLK(CK), .Q(
        n8337), .QN(n3832) );
  SDFFX1 DFF_1361_Q_reg ( .D(WX9569), .SI(n8337), .SE(test_se), .CLK(CK), .Q(
        n8336), .QN(n3831) );
  SDFFX1 DFF_1362_Q_reg ( .D(WX9571), .SI(n8336), .SE(test_se), .CLK(CK), .Q(
        n8335), .QN(n3830) );
  SDFFX1 DFF_1363_Q_reg ( .D(WX9573), .SI(n8335), .SE(test_se), .CLK(CK), .Q(
        n8334), .QN(n3829) );
  SDFFX1 DFF_1364_Q_reg ( .D(WX9575), .SI(n8334), .SE(test_se), .CLK(CK), .Q(
        n8333), .QN(n3828) );
  SDFFX1 DFF_1365_Q_reg ( .D(WX9577), .SI(n8333), .SE(test_se), .CLK(CK), .Q(
        n8332), .QN(n3827) );
  SDFFX1 DFF_1366_Q_reg ( .D(WX9579), .SI(n8332), .SE(test_se), .CLK(CK), .Q(
        n8331), .QN(n3826) );
  SDFFX1 DFF_1367_Q_reg ( .D(WX9581), .SI(n8331), .SE(test_se), .CLK(CK), .Q(
        n8330), .QN(n3825) );
  SDFFX1 DFF_1368_Q_reg ( .D(WX9583), .SI(n8330), .SE(test_se), .CLK(CK), .Q(
        n8329), .QN(n3824) );
  SDFFX1 DFF_1369_Q_reg ( .D(WX9585), .SI(n8329), .SE(test_se), .CLK(CK), .Q(
        n8328), .QN(n3823) );
  SDFFX1 DFF_1370_Q_reg ( .D(WX9587), .SI(n8328), .SE(test_se), .CLK(CK), .Q(
        test_so79), .QN(n3822) );
  SDFFX1 DFF_1371_Q_reg ( .D(WX9589), .SI(test_si80), .SE(test_se), .CLK(CK), 
        .Q(n8325), .QN(n3821) );
  SDFFX1 DFF_1372_Q_reg ( .D(WX9591), .SI(n8325), .SE(test_se), .CLK(CK), .Q(
        n8324), .QN(n3820) );
  SDFFX1 DFF_1373_Q_reg ( .D(WX9593), .SI(n8324), .SE(test_se), .CLK(CK), .Q(
        n8323), .QN(n3819) );
  SDFFX1 DFF_1374_Q_reg ( .D(WX9595), .SI(n8323), .SE(test_se), .CLK(CK), .Q(
        n8322), .QN(n3818) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(test_se), .CLK(CK), .Q(
        n8321), .QN(n3817) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(test_se), .CLK(CK), .Q(
        n8320), .QN(n3339) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(test_se), .CLK(CK), .Q(
        n8319), .QN(n3375) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(test_se), .CLK(CK), .Q(
        n8318), .QN(n3374) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(test_se), .CLK(CK), .Q(
        n8317), .QN(n3373) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(test_se), .CLK(CK), .Q(
        n8316), .QN(n3372) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(test_se), .CLK(CK), .Q(
        n8315), .QN(n3371) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(test_se), .CLK(CK), .Q(
        n8314), .QN(n3370) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(test_se), .CLK(CK), .Q(
        n8313), .QN(n3369) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(test_se), .CLK(CK), .Q(
        n8312), .QN(n3368) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(test_se), .CLK(CK), .Q(
        n8311), .QN(n3367) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(test_se), .CLK(CK), .Q(
        n8310), .QN(n3366) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(test_se), .CLK(CK), .Q(
        test_so80), .QN(n3365) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(test_se), .CLK(CK), 
        .Q(n8307), .QN(n3364) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(test_se), .CLK(CK), .Q(
        n8306), .QN(n3363) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(test_se), .CLK(CK), .Q(
        n8305), .QN(n3362) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(test_se), .CLK(CK), .Q(
        n8304), .QN(n3361) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(test_se), .CLK(CK), .Q(
        WX9728), .QN() );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(test_se), .CLK(CK), .Q(
        WX9730), .QN() );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(test_se), .CLK(CK), .Q(
        WX9732), .QN() );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(test_se), .CLK(CK), .Q(
        WX9734), .QN() );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(test_se), .CLK(CK), .Q(
        WX9736), .QN() );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(test_se), .CLK(CK), .Q(
        WX9738), .QN() );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(test_se), .CLK(CK), .Q(
        WX9740), .QN() );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(test_se), .CLK(CK), .Q(
        WX9742), .QN() );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(test_se), .CLK(CK), .Q(
        WX9744), .QN() );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(test_se), .CLK(CK), .Q(
        WX9746), .QN() );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(test_se), .CLK(CK), .Q(
        WX9748), .QN() );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(test_se), .CLK(CK), .Q(
        WX9750), .QN() );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(test_se), .CLK(CK), .Q(
        test_so81), .QN() );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(test_se), .CLK(CK), 
        .Q(WX9754), .QN() );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(test_se), .CLK(CK), .Q(
        WX9756), .QN() );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(test_se), .CLK(CK), .Q(
        WX9758), .QN() );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(test_se), .CLK(CK), .Q(
        WX9760), .QN() );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(test_se), .CLK(CK), .Q(
        WX9762), .QN() );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(test_se), .CLK(CK), .Q(
        WX9764), .QN() );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(test_se), .CLK(CK), .Q(
        WX9766), .QN() );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(test_se), .CLK(CK), .Q(
        WX9768), .QN() );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(test_se), .CLK(CK), .Q(
        WX9770), .QN() );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(test_se), .CLK(CK), .Q(
        WX9772), .QN() );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(test_se), .CLK(CK), .Q(
        WX9774), .QN() );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(test_se), .CLK(CK), .Q(
        WX9776), .QN() );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(test_se), .CLK(CK), .Q(
        WX9778), .QN() );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(test_se), .CLK(CK), .Q(
        WX9780), .QN() );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(test_se), .CLK(CK), .Q(
        WX9782), .QN() );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(test_se), .CLK(CK), .Q(
        WX9784), .QN() );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(test_se), .CLK(CK), .Q(
        test_so82), .QN() );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(test_se), .CLK(CK), 
        .Q(WX9788), .QN() );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(test_se), .CLK(CK), .Q(
        WX9790), .QN() );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(test_se), .CLK(CK), .Q(
        WX9792), .QN(n3593) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(test_se), .CLK(CK), .Q(
        WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(test_se), .CLK(CK), .Q(
        WX9796), .QN(n3589) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(test_se), .CLK(CK), .Q(
        WX9798), .QN(n3587) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(test_se), .CLK(CK), .Q(
        WX9800), .QN(n3585) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(test_se), .CLK(CK), .Q(
        WX9802), .QN(n3583) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(test_se), .CLK(CK), .Q(
        WX9804), .QN(n3581) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(test_se), .CLK(CK), .Q(
        WX9806), .QN(n3579) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(test_se), .CLK(CK), .Q(
        WX9808), .QN(n3577) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(test_se), .CLK(CK), .Q(
        WX9810), .QN(n3575) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(test_se), .CLK(CK), .Q(
        WX9812), .QN(n3573) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(test_se), .CLK(CK), .Q(
        WX9814), .QN(n3571) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(test_se), .CLK(CK), .Q(
        WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(test_se), .CLK(CK), .Q(
        WX9818), .QN(n3567) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(test_se), .CLK(CK), .Q(
        test_so83), .QN(n3565) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(test_se), .CLK(CK), 
        .Q(WX9822), .QN(n3563) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(test_se), .CLK(CK), .Q(
        WX9824), .QN() );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(test_se), .CLK(CK), .Q(
        WX9826), .QN() );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(test_se), .CLK(CK), .Q(
        WX9828), .QN() );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(test_se), .CLK(CK), .Q(
        WX9830), .QN() );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(test_se), .CLK(CK), .Q(
        WX9832), .QN() );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(test_se), .CLK(CK), .Q(
        WX9834), .QN() );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(test_se), .CLK(CK), .Q(
        WX9836), .QN() );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(test_se), .CLK(CK), .Q(
        WX9838), .QN() );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(test_se), .CLK(CK), .Q(
        WX9840), .QN() );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(test_se), .CLK(CK), .Q(
        WX9842), .QN() );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(test_se), .CLK(CK), .Q(
        WX9844), .QN() );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(test_se), .CLK(CK), .Q(
        WX9846), .QN() );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(test_se), .CLK(CK), .Q(
        WX9848), .QN() );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(test_se), .CLK(CK), .Q(
        WX9850), .QN() );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(test_se), .CLK(CK), .Q(
        WX9852), .QN() );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(test_se), .CLK(CK), .Q(
        test_so84), .QN() );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(test_se), .CLK(CK), 
        .Q(WX9856), .QN() );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(test_se), .CLK(CK), .Q(
        WX9858), .QN() );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(test_se), .CLK(CK), .Q(
        WX9860), .QN() );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(test_se), .CLK(CK), .Q(
        WX9862), .QN() );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(test_se), .CLK(CK), .Q(
        WX9864), .QN() );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(test_se), .CLK(CK), .Q(
        WX9866), .QN() );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(test_se), .CLK(CK), .Q(
        WX9868), .QN() );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(test_se), .CLK(CK), .Q(
        WX9870), .QN() );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(test_se), .CLK(CK), .Q(
        WX9872), .QN() );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(test_se), .CLK(CK), .Q(
        WX9874), .QN() );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(test_se), .CLK(CK), .Q(
        WX9876), .QN() );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(test_se), .CLK(CK), .Q(
        WX9878), .QN() );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(test_se), .CLK(CK), .Q(
        WX9880), .QN() );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(test_se), .CLK(CK), .Q(
        WX9882), .QN() );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(test_se), .CLK(CK), .Q(
        WX9884), .QN() );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(test_se), .CLK(CK), .Q(
        WX9886), .QN() );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(test_se), .CLK(CK), .Q(
        test_so85), .QN() );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(test_se), .CLK(CK), 
        .Q(WX9890), .QN() );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(test_se), .CLK(CK), .Q(
        WX9892), .QN() );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(test_se), .CLK(CK), .Q(
        WX9894), .QN() );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(test_se), .CLK(CK), .Q(
        WX9896), .QN() );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(test_se), .CLK(CK), .Q(
        WX9898), .QN() );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(test_se), .CLK(CK), .Q(
        WX9900), .QN() );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(test_se), .CLK(CK), .Q(
        WX9902), .QN() );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(test_se), .CLK(CK), .Q(
        WX9904), .QN() );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(test_se), .CLK(CK), .Q(
        WX9906), .QN() );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(test_se), .CLK(CK), .Q(
        WX9908), .QN() );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(test_se), .CLK(CK), .Q(
        WX9910), .QN() );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(test_se), .CLK(CK), .Q(
        WX9912), .QN() );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(test_se), .CLK(CK), .Q(
        WX9914), .QN() );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(test_se), .CLK(CK), .Q(
        WX9916), .QN() );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(test_se), .CLK(CK), .Q(
        WX9918), .QN() );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(test_se), .CLK(CK), .Q(
        WX9920), .QN() );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(test_se), .CLK(CK), .Q(
        test_so86), .QN() );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(test_se), .CLK(CK), 
        .Q(WX9924), .QN() );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(test_se), .CLK(CK), .Q(
        WX9926), .QN() );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(test_se), .CLK(CK), .Q(
        WX9928), .QN() );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(test_se), .CLK(CK), .Q(
        WX9930), .QN() );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(test_se), .CLK(CK), .Q(
        WX9932), .QN() );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(test_se), .CLK(CK), .Q(
        WX9934), .QN() );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(test_se), .CLK(CK), .Q(
        WX9936), .QN() );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(test_se), .CLK(CK), .Q(
        WX9938), .QN() );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(test_se), .CLK(CK), .Q(
        WX9940), .QN() );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(test_se), .CLK(CK), .Q(
        WX9942), .QN() );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(test_se), .CLK(CK), .Q(
        WX9944), .QN() );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(test_se), .CLK(CK), .Q(
        WX9946), .QN() );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(test_se), .CLK(CK), .Q(
        WX9948), .QN() );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(test_se), .CLK(CK), .Q(
        WX9950), .QN() );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_2), .QN(DFF_1506_n1) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(test_se), .CLK(CK), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_19), .QN(DFF_1523_n1) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(WX10828), .SI(CRC_OUT_2_31), .SE(test_se), .CLK(
        CK), .Q(WX10829), .QN() );
  SDFFX1 DFF_1537_Q_reg ( .D(WX10830), .SI(WX10829), .SE(test_se), .CLK(CK), 
        .Q(n8295), .QN(n3816) );
  SDFFX1 DFF_1538_Q_reg ( .D(WX10832), .SI(n8295), .SE(test_se), .CLK(CK), .Q(
        n8294), .QN(n3815) );
  SDFFX1 DFF_1539_Q_reg ( .D(WX10834), .SI(n8294), .SE(test_se), .CLK(CK), .Q(
        n8293), .QN(n3814) );
  SDFFX1 DFF_1540_Q_reg ( .D(WX10836), .SI(n8293), .SE(test_se), .CLK(CK), .Q(
        test_so89), .QN(n3813) );
  SDFFX1 DFF_1541_Q_reg ( .D(WX10838), .SI(test_si90), .SE(test_se), .CLK(CK), 
        .Q(n8290), .QN(n3812) );
  SDFFX1 DFF_1542_Q_reg ( .D(WX10840), .SI(n8290), .SE(test_se), .CLK(CK), .Q(
        n8289), .QN(n3811) );
  SDFFX1 DFF_1543_Q_reg ( .D(WX10842), .SI(n8289), .SE(test_se), .CLK(CK), .Q(
        n8288), .QN(n3810) );
  SDFFX1 DFF_1544_Q_reg ( .D(WX10844), .SI(n8288), .SE(test_se), .CLK(CK), .Q(
        n8287), .QN(n3809) );
  SDFFX1 DFF_1545_Q_reg ( .D(WX10846), .SI(n8287), .SE(test_se), .CLK(CK), .Q(
        n8286), .QN(n3808) );
  SDFFX1 DFF_1546_Q_reg ( .D(WX10848), .SI(n8286), .SE(test_se), .CLK(CK), .Q(
        n8285), .QN(n3807) );
  SDFFX1 DFF_1547_Q_reg ( .D(WX10850), .SI(n8285), .SE(test_se), .CLK(CK), .Q(
        n8284), .QN(n3806) );
  SDFFX1 DFF_1548_Q_reg ( .D(WX10852), .SI(n8284), .SE(test_se), .CLK(CK), .Q(
        n8283), .QN(n3805) );
  SDFFX1 DFF_1549_Q_reg ( .D(WX10854), .SI(n8283), .SE(test_se), .CLK(CK), .Q(
        n8282), .QN(n3804) );
  SDFFX1 DFF_1550_Q_reg ( .D(WX10856), .SI(n8282), .SE(test_se), .CLK(CK), .Q(
        n8281), .QN(n3803) );
  SDFFX1 DFF_1551_Q_reg ( .D(WX10858), .SI(n8281), .SE(test_se), .CLK(CK), .Q(
        n8280), .QN(n3802) );
  SDFFX1 DFF_1552_Q_reg ( .D(WX10860), .SI(n8280), .SE(test_se), .CLK(CK), .Q(
        n8279), .QN(n3801) );
  SDFFX1 DFF_1553_Q_reg ( .D(WX10862), .SI(n8279), .SE(test_se), .CLK(CK), .Q(
        n8278), .QN(n3800) );
  SDFFX1 DFF_1554_Q_reg ( .D(WX10864), .SI(n8278), .SE(test_se), .CLK(CK), .Q(
        n8277), .QN(n3799) );
  SDFFX1 DFF_1555_Q_reg ( .D(WX10866), .SI(n8277), .SE(test_se), .CLK(CK), .Q(
        n8276), .QN(n3798) );
  SDFFX1 DFF_1556_Q_reg ( .D(WX10868), .SI(n8276), .SE(test_se), .CLK(CK), .Q(
        n8275), .QN(n3797) );
  SDFFX1 DFF_1557_Q_reg ( .D(WX10870), .SI(n8275), .SE(test_se), .CLK(CK), .Q(
        test_so90), .QN(n3796) );
  SDFFX1 DFF_1558_Q_reg ( .D(WX10872), .SI(test_si91), .SE(test_se), .CLK(CK), 
        .Q(n8272), .QN(n3795) );
  SDFFX1 DFF_1559_Q_reg ( .D(WX10874), .SI(n8272), .SE(test_se), .CLK(CK), .Q(
        n8271), .QN(n3794) );
  SDFFX1 DFF_1560_Q_reg ( .D(WX10876), .SI(n8271), .SE(test_se), .CLK(CK), .Q(
        n8270), .QN(n3793) );
  SDFFX1 DFF_1561_Q_reg ( .D(WX10878), .SI(n8270), .SE(test_se), .CLK(CK), .Q(
        n8269), .QN(n3792) );
  SDFFX1 DFF_1562_Q_reg ( .D(WX10880), .SI(n8269), .SE(test_se), .CLK(CK), .Q(
        n8268), .QN(n3791) );
  SDFFX1 DFF_1563_Q_reg ( .D(WX10882), .SI(n8268), .SE(test_se), .CLK(CK), .Q(
        n8267), .QN(n3790) );
  SDFFX1 DFF_1564_Q_reg ( .D(WX10884), .SI(n8267), .SE(test_se), .CLK(CK), .Q(
        n8266), .QN(n3789) );
  SDFFX1 DFF_1565_Q_reg ( .D(WX10886), .SI(n8266), .SE(test_se), .CLK(CK), .Q(
        n8265), .QN(n3788) );
  SDFFX1 DFF_1566_Q_reg ( .D(WX10888), .SI(n8265), .SE(test_se), .CLK(CK), .Q(
        n8264), .QN(n3787) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(test_se), .CLK(CK), .Q(
        n8263), .QN(n3786) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(test_se), .CLK(CK), .Q(
        n8262), .QN(n3338) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(test_se), .CLK(CK), .Q(
        n8261), .QN(n3360) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(test_se), .CLK(CK), .Q(
        n8260), .QN(n3359) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(test_se), .CLK(CK), .Q(
        n8259), .QN(n3358) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(test_se), .CLK(CK), .Q(
        n8258), .QN(n3357) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(test_se), .CLK(CK), .Q(
        n8257), .QN(n3356) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(test_se), .CLK(CK), .Q(
        test_so91), .QN(n3355) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(test_se), .CLK(CK), 
        .Q(n8254), .QN(n3354) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(test_se), .CLK(CK), .Q(
        n8253), .QN(n3353) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(test_se), .CLK(CK), .Q(
        n8252), .QN(n3352) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(test_se), .CLK(CK), .Q(
        n8251), .QN(n3351) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(test_se), .CLK(CK), .Q(
        n8250), .QN(n3350) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(test_se), .CLK(CK), .Q(
        n8249), .QN(n3349) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(test_se), .CLK(CK), .Q(
        n8248), .QN(n3348) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(test_se), .CLK(CK), .Q(
        n8247), .QN(n3347) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(test_se), .CLK(CK), .Q(
        n8246), .QN(n3346) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(test_se), .CLK(CK), .Q(
        WX11021), .QN() );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(test_se), .CLK(CK), 
        .Q(WX11023), .QN() );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(test_se), .CLK(CK), 
        .Q(WX11025), .QN() );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(test_se), .CLK(CK), 
        .Q(WX11027), .QN() );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(test_se), .CLK(CK), 
        .Q(WX11029), .QN() );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(test_se), .CLK(CK), 
        .Q(WX11031), .QN() );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(test_se), .CLK(CK), 
        .Q(WX11033), .QN() );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(test_se), .CLK(CK), 
        .Q(test_so92), .QN() );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(test_se), .CLK(CK), 
        .Q(WX11037), .QN() );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(test_se), .CLK(CK), 
        .Q(WX11039), .QN() );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(test_se), .CLK(CK), 
        .Q(WX11041), .QN() );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(test_se), .CLK(CK), 
        .Q(WX11043), .QN() );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(test_se), .CLK(CK), 
        .Q(WX11045), .QN() );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(test_se), .CLK(CK), 
        .Q(WX11047), .QN() );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(test_se), .CLK(CK), 
        .Q(WX11049), .QN() );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(test_se), .CLK(CK), 
        .Q(WX11051), .QN() );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(test_se), .CLK(CK), 
        .Q(WX11053), .QN() );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(test_se), .CLK(CK), 
        .Q(WX11055), .QN() );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(test_se), .CLK(CK), 
        .Q(WX11057), .QN() );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(test_se), .CLK(CK), 
        .Q(WX11059), .QN() );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(test_se), .CLK(CK), 
        .Q(WX11061), .QN() );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(test_se), .CLK(CK), 
        .Q(WX11063), .QN() );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(test_se), .CLK(CK), 
        .Q(WX11065), .QN() );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(test_se), .CLK(CK), 
        .Q(WX11067), .QN() );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(test_se), .CLK(CK), 
        .Q(test_so93), .QN() );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(test_se), .CLK(CK), 
        .Q(WX11071), .QN() );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(test_se), .CLK(CK), 
        .Q(WX11073), .QN() );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(test_se), .CLK(CK), 
        .Q(WX11075), .QN() );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(test_se), .CLK(CK), 
        .Q(WX11077), .QN() );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(test_se), .CLK(CK), 
        .Q(WX11079), .QN() );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(test_se), .CLK(CK), 
        .Q(WX11081), .QN() );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(test_se), .CLK(CK), 
        .Q(WX11083), .QN() );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(test_se), .CLK(CK), 
        .Q(WX11085), .QN(n3561) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(test_se), .CLK(CK), 
        .Q(WX11087), .QN(n3559) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(test_se), .CLK(CK), 
        .Q(WX11089), .QN(n3557) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(test_se), .CLK(CK), 
        .Q(WX11091), .QN(n3555) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(test_se), .CLK(CK), 
        .Q(WX11093), .QN(n3553) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(test_se), .CLK(CK), 
        .Q(WX11095), .QN(n3551) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(test_se), .CLK(CK), 
        .Q(WX11097), .QN(n3549) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(test_se), .CLK(CK), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(test_se), .CLK(CK), 
        .Q(WX11101), .QN(n3545) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(test_se), .CLK(CK), 
        .Q(test_so94), .QN(n3543) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(test_se), .CLK(CK), 
        .Q(WX11105), .QN(n3541) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(test_se), .CLK(CK), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(test_se), .CLK(CK), 
        .Q(WX11109), .QN(n3537) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(test_se), .CLK(CK), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(test_se), .CLK(CK), 
        .Q(WX11113), .QN(n3533) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(test_se), .CLK(CK), 
        .Q(WX11115), .QN(n3531) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(test_se), .CLK(CK), 
        .Q(WX11117), .QN() );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(test_se), .CLK(CK), 
        .Q(WX11119), .QN() );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(test_se), .CLK(CK), 
        .Q(WX11121), .QN() );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(test_se), .CLK(CK), 
        .Q(WX11123), .QN() );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(test_se), .CLK(CK), 
        .Q(WX11125), .QN() );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(test_se), .CLK(CK), 
        .Q(WX11127), .QN() );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(test_se), .CLK(CK), 
        .Q(WX11129), .QN() );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(test_se), .CLK(CK), 
        .Q(WX11131), .QN() );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(test_se), .CLK(CK), 
        .Q(WX11133), .QN() );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(test_se), .CLK(CK), 
        .Q(WX11135), .QN() );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(test_se), .CLK(CK), 
        .Q(test_so95), .QN() );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(test_se), .CLK(CK), 
        .Q(WX11139), .QN() );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(test_se), .CLK(CK), 
        .Q(WX11141), .QN() );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(test_se), .CLK(CK), 
        .Q(WX11143), .QN() );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(test_se), .CLK(CK), 
        .Q(WX11145), .QN() );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(test_se), .CLK(CK), 
        .Q(WX11147), .QN() );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(test_se), .CLK(CK), 
        .Q(WX11149), .QN() );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(test_se), .CLK(CK), 
        .Q(WX11151), .QN() );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(test_se), .CLK(CK), 
        .Q(WX11153), .QN() );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(test_se), .CLK(CK), 
        .Q(WX11155), .QN() );

  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155_Tj_Payload), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11157), .QN() );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11159), .QN() );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11161), .QN() );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11163), .QN() );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11165), .QN() );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11167), .QN() );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(test_se_Trojan), .CLK(CK), 
        .Q(WX11169), .QN() );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(test_se_Trojan), .CLK(CK), 
        .Q(test_so96), .QN() );


  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(test_se), .CLK(CK), 
        .Q(WX11173), .QN() );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(test_se), .CLK(CK), 
        .Q(WX11175), .QN() );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(test_se), .CLK(CK), 
        .Q(WX11177), .QN() );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(test_se), .CLK(CK), 
        .Q(WX11179), .QN() );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(test_se), .CLK(CK), 
        .Q(WX11181), .QN() );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(test_se), .CLK(CK), 
        .Q(WX11183), .QN() );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(test_se), .CLK(CK), 
        .Q(WX11185), .QN() );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(test_se), .CLK(CK), 
        .Q(WX11187), .QN() );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(test_se), .CLK(CK), 
        .Q(WX11189), .QN() );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(test_se), .CLK(CK), 
        .Q(WX11191), .QN() );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(test_se), .CLK(CK), 
        .Q(WX11193), .QN() );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(test_se), .CLK(CK), 
        .Q(WX11195), .QN() );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(test_se), .CLK(CK), 
        .Q(WX11197), .QN() );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(test_se), .CLK(CK), 
        .Q(WX11199), .QN() );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(test_se), .CLK(CK), 
        .Q(WX11201), .QN() );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(test_se), .CLK(CK), 
        .Q(WX11203), .QN() );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(test_se), .CLK(CK), 
        .Q(test_so97), .QN() );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(test_se), .CLK(CK), 
        .Q(WX11207), .QN() );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(test_se), .CLK(CK), 
        .Q(WX11209), .QN() );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(test_se), .CLK(CK), 
        .Q(WX11211), .QN() );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(test_se), .CLK(CK), 
        .Q(WX11213), .QN() );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(test_se), .CLK(CK), 
        .Q(WX11215), .QN() );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(test_se), .CLK(CK), 
        .Q(WX11217), .QN() );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(test_se), .CLK(CK), 
        .Q(WX11219), .QN() );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(test_se), .CLK(CK), 
        .Q(WX11221), .QN() );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(test_se), .CLK(CK), 
        .Q(WX11223), .QN() );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(test_se), .CLK(CK), 
        .Q(WX11225), .QN() );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(test_se), .CLK(CK), 
        .Q(WX11227), .QN() );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(test_se), .CLK(CK), 
        .Q(WX11229), .QN() );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(test_se), .CLK(CK), 
        .Q(WX11231), .QN() );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(test_se), .CLK(CK), 
        .Q(WX11233), .QN() );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(test_se), .CLK(CK), 
        .Q(WX11235), .QN() );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(test_se), .CLK(CK), 
        .Q(WX11237), .QN() );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(test_se), .CLK(CK), 
        .Q(test_so98), .QN() );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(test_se), .CLK(CK), 
        .Q(WX11241), .QN() );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(test_se), .CLK(CK), 
        .Q(WX11243), .QN() );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(test_se), .CLK(CK), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_14), .QN(DFF_1710_n1) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(test_se), .CLK(CK), 
        .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(test_se), .CLK(
        CK), .Q(CRC_OUT_1_31), .QN(DFF_1727_n1) );
  NBUFFX2 U3370 ( .IN(n4117), .Q(n4040) );
  NBUFFX2 U3371 ( .IN(n4117), .Q(n4041) );
  NBUFFX2 U3372 ( .IN(n4118), .Q(n4038) );
  NBUFFX2 U3373 ( .IN(n4118), .Q(n4039) );
  NBUFFX2 U3374 ( .IN(n4105), .Q(n4064) );
  NBUFFX2 U3375 ( .IN(n4105), .Q(n4065) );
  NBUFFX2 U3376 ( .IN(n4104), .Q(n4066) );
  NBUFFX2 U3377 ( .IN(n4104), .Q(n4067) );
  NBUFFX2 U3378 ( .IN(n4103), .Q(n4068) );
  NBUFFX2 U3379 ( .IN(n4103), .Q(n4069) );
  NBUFFX2 U3380 ( .IN(n4102), .Q(n4070) );
  NBUFFX2 U3381 ( .IN(n4102), .Q(n4071) );
  NBUFFX2 U3382 ( .IN(n4101), .Q(n4072) );
  NBUFFX2 U3383 ( .IN(n4101), .Q(n4073) );
  NBUFFX2 U3384 ( .IN(n4100), .Q(n4074) );
  NBUFFX2 U3385 ( .IN(n4100), .Q(n4075) );
  NBUFFX2 U3386 ( .IN(n4099), .Q(n4076) );
  NBUFFX2 U3387 ( .IN(n4099), .Q(n4077) );
  NBUFFX2 U3388 ( .IN(n4098), .Q(n4078) );
  NBUFFX2 U3389 ( .IN(n4098), .Q(n4079) );
  NBUFFX2 U3390 ( .IN(n4097), .Q(n4080) );
  NBUFFX2 U3391 ( .IN(n4093), .Q(n4088) );
  NBUFFX2 U3392 ( .IN(n4093), .Q(n4089) );
  NBUFFX2 U3393 ( .IN(n4116), .Q(n4042) );
  NBUFFX2 U3394 ( .IN(n4116), .Q(n4043) );
  NBUFFX2 U3395 ( .IN(n4115), .Q(n4044) );
  NBUFFX2 U3396 ( .IN(n4115), .Q(n4045) );
  NBUFFX2 U3397 ( .IN(n4114), .Q(n4046) );
  NBUFFX2 U3398 ( .IN(n4114), .Q(n4047) );
  NBUFFX2 U3399 ( .IN(n4113), .Q(n4048) );
  NBUFFX2 U3400 ( .IN(n4113), .Q(n4049) );
  NBUFFX2 U3401 ( .IN(n4112), .Q(n4050) );
  NBUFFX2 U3402 ( .IN(n4112), .Q(n4051) );
  NBUFFX2 U3403 ( .IN(n4111), .Q(n4052) );
  NBUFFX2 U3404 ( .IN(n4111), .Q(n4053) );
  NBUFFX2 U3405 ( .IN(n4110), .Q(n4054) );
  NBUFFX2 U3406 ( .IN(n4110), .Q(n4055) );
  NBUFFX2 U3407 ( .IN(n4109), .Q(n4056) );
  NBUFFX2 U3408 ( .IN(n4109), .Q(n4057) );
  NBUFFX2 U3409 ( .IN(n4108), .Q(n4058) );
  NBUFFX2 U3410 ( .IN(n4108), .Q(n4059) );
  NBUFFX2 U3411 ( .IN(n4107), .Q(n4060) );
  NBUFFX2 U3412 ( .IN(n4107), .Q(n4061) );
  NBUFFX2 U3413 ( .IN(n4106), .Q(n4062) );
  NBUFFX2 U3414 ( .IN(n4106), .Q(n4063) );
  NBUFFX2 U3415 ( .IN(n4097), .Q(n4081) );
  NBUFFX2 U3416 ( .IN(n4096), .Q(n4082) );
  NBUFFX2 U3417 ( .IN(n4096), .Q(n4083) );
  NBUFFX2 U3418 ( .IN(n4095), .Q(n4084) );
  NBUFFX2 U3419 ( .IN(n4095), .Q(n4085) );
  NBUFFX2 U3420 ( .IN(n4094), .Q(n4086) );
  NBUFFX2 U3421 ( .IN(n4094), .Q(n4087) );
  NBUFFX2 U3422 ( .IN(n4237), .Q(n4172) );
  NBUFFX2 U3423 ( .IN(n4237), .Q(n4173) );
  NBUFFX2 U3424 ( .IN(n4236), .Q(n4174) );
  NBUFFX2 U3425 ( .IN(n4236), .Q(n4175) );
  NBUFFX2 U3426 ( .IN(n4235), .Q(n4176) );
  NBUFFX2 U3427 ( .IN(n4235), .Q(n4177) );
  NBUFFX2 U3428 ( .IN(n4234), .Q(n4178) );
  NBUFFX2 U3429 ( .IN(n4233), .Q(n4180) );
  NBUFFX2 U3430 ( .IN(n4233), .Q(n4181) );
  NBUFFX2 U3431 ( .IN(n4232), .Q(n4182) );
  NBUFFX2 U3432 ( .IN(n4232), .Q(n4183) );
  NBUFFX2 U3433 ( .IN(n4231), .Q(n4184) );
  NBUFFX2 U3434 ( .IN(n4231), .Q(n4185) );
  NBUFFX2 U3435 ( .IN(n4230), .Q(n4186) );
  NBUFFX2 U3436 ( .IN(n4230), .Q(n4187) );
  NBUFFX2 U3437 ( .IN(n4229), .Q(n4188) );
  NBUFFX2 U3438 ( .IN(n4229), .Q(n4189) );
  NBUFFX2 U3439 ( .IN(n4228), .Q(n4190) );
  NBUFFX2 U3440 ( .IN(n4228), .Q(n4191) );
  NBUFFX2 U3441 ( .IN(n4227), .Q(n4192) );
  NBUFFX2 U3442 ( .IN(n4227), .Q(n4193) );
  NBUFFX2 U3443 ( .IN(n4226), .Q(n4194) );
  NBUFFX2 U3444 ( .IN(n4226), .Q(n4195) );
  NBUFFX2 U3445 ( .IN(n4225), .Q(n4196) );
  NBUFFX2 U3446 ( .IN(n4224), .Q(n4198) );
  NBUFFX2 U3447 ( .IN(n4225), .Q(n4197) );
  NBUFFX2 U3448 ( .IN(n4224), .Q(n4199) );
  NBUFFX2 U3449 ( .IN(n4223), .Q(n4200) );
  NBUFFX2 U3450 ( .IN(n4251), .Q(n4144) );
  NBUFFX2 U3451 ( .IN(n4251), .Q(n4145) );
  NBUFFX2 U3452 ( .IN(n4250), .Q(n4146) );
  NBUFFX2 U3453 ( .IN(n4250), .Q(n4147) );
  NBUFFX2 U3454 ( .IN(n4249), .Q(n4148) );
  NBUFFX2 U3455 ( .IN(n4249), .Q(n4149) );
  NBUFFX2 U3456 ( .IN(n4248), .Q(n4150) );
  NBUFFX2 U3457 ( .IN(n4248), .Q(n4151) );
  NBUFFX2 U3458 ( .IN(n4247), .Q(n4152) );
  NBUFFX2 U3459 ( .IN(n4247), .Q(n4153) );
  NBUFFX2 U3460 ( .IN(n4246), .Q(n4154) );
  NBUFFX2 U3461 ( .IN(n4246), .Q(n4155) );
  NBUFFX2 U3462 ( .IN(n4245), .Q(n4156) );
  NBUFFX2 U3463 ( .IN(n4245), .Q(n4157) );
  NBUFFX2 U3464 ( .IN(n4244), .Q(n4158) );
  NBUFFX2 U3465 ( .IN(n4244), .Q(n4159) );
  NBUFFX2 U3466 ( .IN(n4243), .Q(n4160) );
  NBUFFX2 U3467 ( .IN(n4243), .Q(n4161) );
  NBUFFX2 U3468 ( .IN(n4234), .Q(n4179) );
  NBUFFX2 U3469 ( .IN(n4242), .Q(n4162) );
  NBUFFX2 U3470 ( .IN(n4242), .Q(n4163) );
  NBUFFX2 U3471 ( .IN(n4241), .Q(n4164) );
  NBUFFX2 U3472 ( .IN(n4241), .Q(n4165) );
  NBUFFX2 U3473 ( .IN(n4240), .Q(n4166) );
  NBUFFX2 U3474 ( .IN(n4240), .Q(n4167) );
  NBUFFX2 U3475 ( .IN(n4239), .Q(n4168) );
  NBUFFX2 U3476 ( .IN(n4239), .Q(n4169) );
  NBUFFX2 U3477 ( .IN(n4238), .Q(n4170) );
  NBUFFX2 U3478 ( .IN(n4238), .Q(n4171) );
  NBUFFX2 U3479 ( .IN(n4223), .Q(n4201) );
  NBUFFX2 U3480 ( .IN(n4222), .Q(n4203) );
  NBUFFX2 U3481 ( .IN(n4222), .Q(n4202) );
  NBUFFX2 U3482 ( .IN(n4221), .Q(n4204) );
  NBUFFX2 U3483 ( .IN(n4220), .Q(n4207) );
  NBUFFX2 U3484 ( .IN(n4220), .Q(n4206) );
  NBUFFX2 U3485 ( .IN(n4221), .Q(n4205) );
  NBUFFX2 U3486 ( .IN(n4120), .Q(n4034) );
  NBUFFX2 U3487 ( .IN(n4120), .Q(n4035) );
  NBUFFX2 U3488 ( .IN(n4119), .Q(n4036) );
  NBUFFX2 U3489 ( .IN(n4119), .Q(n4037) );
  NBUFFX2 U3490 ( .IN(n4092), .Q(n4090) );
  NBUFFX2 U3491 ( .IN(n4217), .Q(n4212) );
  NBUFFX2 U3492 ( .IN(n4218), .Q(n4211) );
  NBUFFX2 U3493 ( .IN(n4219), .Q(n4209) );
  NBUFFX2 U3494 ( .IN(n4219), .Q(n4208) );
  NBUFFX2 U3495 ( .IN(n4218), .Q(n4210) );
  NBUFFX2 U3496 ( .IN(n4217), .Q(n4213) );
  NBUFFX2 U3497 ( .IN(n4216), .Q(n4214) );
  NBUFFX2 U3498 ( .IN(n4216), .Q(n4215) );
  NBUFFX2 U3499 ( .IN(n4092), .Q(n4091) );
  NBUFFX2 U3500 ( .IN(n4259), .Q(n4237) );
  NBUFFX2 U3501 ( .IN(n4259), .Q(n4236) );
  NBUFFX2 U3502 ( .IN(n4122), .Q(n4117) );
  NBUFFX2 U3503 ( .IN(n4260), .Q(n4235) );
  NBUFFX2 U3504 ( .IN(n4122), .Q(n4118) );
  NBUFFX2 U3505 ( .IN(n4261), .Q(n4233) );
  NBUFFX2 U3506 ( .IN(n4128), .Q(n4105) );
  NBUFFX2 U3507 ( .IN(n4261), .Q(n4232) );
  NBUFFX2 U3508 ( .IN(n4129), .Q(n4104) );
  NBUFFX2 U3509 ( .IN(n4262), .Q(n4231) );
  NBUFFX2 U3510 ( .IN(n4129), .Q(n4103) );
  NBUFFX2 U3511 ( .IN(n4262), .Q(n4230) );
  NBUFFX2 U3512 ( .IN(n4263), .Q(n4229) );
  NBUFFX2 U3513 ( .IN(n4130), .Q(n4102) );
  NBUFFX2 U3514 ( .IN(n4263), .Q(n4228) );
  NBUFFX2 U3515 ( .IN(n4130), .Q(n4101) );
  NBUFFX2 U3516 ( .IN(n4264), .Q(n4227) );
  NBUFFX2 U3517 ( .IN(n4131), .Q(n4100) );
  NBUFFX2 U3518 ( .IN(n4264), .Q(n4226) );
  NBUFFX2 U3519 ( .IN(n4131), .Q(n4099) );
  NBUFFX2 U3520 ( .IN(n4265), .Q(n4225) );
  NBUFFX2 U3521 ( .IN(n4265), .Q(n4224) );
  NBUFFX2 U3522 ( .IN(n4132), .Q(n4098) );
  NBUFFX2 U3523 ( .IN(n4134), .Q(n4093) );
  NBUFFX2 U3524 ( .IN(n4252), .Q(n4251) );
  NBUFFX2 U3525 ( .IN(n4252), .Q(n4250) );
  NBUFFX2 U3526 ( .IN(n4123), .Q(n4116) );
  NBUFFX2 U3527 ( .IN(n4253), .Q(n4249) );
  NBUFFX2 U3528 ( .IN(n4123), .Q(n4115) );
  NBUFFX2 U3529 ( .IN(n4253), .Q(n4248) );
  NBUFFX2 U3530 ( .IN(n4124), .Q(n4114) );
  NBUFFX2 U3531 ( .IN(n4254), .Q(n4247) );
  NBUFFX2 U3532 ( .IN(n4124), .Q(n4113) );
  NBUFFX2 U3533 ( .IN(n4254), .Q(n4246) );
  NBUFFX2 U3534 ( .IN(n4125), .Q(n4112) );
  NBUFFX2 U3535 ( .IN(n4255), .Q(n4245) );
  NBUFFX2 U3536 ( .IN(n4125), .Q(n4111) );
  NBUFFX2 U3537 ( .IN(n4255), .Q(n4244) );
  NBUFFX2 U3538 ( .IN(n4256), .Q(n4243) );
  NBUFFX2 U3539 ( .IN(n4260), .Q(n4234) );
  NBUFFX2 U3540 ( .IN(n4126), .Q(n4110) );
  NBUFFX2 U3541 ( .IN(n4256), .Q(n4242) );
  NBUFFX2 U3542 ( .IN(n4126), .Q(n4109) );
  NBUFFX2 U3543 ( .IN(n4257), .Q(n4241) );
  NBUFFX2 U3544 ( .IN(n4127), .Q(n4108) );
  NBUFFX2 U3545 ( .IN(n4257), .Q(n4240) );
  NBUFFX2 U3546 ( .IN(n4258), .Q(n4239) );
  NBUFFX2 U3547 ( .IN(n4127), .Q(n4107) );
  NBUFFX2 U3548 ( .IN(n4258), .Q(n4238) );
  NBUFFX2 U3549 ( .IN(n4128), .Q(n4106) );
  NBUFFX2 U3550 ( .IN(n4266), .Q(n4223) );
  NBUFFX2 U3551 ( .IN(n4132), .Q(n4097) );
  NBUFFX2 U3552 ( .IN(n4266), .Q(n4222) );
  NBUFFX2 U3553 ( .IN(n4133), .Q(n4096) );
  NBUFFX2 U3554 ( .IN(n4133), .Q(n4095) );
  NBUFFX2 U3555 ( .IN(n4267), .Q(n4220) );
  NBUFFX2 U3556 ( .IN(n4267), .Q(n4221) );
  NBUFFX2 U3557 ( .IN(n4134), .Q(n4094) );
  ISOLANDX1 U3558 ( .D(n4479), .ISO(n4586), .Q(n2245) );
  NBUFFX2 U3559 ( .IN(n4482), .Q(n4474) );
  NBUFFX2 U3560 ( .IN(n4482), .Q(n4475) );
  NBUFFX2 U3561 ( .IN(n4481), .Q(n4476) );
  NBUFFX2 U3562 ( .IN(n4481), .Q(n4477) );
  NBUFFX2 U3563 ( .IN(n4480), .Q(n4478) );
  NBUFFX2 U3564 ( .IN(n4507), .Q(n4424) );
  NBUFFX2 U3565 ( .IN(n4507), .Q(n4425) );
  NBUFFX2 U3566 ( .IN(n4506), .Q(n4426) );
  NBUFFX2 U3567 ( .IN(n4506), .Q(n4427) );
  NBUFFX2 U3568 ( .IN(n4505), .Q(n4428) );
  NBUFFX2 U3569 ( .IN(n4505), .Q(n4429) );
  NBUFFX2 U3570 ( .IN(n4504), .Q(n4430) );
  NBUFFX2 U3571 ( .IN(n4504), .Q(n4431) );
  NBUFFX2 U3572 ( .IN(n4503), .Q(n4432) );
  NBUFFX2 U3573 ( .IN(n4503), .Q(n4433) );
  NBUFFX2 U3574 ( .IN(n4502), .Q(n4434) );
  NBUFFX2 U3575 ( .IN(n4502), .Q(n4435) );
  NBUFFX2 U3576 ( .IN(n4501), .Q(n4436) );
  NBUFFX2 U3577 ( .IN(n4501), .Q(n4437) );
  NBUFFX2 U3578 ( .IN(n4500), .Q(n4438) );
  NBUFFX2 U3579 ( .IN(n4500), .Q(n4439) );
  NBUFFX2 U3580 ( .IN(n4499), .Q(n4440) );
  NBUFFX2 U3581 ( .IN(n4499), .Q(n4441) );
  NBUFFX2 U3582 ( .IN(n4495), .Q(n4449) );
  NBUFFX2 U3583 ( .IN(n4494), .Q(n4450) );
  NBUFFX2 U3584 ( .IN(n4494), .Q(n4451) );
  NBUFFX2 U3585 ( .IN(n4493), .Q(n4452) );
  NBUFFX2 U3586 ( .IN(n4493), .Q(n4453) );
  NBUFFX2 U3587 ( .IN(n4492), .Q(n4454) );
  NBUFFX2 U3588 ( .IN(n4492), .Q(n4455) );
  NBUFFX2 U3589 ( .IN(n4491), .Q(n4456) );
  NBUFFX2 U3590 ( .IN(n4491), .Q(n4457) );
  NBUFFX2 U3591 ( .IN(n4490), .Q(n4458) );
  NBUFFX2 U3592 ( .IN(n4490), .Q(n4459) );
  NBUFFX2 U3593 ( .IN(n4489), .Q(n4460) );
  NBUFFX2 U3594 ( .IN(n4489), .Q(n4461) );
  NBUFFX2 U3595 ( .IN(n4488), .Q(n4462) );
  NBUFFX2 U3596 ( .IN(n4488), .Q(n4463) );
  NBUFFX2 U3597 ( .IN(n4487), .Q(n4464) );
  NBUFFX2 U3598 ( .IN(n4487), .Q(n4465) );
  NBUFFX2 U3599 ( .IN(n4486), .Q(n4466) );
  NBUFFX2 U3600 ( .IN(n4486), .Q(n4467) );
  NBUFFX2 U3601 ( .IN(n4485), .Q(n4468) );
  NBUFFX2 U3602 ( .IN(n4485), .Q(n4469) );
  NBUFFX2 U3603 ( .IN(n4484), .Q(n4470) );
  NBUFFX2 U3604 ( .IN(n4484), .Q(n4471) );
  NBUFFX2 U3605 ( .IN(n4483), .Q(n4472) );
  NBUFFX2 U3606 ( .IN(n4483), .Q(n4473) );
  NBUFFX2 U3607 ( .IN(n4498), .Q(n4442) );
  NBUFFX2 U3608 ( .IN(n4498), .Q(n4443) );
  NBUFFX2 U3609 ( .IN(n4497), .Q(n4444) );
  NBUFFX2 U3610 ( .IN(n4497), .Q(n4445) );
  NBUFFX2 U3611 ( .IN(n4496), .Q(n4446) );
  NBUFFX2 U3612 ( .IN(n4496), .Q(n4447) );
  NBUFFX2 U3613 ( .IN(n4495), .Q(n4448) );
  NBUFFX2 U3614 ( .IN(n4480), .Q(n4479) );
  NBUFFX2 U3615 ( .IN(n4275), .Q(n4259) );
  NBUFFX2 U3616 ( .IN(n4142), .Q(n4122) );
  NBUFFX2 U3617 ( .IN(n4274), .Q(n4261) );
  NBUFFX2 U3618 ( .IN(n4139), .Q(n4129) );
  NBUFFX2 U3619 ( .IN(n4273), .Q(n4262) );
  NBUFFX2 U3620 ( .IN(n4273), .Q(n4263) );
  NBUFFX2 U3621 ( .IN(n4138), .Q(n4130) );
  NBUFFX2 U3622 ( .IN(n4272), .Q(n4264) );
  NBUFFX2 U3623 ( .IN(n4138), .Q(n4131) );
  NBUFFX2 U3624 ( .IN(n4272), .Q(n4265) );
  NBUFFX2 U3625 ( .IN(n4278), .Q(n4252) );
  NBUFFX2 U3626 ( .IN(n4142), .Q(n4123) );
  NBUFFX2 U3627 ( .IN(n4278), .Q(n4253) );
  NBUFFX2 U3628 ( .IN(n4141), .Q(n4124) );
  NBUFFX2 U3629 ( .IN(n4277), .Q(n4254) );
  NBUFFX2 U3630 ( .IN(n4141), .Q(n4125) );
  NBUFFX2 U3631 ( .IN(n4277), .Q(n4255) );
  NBUFFX2 U3632 ( .IN(n4274), .Q(n4260) );
  NBUFFX2 U3633 ( .IN(n4276), .Q(n4256) );
  NBUFFX2 U3634 ( .IN(n4140), .Q(n4126) );
  NBUFFX2 U3635 ( .IN(n4276), .Q(n4257) );
  NBUFFX2 U3636 ( .IN(n4140), .Q(n4127) );
  NBUFFX2 U3637 ( .IN(n4275), .Q(n4258) );
  NBUFFX2 U3638 ( .IN(n4139), .Q(n4128) );
  NBUFFX2 U3639 ( .IN(n4137), .Q(n4132) );
  NBUFFX2 U3640 ( .IN(n4271), .Q(n4266) );
  NBUFFX2 U3641 ( .IN(n4137), .Q(n4133) );
  NBUFFX2 U3642 ( .IN(n4271), .Q(n4267) );
  NBUFFX2 U3643 ( .IN(n4136), .Q(n4134) );
  NBUFFX2 U3644 ( .IN(n4121), .Q(n4119) );
  NBUFFX2 U3645 ( .IN(n4121), .Q(n4120) );
  NBUFFX2 U3646 ( .IN(n4269), .Q(n4217) );
  NBUFFX2 U3647 ( .IN(n4135), .Q(n4092) );
  NBUFFX2 U3648 ( .IN(n4136), .Q(n4135) );
  NBUFFX2 U3649 ( .IN(n4268), .Q(n4219) );
  NBUFFX2 U3650 ( .IN(n4268), .Q(n4218) );
  NBUFFX2 U3651 ( .IN(n4269), .Q(n4216) );
  NBUFFX2 U3652 ( .IN(n4679), .Q(n4558) );
  NBUFFX2 U3653 ( .IN(n4377), .Q(n4312) );
  NBUFFX2 U3654 ( .IN(n4377), .Q(n4313) );
  NBUFFX2 U3655 ( .IN(n4376), .Q(n4314) );
  NBUFFX2 U3656 ( .IN(n4376), .Q(n4315) );
  NBUFFX2 U3657 ( .IN(n4375), .Q(n4316) );
  NBUFFX2 U3658 ( .IN(n4375), .Q(n4317) );
  NBUFFX2 U3659 ( .IN(n4374), .Q(n4318) );
  NBUFFX2 U3660 ( .IN(n4373), .Q(n4320) );
  NBUFFX2 U3661 ( .IN(n4373), .Q(n4321) );
  NBUFFX2 U3662 ( .IN(n4372), .Q(n4322) );
  NBUFFX2 U3663 ( .IN(n4372), .Q(n4323) );
  NBUFFX2 U3664 ( .IN(n4371), .Q(n4324) );
  NBUFFX2 U3665 ( .IN(n4371), .Q(n4325) );
  NBUFFX2 U3666 ( .IN(n4370), .Q(n4326) );
  NBUFFX2 U3667 ( .IN(n4370), .Q(n4327) );
  NBUFFX2 U3668 ( .IN(n4369), .Q(n4328) );
  NBUFFX2 U3669 ( .IN(n4369), .Q(n4329) );
  NBUFFX2 U3670 ( .IN(n4368), .Q(n4330) );
  NBUFFX2 U3671 ( .IN(n4368), .Q(n4331) );
  NBUFFX2 U3672 ( .IN(n4367), .Q(n4332) );
  NBUFFX2 U3673 ( .IN(n4367), .Q(n4333) );
  NBUFFX2 U3674 ( .IN(n4366), .Q(n4334) );
  NBUFFX2 U3675 ( .IN(n4366), .Q(n4335) );
  NBUFFX2 U3676 ( .IN(n4365), .Q(n4336) );
  NBUFFX2 U3677 ( .IN(n4364), .Q(n4338) );
  NBUFFX2 U3678 ( .IN(n4365), .Q(n4337) );
  NBUFFX2 U3679 ( .IN(n4364), .Q(n4339) );
  NBUFFX2 U3680 ( .IN(n4363), .Q(n4340) );
  NBUFFX2 U3681 ( .IN(n4391), .Q(n4284) );
  NBUFFX2 U3682 ( .IN(n4391), .Q(n4285) );
  NBUFFX2 U3683 ( .IN(n4390), .Q(n4286) );
  NBUFFX2 U3684 ( .IN(n4390), .Q(n4287) );
  NBUFFX2 U3685 ( .IN(n4389), .Q(n4288) );
  NBUFFX2 U3686 ( .IN(n4389), .Q(n4289) );
  NBUFFX2 U3687 ( .IN(n4388), .Q(n4290) );
  NBUFFX2 U3688 ( .IN(n4388), .Q(n4291) );
  NBUFFX2 U3689 ( .IN(n4387), .Q(n4292) );
  NBUFFX2 U3690 ( .IN(n4387), .Q(n4293) );
  NBUFFX2 U3691 ( .IN(n4386), .Q(n4294) );
  NBUFFX2 U3692 ( .IN(n4386), .Q(n4295) );
  NBUFFX2 U3693 ( .IN(n4385), .Q(n4296) );
  NBUFFX2 U3694 ( .IN(n4385), .Q(n4297) );
  NBUFFX2 U3695 ( .IN(n4384), .Q(n4298) );
  NBUFFX2 U3696 ( .IN(n4384), .Q(n4299) );
  NBUFFX2 U3697 ( .IN(n4383), .Q(n4300) );
  NBUFFX2 U3698 ( .IN(n4383), .Q(n4301) );
  NBUFFX2 U3699 ( .IN(n4374), .Q(n4319) );
  NBUFFX2 U3700 ( .IN(n4382), .Q(n4302) );
  NBUFFX2 U3701 ( .IN(n4382), .Q(n4303) );
  NBUFFX2 U3702 ( .IN(n4381), .Q(n4304) );
  NBUFFX2 U3703 ( .IN(n4381), .Q(n4305) );
  NBUFFX2 U3704 ( .IN(n4380), .Q(n4306) );
  NBUFFX2 U3705 ( .IN(n4380), .Q(n4307) );
  NBUFFX2 U3706 ( .IN(n4379), .Q(n4308) );
  NBUFFX2 U3707 ( .IN(n4379), .Q(n4309) );
  NBUFFX2 U3708 ( .IN(n4378), .Q(n4310) );
  NBUFFX2 U3709 ( .IN(n4378), .Q(n4311) );
  NBUFFX2 U3710 ( .IN(n4363), .Q(n4341) );
  NBUFFX2 U3711 ( .IN(n4362), .Q(n4343) );
  NBUFFX2 U3712 ( .IN(n4362), .Q(n4342) );
  NBUFFX2 U3713 ( .IN(n4361), .Q(n4344) );
  NBUFFX2 U3714 ( .IN(n4360), .Q(n4347) );
  NBUFFX2 U3715 ( .IN(n4360), .Q(n4346) );
  NBUFFX2 U3716 ( .IN(n4361), .Q(n4345) );
  NBUFFX2 U3717 ( .IN(n2153), .Q(n4138) );
  NBUFFX2 U3718 ( .IN(n2153), .Q(n4142) );
  NBUFFX2 U3719 ( .IN(n2153), .Q(n4141) );
  NBUFFX2 U3720 ( .IN(n2153), .Q(n4140) );
  NBUFFX2 U3721 ( .IN(n2153), .Q(n4139) );
  NBUFFX2 U3722 ( .IN(n2153), .Q(n4137) );
  NBUFFX2 U3723 ( .IN(n2153), .Q(n4136) );
  NBUFFX2 U3724 ( .IN(n4281), .Q(n4273) );
  NBUFFX2 U3725 ( .IN(n4282), .Q(n4272) );
  NBUFFX2 U3726 ( .IN(n4279), .Q(n4278) );
  NBUFFX2 U3727 ( .IN(n4279), .Q(n4277) );
  NBUFFX2 U3728 ( .IN(n4281), .Q(n4274) );
  NBUFFX2 U3729 ( .IN(n4280), .Q(n4276) );
  NBUFFX2 U3730 ( .IN(n4280), .Q(n4275) );
  NBUFFX2 U3731 ( .IN(n4282), .Q(n4271) );
  NBUFFX2 U3732 ( .IN(n4143), .Q(n4121) );
  NBUFFX2 U3733 ( .IN(n2153), .Q(n4143) );
  NBUFFX2 U3734 ( .IN(n4270), .Q(n4268) );
  NBUFFX2 U3735 ( .IN(n4270), .Q(n4269) );
  NBUFFX2 U3736 ( .IN(n4521), .Q(n4480) );
  NBUFFX2 U3737 ( .IN(n4520), .Q(n4482) );
  NBUFFX2 U3738 ( .IN(n4521), .Q(n4481) );
  NBUFFX2 U3739 ( .IN(n4508), .Q(n4507) );
  NBUFFX2 U3740 ( .IN(n4508), .Q(n4506) );
  NBUFFX2 U3741 ( .IN(n4509), .Q(n4505) );
  NBUFFX2 U3742 ( .IN(n4509), .Q(n4504) );
  NBUFFX2 U3743 ( .IN(n4510), .Q(n4503) );
  NBUFFX2 U3744 ( .IN(n4510), .Q(n4502) );
  NBUFFX2 U3745 ( .IN(n4511), .Q(n4501) );
  NBUFFX2 U3746 ( .IN(n4511), .Q(n4500) );
  NBUFFX2 U3747 ( .IN(n4512), .Q(n4499) );
  NBUFFX2 U3748 ( .IN(n4514), .Q(n4494) );
  NBUFFX2 U3749 ( .IN(n4515), .Q(n4493) );
  NBUFFX2 U3750 ( .IN(n4515), .Q(n4492) );
  NBUFFX2 U3751 ( .IN(n4516), .Q(n4491) );
  NBUFFX2 U3752 ( .IN(n4516), .Q(n4490) );
  NBUFFX2 U3753 ( .IN(n4517), .Q(n4489) );
  NBUFFX2 U3754 ( .IN(n4517), .Q(n4488) );
  NBUFFX2 U3755 ( .IN(n4518), .Q(n4487) );
  NBUFFX2 U3756 ( .IN(n4518), .Q(n4486) );
  NBUFFX2 U3757 ( .IN(n4519), .Q(n4485) );
  NBUFFX2 U3758 ( .IN(n4519), .Q(n4484) );
  NBUFFX2 U3759 ( .IN(n4520), .Q(n4483) );
  NBUFFX2 U3760 ( .IN(n4512), .Q(n4498) );
  NBUFFX2 U3761 ( .IN(n4513), .Q(n4497) );
  NBUFFX2 U3762 ( .IN(n4513), .Q(n4496) );
  NBUFFX2 U3763 ( .IN(n4514), .Q(n4495) );
  NBUFFX2 U3764 ( .IN(n4667), .Q(n4581) );
  NBUFFX2 U3765 ( .IN(n4667), .Q(n4582) );
  NBUFFX2 U3766 ( .IN(n4666), .Q(n4583) );
  NBUFFX2 U3767 ( .IN(n4665), .Q(n4585) );
  NBUFFX2 U3768 ( .IN(n4665), .Q(n4586) );
  NBUFFX2 U3769 ( .IN(n4664), .Q(n4587) );
  NBUFFX2 U3770 ( .IN(n4654), .Q(n4608) );
  NBUFFX2 U3771 ( .IN(n4653), .Q(n4609) );
  NBUFFX2 U3772 ( .IN(n4653), .Q(n4610) );
  NBUFFX2 U3773 ( .IN(n4652), .Q(n4611) );
  NBUFFX2 U3774 ( .IN(n4652), .Q(n4612) );
  NBUFFX2 U3775 ( .IN(n4651), .Q(n4613) );
  NBUFFX2 U3776 ( .IN(n4654), .Q(n4607) );
  NBUFFX2 U3777 ( .IN(n4641), .Q(n4634) );
  NBUFFX2 U3778 ( .IN(n4640), .Q(n4635) );
  NBUFFX2 U3779 ( .IN(n4640), .Q(n4636) );
  NBUFFX2 U3780 ( .IN(n4649), .Q(n4617) );
  NBUFFX2 U3781 ( .IN(n4649), .Q(n4618) );
  NBUFFX2 U3782 ( .IN(n4648), .Q(n4619) );
  NBUFFX2 U3783 ( .IN(n4648), .Q(n4620) );
  NBUFFX2 U3784 ( .IN(n4647), .Q(n4621) );
  NBUFFX2 U3785 ( .IN(n4645), .Q(n4625) );
  NBUFFX2 U3786 ( .IN(n4645), .Q(n4626) );
  NBUFFX2 U3787 ( .IN(n4644), .Q(n4627) );
  NBUFFX2 U3788 ( .IN(n4669), .Q(n4578) );
  NBUFFX2 U3789 ( .IN(n4669), .Q(n4577) );
  NBUFFX2 U3790 ( .IN(n4670), .Q(n4576) );
  NBUFFX2 U3791 ( .IN(n4670), .Q(n4575) );
  NBUFFX2 U3792 ( .IN(n4671), .Q(n4573) );
  NBUFFX2 U3793 ( .IN(n4672), .Q(n4572) );
  NBUFFX2 U3794 ( .IN(n4671), .Q(n4574) );
  NBUFFX2 U3795 ( .IN(n4664), .Q(n4588) );
  NBUFFX2 U3796 ( .IN(n4663), .Q(n4589) );
  NBUFFX2 U3797 ( .IN(n4663), .Q(n4590) );
  NBUFFX2 U3798 ( .IN(n4662), .Q(n4591) );
  NBUFFX2 U3799 ( .IN(n4662), .Q(n4592) );
  NBUFFX2 U3800 ( .IN(n4661), .Q(n4593) );
  NBUFFX2 U3801 ( .IN(n4661), .Q(n4594) );
  NBUFFX2 U3802 ( .IN(n4660), .Q(n4595) );
  NBUFFX2 U3803 ( .IN(n4666), .Q(n4584) );
  NBUFFX2 U3804 ( .IN(n4668), .Q(n4579) );
  NBUFFX2 U3805 ( .IN(n4668), .Q(n4580) );
  NBUFFX2 U3806 ( .IN(n4651), .Q(n4614) );
  NBUFFX2 U3807 ( .IN(n4650), .Q(n4615) );
  NBUFFX2 U3808 ( .IN(n4650), .Q(n4616) );
  NBUFFX2 U3809 ( .IN(n4660), .Q(n4596) );
  NBUFFX2 U3810 ( .IN(n4659), .Q(n4597) );
  NBUFFX2 U3811 ( .IN(n4659), .Q(n4598) );
  NBUFFX2 U3812 ( .IN(n4658), .Q(n4599) );
  NBUFFX2 U3813 ( .IN(n4658), .Q(n4600) );
  NBUFFX2 U3814 ( .IN(n4657), .Q(n4601) );
  NBUFFX2 U3815 ( .IN(n4657), .Q(n4602) );
  NBUFFX2 U3816 ( .IN(n4656), .Q(n4603) );
  NBUFFX2 U3817 ( .IN(n4656), .Q(n4604) );
  NBUFFX2 U3818 ( .IN(n4655), .Q(n4605) );
  NBUFFX2 U3819 ( .IN(n4655), .Q(n4606) );
  NBUFFX2 U3820 ( .IN(n4644), .Q(n4628) );
  NBUFFX2 U3821 ( .IN(n4643), .Q(n4629) );
  NBUFFX2 U3822 ( .IN(n4643), .Q(n4630) );
  NBUFFX2 U3823 ( .IN(n4642), .Q(n4631) );
  NBUFFX2 U3824 ( .IN(n4642), .Q(n4632) );
  NBUFFX2 U3825 ( .IN(n4641), .Q(n4633) );
  NBUFFX2 U3826 ( .IN(n4647), .Q(n4622) );
  NBUFFX2 U3827 ( .IN(n4646), .Q(n4623) );
  NBUFFX2 U3828 ( .IN(n4646), .Q(n4624) );
  NBUFFX2 U3829 ( .IN(n4678), .Q(n4559) );
  NBUFFX2 U3830 ( .IN(n4677), .Q(n4561) );
  NBUFFX2 U3831 ( .IN(n4679), .Q(n4557) );
  NBUFFX2 U3832 ( .IN(n4675), .Q(n4565) );
  NBUFFX2 U3833 ( .IN(n4676), .Q(n4564) );
  NBUFFX2 U3834 ( .IN(n4680), .Q(n4556) );
  NBUFFX2 U3835 ( .IN(n4676), .Q(n4563) );
  NBUFFX2 U3836 ( .IN(n4677), .Q(n4562) );
  NBUFFX2 U3837 ( .IN(n4678), .Q(n4560) );
  NBUFFX2 U3838 ( .IN(n4674), .Q(n4568) );
  NBUFFX2 U3839 ( .IN(n4673), .Q(n4570) );
  NBUFFX2 U3840 ( .IN(n4673), .Q(n4569) );
  NBUFFX2 U3841 ( .IN(n4675), .Q(n4566) );
  NBUFFX2 U3842 ( .IN(n4674), .Q(n4567) );
  NBUFFX2 U3843 ( .IN(n4692), .Q(n4532) );
  NBUFFX2 U3844 ( .IN(n4692), .Q(n4531) );
  NBUFFX2 U3845 ( .IN(n4683), .Q(n4549) );
  NBUFFX2 U3846 ( .IN(n4683), .Q(n4550) );
  NBUFFX2 U3847 ( .IN(n4682), .Q(n4551) );
  NBUFFX2 U3848 ( .IN(n4688), .Q(n4540) );
  NBUFFX2 U3849 ( .IN(n4687), .Q(n4541) );
  NBUFFX2 U3850 ( .IN(n4684), .Q(n4547) );
  NBUFFX2 U3851 ( .IN(n4685), .Q(n4545) );
  NBUFFX2 U3852 ( .IN(n4693), .Q(n4529) );
  NBUFFX2 U3853 ( .IN(n4680), .Q(n4555) );
  NBUFFX2 U3854 ( .IN(n4682), .Q(n4552) );
  NBUFFX2 U3855 ( .IN(n4681), .Q(n4554) );
  NBUFFX2 U3856 ( .IN(n4681), .Q(n4553) );
  NBUFFX2 U3857 ( .IN(n4684), .Q(n4548) );
  NBUFFX2 U3858 ( .IN(n4693), .Q(n4530) );
  NBUFFX2 U3859 ( .IN(n4689), .Q(n4537) );
  NBUFFX2 U3860 ( .IN(n4689), .Q(n4538) );
  NBUFFX2 U3861 ( .IN(n4685), .Q(n4546) );
  NBUFFX2 U3862 ( .IN(n4686), .Q(n4544) );
  NBUFFX2 U3863 ( .IN(n4686), .Q(n4543) );
  NBUFFX2 U3864 ( .IN(n4687), .Q(n4542) );
  NBUFFX2 U3865 ( .IN(n4688), .Q(n4539) );
  NBUFFX2 U3866 ( .IN(n4690), .Q(n4535) );
  NBUFFX2 U3867 ( .IN(n4691), .Q(n4534) );
  NBUFFX2 U3868 ( .IN(n4691), .Q(n4533) );
  NBUFFX2 U3869 ( .IN(n4690), .Q(n4536) );
  NBUFFX2 U3870 ( .IN(n4672), .Q(n4571) );
  ISOLANDX1 U3871 ( .D(n3278), .ISO(n4766), .Q(n2153) );
  NOR2X0 U3872 ( .IN1(n4558), .IN2(n4743), .QN(n3278) );
  NBUFFX2 U3873 ( .IN(n4357), .Q(n4352) );
  NBUFFX2 U3874 ( .IN(n4358), .Q(n4351) );
  NBUFFX2 U3875 ( .IN(n4359), .Q(n4349) );
  NBUFFX2 U3876 ( .IN(n4359), .Q(n4348) );
  NBUFFX2 U3877 ( .IN(n4358), .Q(n4350) );
  NBUFFX2 U3878 ( .IN(n4357), .Q(n4353) );
  NBUFFX2 U3879 ( .IN(n4356), .Q(n4354) );
  NBUFFX2 U3880 ( .IN(n4356), .Q(n4355) );
  NBUFFX2 U3881 ( .IN(n4283), .Q(n4270) );
  NBUFFX2 U3882 ( .IN(n2152), .Q(n4283) );
  NBUFFX2 U3883 ( .IN(n4522), .Q(n4521) );
  NBUFFX2 U3884 ( .IN(n4528), .Q(n4508) );
  NBUFFX2 U3885 ( .IN(n4528), .Q(n4509) );
  NBUFFX2 U3886 ( .IN(n4527), .Q(n4510) );
  NBUFFX2 U3887 ( .IN(n4527), .Q(n4511) );
  NBUFFX2 U3888 ( .IN(n4525), .Q(n4515) );
  NBUFFX2 U3889 ( .IN(n4524), .Q(n4516) );
  NBUFFX2 U3890 ( .IN(n4524), .Q(n4517) );
  NBUFFX2 U3891 ( .IN(n4523), .Q(n4518) );
  NBUFFX2 U3892 ( .IN(n4523), .Q(n4519) );
  NBUFFX2 U3893 ( .IN(n4522), .Q(n4520) );
  NBUFFX2 U3894 ( .IN(n4526), .Q(n4512) );
  NBUFFX2 U3895 ( .IN(n4526), .Q(n4513) );
  NBUFFX2 U3896 ( .IN(n4525), .Q(n4514) );
  NBUFFX2 U3897 ( .IN(n4399), .Q(n4377) );
  NBUFFX2 U3898 ( .IN(n4399), .Q(n4376) );
  NBUFFX2 U3899 ( .IN(n4400), .Q(n4375) );
  NBUFFX2 U3900 ( .IN(n4401), .Q(n4373) );
  NBUFFX2 U3901 ( .IN(n4401), .Q(n4372) );
  NBUFFX2 U3902 ( .IN(n4402), .Q(n4371) );
  NBUFFX2 U3903 ( .IN(n4402), .Q(n4370) );
  NBUFFX2 U3904 ( .IN(n4403), .Q(n4369) );
  NBUFFX2 U3905 ( .IN(n4403), .Q(n4368) );
  NBUFFX2 U3906 ( .IN(n4404), .Q(n4367) );
  NBUFFX2 U3907 ( .IN(n4404), .Q(n4366) );
  NBUFFX2 U3908 ( .IN(n4405), .Q(n4365) );
  NBUFFX2 U3909 ( .IN(n4405), .Q(n4364) );
  NBUFFX2 U3910 ( .IN(n4392), .Q(n4391) );
  NBUFFX2 U3911 ( .IN(n4392), .Q(n4390) );
  NBUFFX2 U3912 ( .IN(n4393), .Q(n4389) );
  NBUFFX2 U3913 ( .IN(n4393), .Q(n4388) );
  NBUFFX2 U3914 ( .IN(n4394), .Q(n4387) );
  NBUFFX2 U3915 ( .IN(n4394), .Q(n4386) );
  NBUFFX2 U3916 ( .IN(n4701), .Q(n4679) );
  NBUFFX2 U3917 ( .IN(n4395), .Q(n4385) );
  NBUFFX2 U3918 ( .IN(n4395), .Q(n4384) );
  NBUFFX2 U3919 ( .IN(n4396), .Q(n4383) );
  NBUFFX2 U3920 ( .IN(n4400), .Q(n4374) );
  NBUFFX2 U3921 ( .IN(n4396), .Q(n4382) );
  NBUFFX2 U3922 ( .IN(n4397), .Q(n4381) );
  NBUFFX2 U3923 ( .IN(n4397), .Q(n4380) );
  NBUFFX2 U3924 ( .IN(n4398), .Q(n4379) );
  NBUFFX2 U3925 ( .IN(n4398), .Q(n4378) );
  NBUFFX2 U3926 ( .IN(n4406), .Q(n4363) );
  NBUFFX2 U3927 ( .IN(n4406), .Q(n4362) );
  NBUFFX2 U3928 ( .IN(n4407), .Q(n4360) );
  NBUFFX2 U3929 ( .IN(n4407), .Q(n4361) );
  NBUFFX2 U3930 ( .IN(n2152), .Q(n4279) );
  NBUFFX2 U3931 ( .IN(n2152), .Q(n4281) );
  NBUFFX2 U3932 ( .IN(n2152), .Q(n4280) );
  NBUFFX2 U3933 ( .IN(n2152), .Q(n4282) );
  NBUFFX2 U3934 ( .IN(n4639), .Q(n4637) );
  NBUFFX2 U3935 ( .IN(n4639), .Q(n4638) );
  NBUFFX2 U3936 ( .IN(n4694), .Q(n4692) );
  NBUFFX2 U3937 ( .IN(n4707), .Q(n4667) );
  NBUFFX2 U3938 ( .IN(n4708), .Q(n4665) );
  NBUFFX2 U3939 ( .IN(n4714), .Q(n4653) );
  NBUFFX2 U3940 ( .IN(n4714), .Q(n4652) );
  NBUFFX2 U3941 ( .IN(n4699), .Q(n4683) );
  NBUFFX2 U3942 ( .IN(n4713), .Q(n4654) );
  NBUFFX2 U3943 ( .IN(n4720), .Q(n4640) );
  NBUFFX2 U3944 ( .IN(n4716), .Q(n4649) );
  NBUFFX2 U3945 ( .IN(n4716), .Q(n4648) );
  NBUFFX2 U3946 ( .IN(n4699), .Q(n4682) );
  NBUFFX2 U3947 ( .IN(n4700), .Q(n4681) );
  NBUFFX2 U3948 ( .IN(n4718), .Q(n4645) );
  NBUFFX2 U3949 ( .IN(n4698), .Q(n4684) );
  NBUFFX2 U3950 ( .IN(n4694), .Q(n4693) );
  NBUFFX2 U3951 ( .IN(n4696), .Q(n4689) );
  NBUFFX2 U3952 ( .IN(n4706), .Q(n4669) );
  NBUFFX2 U3953 ( .IN(n4705), .Q(n4670) );
  NBUFFX2 U3954 ( .IN(n4705), .Q(n4671) );
  NBUFFX2 U3955 ( .IN(n4700), .Q(n4680) );
  NBUFFX2 U3956 ( .IN(n4702), .Q(n4676) );
  NBUFFX2 U3957 ( .IN(n4702), .Q(n4677) );
  NBUFFX2 U3958 ( .IN(n4698), .Q(n4685) );
  NBUFFX2 U3959 ( .IN(n4708), .Q(n4664) );
  NBUFFX2 U3960 ( .IN(n4697), .Q(n4686) );
  NBUFFX2 U3961 ( .IN(n4701), .Q(n4678) );
  NBUFFX2 U3962 ( .IN(n4697), .Q(n4687) );
  NBUFFX2 U3963 ( .IN(n4709), .Q(n4663) );
  NBUFFX2 U3964 ( .IN(n4709), .Q(n4662) );
  NBUFFX2 U3965 ( .IN(n4710), .Q(n4661) );
  NBUFFX2 U3966 ( .IN(n4704), .Q(n4672) );
  NBUFFX2 U3967 ( .IN(n4704), .Q(n4673) );
  NBUFFX2 U3968 ( .IN(n4696), .Q(n4688) );
  NBUFFX2 U3969 ( .IN(n4707), .Q(n4666) );
  NBUFFX2 U3970 ( .IN(n4706), .Q(n4668) );
  NBUFFX2 U3971 ( .IN(n4703), .Q(n4675) );
  NBUFFX2 U3972 ( .IN(n4703), .Q(n4674) );
  NBUFFX2 U3973 ( .IN(n4695), .Q(n4691) );
  NBUFFX2 U3974 ( .IN(n4715), .Q(n4651) );
  NBUFFX2 U3975 ( .IN(n4715), .Q(n4650) );
  NBUFFX2 U3976 ( .IN(n4710), .Q(n4660) );
  NBUFFX2 U3977 ( .IN(n4711), .Q(n4659) );
  NBUFFX2 U3978 ( .IN(n4711), .Q(n4658) );
  NBUFFX2 U3979 ( .IN(n4712), .Q(n4657) );
  NBUFFX2 U3980 ( .IN(n4712), .Q(n4656) );
  NBUFFX2 U3981 ( .IN(n4713), .Q(n4655) );
  NBUFFX2 U3982 ( .IN(n4718), .Q(n4644) );
  NBUFFX2 U3983 ( .IN(n4719), .Q(n4643) );
  NBUFFX2 U3984 ( .IN(n4719), .Q(n4642) );
  NBUFFX2 U3985 ( .IN(n4720), .Q(n4641) );
  NBUFFX2 U3986 ( .IN(n4695), .Q(n4690) );
  NBUFFX2 U3987 ( .IN(n4717), .Q(n4647) );
  NBUFFX2 U3988 ( .IN(n4717), .Q(n4646) );
  INVX0 U3989 ( .IN(n4753), .QN(n4743) );
  INVX0 U3990 ( .IN(n4771), .QN(n4766) );
  ISOLANDX1 U3991 ( .D(n3278), .ISO(n4774), .Q(n2152) );
  NBUFFX2 U3992 ( .IN(n2148), .Q(n4522) );
  NBUFFX2 U3993 ( .IN(n2148), .Q(n4528) );
  NBUFFX2 U3994 ( .IN(n2148), .Q(n4527) );
  NBUFFX2 U3995 ( .IN(n2148), .Q(n4524) );
  NBUFFX2 U3996 ( .IN(n2148), .Q(n4523) );
  NBUFFX2 U3997 ( .IN(n2148), .Q(n4526) );
  NBUFFX2 U3998 ( .IN(n2148), .Q(n4525) );
  NBUFFX2 U3999 ( .IN(n4415), .Q(n4399) );
  NBUFFX2 U4000 ( .IN(n4414), .Q(n4401) );
  NBUFFX2 U4001 ( .IN(n4413), .Q(n4402) );
  NBUFFX2 U4002 ( .IN(n4413), .Q(n4403) );
  NBUFFX2 U4003 ( .IN(n4409), .Q(n4357) );
  NBUFFX2 U4004 ( .IN(n4412), .Q(n4404) );
  NBUFFX2 U4005 ( .IN(n4412), .Q(n4405) );
  NBUFFX2 U4006 ( .IN(n4418), .Q(n4392) );
  NBUFFX2 U4007 ( .IN(n4418), .Q(n4393) );
  NBUFFX2 U4008 ( .IN(n4417), .Q(n4394) );
  NBUFFX2 U4009 ( .IN(n4417), .Q(n4395) );
  NBUFFX2 U4010 ( .IN(n4414), .Q(n4400) );
  NBUFFX2 U4011 ( .IN(n4732), .Q(n4701) );
  NBUFFX2 U4012 ( .IN(n4416), .Q(n4396) );
  NBUFFX2 U4013 ( .IN(n4416), .Q(n4397) );
  NBUFFX2 U4014 ( .IN(n4415), .Q(n4398) );
  NBUFFX2 U4015 ( .IN(n4411), .Q(n4406) );
  NBUFFX2 U4016 ( .IN(n4411), .Q(n4407) );
  NBUFFX2 U4017 ( .IN(n4409), .Q(n4356) );
  NBUFFX2 U4018 ( .IN(n4408), .Q(n4359) );
  NBUFFX2 U4019 ( .IN(n4408), .Q(n4358) );
  INVX0 U4020 ( .IN(n4754), .QN(n4744) );
  INVX0 U4021 ( .IN(n4755), .QN(n4745) );
  INVX0 U4022 ( .IN(n4756), .QN(n4746) );
  INVX0 U4023 ( .IN(n4757), .QN(n4747) );
  INVX0 U4024 ( .IN(n4758), .QN(n4748) );
  INVX0 U4025 ( .IN(n4759), .QN(n4749) );
  INVX0 U4026 ( .IN(n4772), .QN(n4768) );
  INVX0 U4027 ( .IN(n4770), .QN(n4767) );
  NBUFFX2 U4028 ( .IN(n4725), .Q(n4714) );
  NBUFFX2 U4029 ( .IN(n4724), .Q(n4716) );
  NBUFFX2 U4030 ( .IN(n4733), .Q(n4699) );
  NBUFFX2 U4031 ( .IN(n4735), .Q(n4694) );
  NBUFFX2 U4032 ( .IN(n4730), .Q(n4705) );
  NBUFFX2 U4033 ( .IN(n4732), .Q(n4700) );
  NBUFFX2 U4034 ( .IN(n4731), .Q(n4702) );
  NBUFFX2 U4035 ( .IN(n4733), .Q(n4698) );
  NBUFFX2 U4036 ( .IN(n4728), .Q(n4708) );
  NBUFFX2 U4037 ( .IN(n4734), .Q(n4697) );
  NBUFFX2 U4038 ( .IN(n4728), .Q(n4709) );
  NBUFFX2 U4039 ( .IN(n4730), .Q(n4704) );
  NBUFFX2 U4040 ( .IN(n4734), .Q(n4696) );
  NBUFFX2 U4041 ( .IN(n4729), .Q(n4707) );
  NBUFFX2 U4042 ( .IN(n4729), .Q(n4706) );
  NBUFFX2 U4043 ( .IN(n4731), .Q(n4703) );
  NBUFFX2 U4044 ( .IN(n4725), .Q(n4715) );
  NBUFFX2 U4045 ( .IN(n4727), .Q(n4710) );
  NBUFFX2 U4046 ( .IN(n4727), .Q(n4711) );
  NBUFFX2 U4047 ( .IN(n4726), .Q(n4712) );
  NBUFFX2 U4048 ( .IN(n4726), .Q(n4713) );
  NBUFFX2 U4049 ( .IN(n4723), .Q(n4718) );
  NBUFFX2 U4050 ( .IN(n4723), .Q(n4719) );
  NBUFFX2 U4051 ( .IN(n4722), .Q(n4720) );
  NBUFFX2 U4052 ( .IN(n4735), .Q(n4695) );
  NBUFFX2 U4053 ( .IN(n4724), .Q(n4717) );
  NBUFFX2 U4054 ( .IN(n4721), .Q(n4639) );
  NBUFFX2 U4055 ( .IN(n4722), .Q(n4721) );
  NOR2X0 U4056 ( .IN1(n4752), .IN2(n4775), .QN(n2148) );
  INVX0 U4057 ( .IN(n4779), .QN(n4771) );
  INVX0 U4058 ( .IN(TM0), .QN(n4772) );
  INVX0 U4059 ( .IN(n4779), .QN(n4770) );
  INVX0 U4060 ( .IN(TM1), .QN(n4753) );
  INVX0 U4061 ( .IN(n4763), .QN(n4754) );
  INVX0 U4062 ( .IN(n4763), .QN(n4755) );
  INVX0 U4063 ( .IN(n4764), .QN(n4756) );
  INVX0 U4064 ( .IN(n4764), .QN(n4757) );
  INVX0 U4065 ( .IN(n4763), .QN(n4758) );
  INVX0 U4066 ( .IN(n4763), .QN(n4759) );
  INVX0 U4067 ( .IN(n4778), .QN(n4773) );
  INVX0 U4068 ( .IN(n4778), .QN(n4774) );
  INVX0 U4069 ( .IN(TM1), .QN(n4752) );
  INVX0 U4070 ( .IN(n4778), .QN(n4775) );
  NBUFFX2 U4071 ( .IN(n4421), .Q(n4413) );
  NBUFFX2 U4072 ( .IN(n4422), .Q(n4412) );
  NBUFFX2 U4073 ( .IN(n4419), .Q(n4418) );
  NBUFFX2 U4074 ( .IN(n4419), .Q(n4417) );
  NBUFFX2 U4075 ( .IN(n4421), .Q(n4414) );
  NBUFFX2 U4076 ( .IN(n4737), .Q(n4732) );
  NBUFFX2 U4077 ( .IN(n4420), .Q(n4416) );
  NBUFFX2 U4078 ( .IN(n4420), .Q(n4415) );
  NBUFFX2 U4079 ( .IN(n4422), .Q(n4411) );
  NBUFFX2 U4080 ( .IN(n4410), .Q(n4409) );
  NBUFFX2 U4081 ( .IN(n4410), .Q(n4408) );
  INVX0 U4082 ( .IN(n4760), .QN(n4750) );
  INVX0 U4083 ( .IN(n4776), .QN(n4769) );
  NBUFFX2 U4084 ( .IN(n4737), .Q(n4733) );
  NBUFFX2 U4085 ( .IN(n4739), .Q(n4728) );
  NBUFFX2 U4086 ( .IN(n4738), .Q(n4730) );
  NBUFFX2 U4087 ( .IN(n4736), .Q(n4734) );
  NBUFFX2 U4088 ( .IN(n4739), .Q(n4729) );
  NBUFFX2 U4089 ( .IN(n4738), .Q(n4731) );
  NBUFFX2 U4090 ( .IN(n4741), .Q(n4725) );
  NBUFFX2 U4091 ( .IN(n4740), .Q(n4727) );
  NBUFFX2 U4092 ( .IN(n4740), .Q(n4726) );
  NBUFFX2 U4093 ( .IN(n4742), .Q(n4723) );
  NBUFFX2 U4094 ( .IN(n4742), .Q(n4722) );
  NBUFFX2 U4095 ( .IN(n4736), .Q(n4735) );
  NBUFFX2 U4096 ( .IN(n4741), .Q(n4724) );
  INVX0 U4097 ( .IN(n4762), .QN(n4760) );
  INVX0 U4098 ( .IN(n4778), .QN(n4776) );
  INVX0 U4099 ( .IN(n4778), .QN(n4777) );
  INVX0 U4100 ( .IN(n4780), .QN(n4779) );
  INVX0 U4101 ( .IN(n4780), .QN(n4778) );
  INVX0 U4102 ( .IN(n4760), .QN(n4764) );
  INVX0 U4103 ( .IN(n4752), .QN(n4763) );
  INVX0 U4104 ( .IN(n4761), .QN(n4751) );
  INVX0 U4105 ( .IN(n4762), .QN(n4761) );
  NBUFFX2 U4106 ( .IN(n2149), .Q(n4419) );
  NBUFFX2 U4107 ( .IN(n2149), .Q(n4421) );
  NBUFFX2 U4108 ( .IN(n2149), .Q(n4420) );
  NBUFFX2 U4109 ( .IN(n2149), .Q(n4422) );
  NBUFFX2 U4110 ( .IN(n1729), .Q(n4737) );
  NBUFFX2 U4111 ( .IN(n4423), .Q(n4410) );
  NBUFFX2 U4112 ( .IN(n2149), .Q(n4423) );
  NOR2X0 U4113 ( .IN1(n4568), .IN2(n3346), .QN(WX11082) );
  NOR2X0 U4114 ( .IN1(n4568), .IN2(n3347), .QN(WX11080) );
  NOR2X0 U4115 ( .IN1(n4568), .IN2(n3348), .QN(WX11078) );
  NOR2X0 U4116 ( .IN1(n4557), .IN2(n3349), .QN(WX11076) );
  NOR2X0 U4117 ( .IN1(n4556), .IN2(n3350), .QN(WX11074) );
  NOR2X0 U4118 ( .IN1(n4557), .IN2(n3351), .QN(WX11072) );
  NOR2X0 U4119 ( .IN1(n4558), .IN2(n3352), .QN(WX11070) );
  NOR2X0 U4120 ( .IN1(n4556), .IN2(n3353), .QN(WX11068) );
  NOR2X0 U4121 ( .IN1(n4556), .IN2(n3354), .QN(WX11066) );
  NOR2X0 U4122 ( .IN1(n4556), .IN2(n3355), .QN(WX11064) );
  NOR2X0 U4123 ( .IN1(n4557), .IN2(n3356), .QN(WX11062) );
  NOR2X0 U4124 ( .IN1(n4557), .IN2(n3357), .QN(WX11060) );
  NOR2X0 U4125 ( .IN1(n4557), .IN2(n3358), .QN(WX11058) );
  NOR2X0 U4126 ( .IN1(n4558), .IN2(n3359), .QN(WX11056) );
  NOR2X0 U4127 ( .IN1(n4557), .IN2(n3360), .QN(WX11054) );
  NOR2X0 U4128 ( .IN1(n4557), .IN2(n3338), .QN(WX11052) );
  NOR2X0 U4129 ( .IN1(n4557), .IN2(n3361), .QN(WX9789) );
  NOR2X0 U4130 ( .IN1(n4556), .IN2(n3362), .QN(WX9787) );
  NOR2X0 U4131 ( .IN1(n4556), .IN2(n3363), .QN(WX9785) );
  NOR2X0 U4132 ( .IN1(n4556), .IN2(n3364), .QN(WX9783) );
  NOR2X0 U4133 ( .IN1(n4556), .IN2(n3365), .QN(WX9781) );
  NOR2X0 U4134 ( .IN1(n4563), .IN2(n3366), .QN(WX9779) );
  NOR2X0 U4135 ( .IN1(n4570), .IN2(n3367), .QN(WX9777) );
  NOR2X0 U4136 ( .IN1(n4570), .IN2(n3368), .QN(WX9775) );
  NOR2X0 U4137 ( .IN1(n4570), .IN2(n3370), .QN(WX9771) );
  NOR2X0 U4138 ( .IN1(n4569), .IN2(n3372), .QN(WX9767) );
  NOR2X0 U4139 ( .IN1(n4568), .IN2(n3373), .QN(WX9765) );
  NOR2X0 U4140 ( .IN1(n4569), .IN2(n3374), .QN(WX9763) );
  NOR2X0 U4141 ( .IN1(n4569), .IN2(n3375), .QN(WX9761) );
  NOR2X0 U4142 ( .IN1(n4569), .IN2(n3339), .QN(WX9759) );
  NOR2X0 U4143 ( .IN1(n4566), .IN2(n3376), .QN(WX8496) );
  NOR2X0 U4144 ( .IN1(n4566), .IN2(n3377), .QN(WX8494) );
  NOR2X0 U4145 ( .IN1(n4566), .IN2(n3378), .QN(WX8492) );
  NOR2X0 U4146 ( .IN1(n4566), .IN2(n3379), .QN(WX8490) );
  NOR2X0 U4147 ( .IN1(n4566), .IN2(n3380), .QN(WX8488) );
  NOR2X0 U4148 ( .IN1(n4566), .IN2(n3381), .QN(WX8486) );
  NOR2X0 U4149 ( .IN1(n4566), .IN2(n3382), .QN(WX8484) );
  NOR2X0 U4150 ( .IN1(n4566), .IN2(n3383), .QN(WX8482) );
  NOR2X0 U4151 ( .IN1(n4566), .IN2(n3384), .QN(WX8480) );
  NOR2X0 U4152 ( .IN1(n4565), .IN2(n3385), .QN(WX8478) );
  NOR2X0 U4153 ( .IN1(n4565), .IN2(n3386), .QN(WX8476) );
  NOR2X0 U4154 ( .IN1(n4565), .IN2(n3387), .QN(WX8474) );
  NOR2X0 U4155 ( .IN1(n4565), .IN2(n3388), .QN(WX8472) );
  NOR2X0 U4156 ( .IN1(n4565), .IN2(n3389), .QN(WX8470) );
  NOR2X0 U4157 ( .IN1(n4565), .IN2(n3390), .QN(WX8468) );
  NOR2X0 U4158 ( .IN1(n4565), .IN2(n3340), .QN(WX8466) );
  NOR2X0 U4159 ( .IN1(n4560), .IN2(n3391), .QN(WX7203) );
  NOR2X0 U4160 ( .IN1(n4560), .IN2(n3392), .QN(WX7201) );
  NOR2X0 U4161 ( .IN1(n4560), .IN2(n3393), .QN(WX7199) );
  NOR2X0 U4162 ( .IN1(n4560), .IN2(n3394), .QN(WX7197) );
  NOR2X0 U4163 ( .IN1(n4560), .IN2(n3395), .QN(WX7195) );
  NOR2X0 U4164 ( .IN1(n4560), .IN2(n3396), .QN(WX7193) );
  NOR2X0 U4165 ( .IN1(n4561), .IN2(n3397), .QN(WX7191) );
  NOR2X0 U4166 ( .IN1(n4561), .IN2(n3398), .QN(WX7189) );
  NOR2X0 U4167 ( .IN1(n4561), .IN2(n3399), .QN(WX7187) );
  NOR2X0 U4168 ( .IN1(n4561), .IN2(n3400), .QN(WX7185) );
  NOR2X0 U4169 ( .IN1(n4561), .IN2(n3401), .QN(WX7183) );
  NOR2X0 U4170 ( .IN1(n4561), .IN2(n3402), .QN(WX7181) );
  NOR2X0 U4171 ( .IN1(n4561), .IN2(n3403), .QN(WX7179) );
  NOR2X0 U4172 ( .IN1(n4561), .IN2(n3404), .QN(WX7177) );
  NOR2X0 U4173 ( .IN1(n4561), .IN2(n3405), .QN(WX7175) );
  NOR2X0 U4174 ( .IN1(n4561), .IN2(n3341), .QN(WX7173) );
  NOR2X0 U4175 ( .IN1(n4559), .IN2(n3406), .QN(WX5910) );
  NOR2X0 U4176 ( .IN1(n4559), .IN2(n3407), .QN(WX5908) );
  NOR2X0 U4177 ( .IN1(n4559), .IN2(n3408), .QN(WX5906) );
  NOR2X0 U4178 ( .IN1(n4559), .IN2(n3409), .QN(WX5904) );
  NOR2X0 U4179 ( .IN1(n4559), .IN2(n3410), .QN(WX5902) );
  NOR2X0 U4180 ( .IN1(n4559), .IN2(n3411), .QN(WX5900) );
  NOR2X0 U4181 ( .IN1(n4559), .IN2(n3412), .QN(WX5898) );
  NOR2X0 U4182 ( .IN1(n4559), .IN2(n3413), .QN(WX5896) );
  NOR2X0 U4183 ( .IN1(n4558), .IN2(n3414), .QN(WX5894) );
  NOR2X0 U4184 ( .IN1(n4559), .IN2(n3415), .QN(WX5892) );
  NOR2X0 U4185 ( .IN1(n4558), .IN2(n3416), .QN(WX5890) );
  NOR2X0 U4186 ( .IN1(n4557), .IN2(n3417), .QN(WX5888) );
  NOR2X0 U4187 ( .IN1(n4556), .IN2(n3418), .QN(WX5886) );
  NOR2X0 U4188 ( .IN1(n4568), .IN2(n3420), .QN(WX5882) );
  NOR2X0 U4189 ( .IN1(n4560), .IN2(n3421), .QN(WX4617) );
  NOR2X0 U4190 ( .IN1(n4558), .IN2(n3422), .QN(WX4615) );
  NOR2X0 U4191 ( .IN1(n4558), .IN2(n3423), .QN(WX4613) );
  NOR2X0 U4192 ( .IN1(n4559), .IN2(n3424), .QN(WX4611) );
  NOR2X0 U4193 ( .IN1(n4558), .IN2(n3425), .QN(WX4609) );
  NOR2X0 U4194 ( .IN1(n4568), .IN2(n3426), .QN(WX4607) );
  NOR2X0 U4195 ( .IN1(n4568), .IN2(n3427), .QN(WX4605) );
  NOR2X0 U4196 ( .IN1(n4565), .IN2(n3428), .QN(WX4603) );
  NOR2X0 U4197 ( .IN1(n4564), .IN2(n3429), .QN(WX4601) );
  NOR2X0 U4198 ( .IN1(n4564), .IN2(n3430), .QN(WX4599) );
  NOR2X0 U4199 ( .IN1(n4564), .IN2(n3431), .QN(WX4597) );
  NOR2X0 U4200 ( .IN1(n4564), .IN2(n3432), .QN(WX4595) );
  NOR2X0 U4201 ( .IN1(n4564), .IN2(n3433), .QN(WX4593) );
  NOR2X0 U4202 ( .IN1(n4564), .IN2(n3434), .QN(WX4591) );
  NOR2X0 U4203 ( .IN1(n4564), .IN2(n3435), .QN(WX4589) );
  NOR2X0 U4204 ( .IN1(n4565), .IN2(n3343), .QN(WX4587) );
  NOR2X0 U4205 ( .IN1(n4562), .IN2(n3436), .QN(WX3324) );
  NOR2X0 U4206 ( .IN1(n4562), .IN2(n3437), .QN(WX3322) );
  NOR2X0 U4207 ( .IN1(n4564), .IN2(n3438), .QN(WX3320) );
  NOR2X0 U4208 ( .IN1(n4562), .IN2(n3439), .QN(WX3318) );
  NOR2X0 U4209 ( .IN1(n4562), .IN2(n3440), .QN(WX3316) );
  NOR2X0 U4210 ( .IN1(n4562), .IN2(n3441), .QN(WX3314) );
  NOR2X0 U4211 ( .IN1(n4563), .IN2(n3442), .QN(WX3312) );
  NOR2X0 U4212 ( .IN1(n4564), .IN2(n3443), .QN(WX3310) );
  NOR2X0 U4213 ( .IN1(n4556), .IN2(n3444), .QN(WX3308) );
  NOR2X0 U4214 ( .IN1(n4563), .IN2(n3445), .QN(WX3306) );
  NOR2X0 U4215 ( .IN1(n4563), .IN2(n3446), .QN(WX3304) );
  NOR2X0 U4216 ( .IN1(n4563), .IN2(n3447), .QN(WX3302) );
  NOR2X0 U4217 ( .IN1(n4563), .IN2(n3448), .QN(WX3300) );
  NOR2X0 U4218 ( .IN1(n4563), .IN2(n3449), .QN(WX3298) );
  NOR2X0 U4219 ( .IN1(n4563), .IN2(n3450), .QN(WX3296) );
  NOR2X0 U4220 ( .IN1(n4562), .IN2(n3344), .QN(WX3294) );
  NOR2X0 U4221 ( .IN1(n4570), .IN2(n3451), .QN(WX2031) );
  NOR2X0 U4222 ( .IN1(n4569), .IN2(n3453), .QN(WX2027) );
  NOR2X0 U4223 ( .IN1(n4568), .IN2(n3454), .QN(WX2025) );
  NOR2X0 U4224 ( .IN1(n4570), .IN2(n3455), .QN(WX2023) );
  NOR2X0 U4225 ( .IN1(n4569), .IN2(n3456), .QN(WX2021) );
  NOR2X0 U4226 ( .IN1(n4570), .IN2(n3457), .QN(WX2019) );
  NOR2X0 U4227 ( .IN1(n4570), .IN2(n3458), .QN(WX2017) );
  NOR2X0 U4228 ( .IN1(n4569), .IN2(n3459), .QN(WX2015) );
  NOR2X0 U4229 ( .IN1(n4570), .IN2(n3460), .QN(WX2013) );
  NOR2X0 U4230 ( .IN1(n4568), .IN2(n3461), .QN(WX2011) );
  NOR2X0 U4231 ( .IN1(n4569), .IN2(n3462), .QN(WX2009) );
  NOR2X0 U4232 ( .IN1(n4570), .IN2(n3463), .QN(WX2007) );
  NOR2X0 U4233 ( .IN1(n4570), .IN2(n3464), .QN(WX2005) );
  NOR2X0 U4234 ( .IN1(n4569), .IN2(n3465), .QN(WX2003) );
  NOR2X0 U4235 ( .IN1(n4569), .IN2(n3345), .QN(WX2001) );
  NOR2X0 U4236 ( .IN1(n4571), .IN2(n3369), .QN(WX9773) );
  NOR2X0 U4237 ( .IN1(n4571), .IN2(n3371), .QN(WX9769) );
  NOR2X0 U4238 ( .IN1(n4571), .IN2(n3419), .QN(WX5884) );
  NOR2X0 U4239 ( .IN1(n4571), .IN2(n3342), .QN(WX5880) );
  NOR2X0 U4240 ( .IN1(n4571), .IN2(n3452), .QN(WX2029) );
  NBUFFX2 U4241 ( .IN(n1729), .Q(n4739) );
  NBUFFX2 U4242 ( .IN(n1729), .Q(n4738) );
  NBUFFX2 U4243 ( .IN(n1729), .Q(n4740) );
  NBUFFX2 U4244 ( .IN(n1729), .Q(n4742) );
  NBUFFX2 U4245 ( .IN(n1729), .Q(n4736) );
  NBUFFX2 U4246 ( .IN(n1729), .Q(n4741) );
  XNOR2X1 U4247 ( .IN1(n3179), .IN2(n2532), .Q(DATA_9_9) );
  NAND2X0 U4248 ( .IN1(WX529), .IN2(n4767), .QN(n3179) );
  XNOR2X1 U4249 ( .IN1(n3161), .IN2(n2529), .Q(DATA_9_8) );
  NAND2X0 U4250 ( .IN1(WX531), .IN2(n4766), .QN(n3161) );
  XNOR2X1 U4251 ( .IN1(n3159), .IN2(n2526), .Q(DATA_9_7) );
  NAND2X0 U4252 ( .IN1(WX533), .IN2(n4766), .QN(n3159) );
  XNOR2X1 U4253 ( .IN1(n3157), .IN2(n2523), .Q(DATA_9_6) );
  NAND2X0 U4254 ( .IN1(WX535), .IN2(n4766), .QN(n3157) );
  XNOR2X1 U4255 ( .IN1(n3155), .IN2(n2520), .Q(DATA_9_5) );
  NAND2X0 U4256 ( .IN1(WX537), .IN2(n4766), .QN(n3155) );
  XNOR2X1 U4257 ( .IN1(n3153), .IN2(n2517), .Q(DATA_9_4) );
  NAND2X0 U4258 ( .IN1(WX539), .IN2(n4766), .QN(n3153) );
  XNOR2X1 U4259 ( .IN1(n3336), .IN2(n2630), .Q(DATA_9_31) );
  NAND2X0 U4260 ( .IN1(WX485), .IN2(n4766), .QN(n3336) );
  XNOR2X1 U4261 ( .IN1(n3334), .IN2(n2615), .Q(DATA_9_30) );
  NAND2X0 U4262 ( .IN1(WX487), .IN2(n4769), .QN(n3334) );
  XNOR2X1 U4263 ( .IN1(n3151), .IN2(n2514), .Q(DATA_9_3) );
  NAND2X0 U4264 ( .IN1(WX541), .IN2(n4766), .QN(n3151) );
  XNOR2X1 U4265 ( .IN1(n3332), .IN2(n2602), .Q(DATA_9_29) );
  NAND2X0 U4266 ( .IN1(WX489), .IN2(n4769), .QN(n3332) );
  XNOR2X1 U4267 ( .IN1(n3330), .IN2(n2589), .Q(DATA_9_28) );
  NAND2X0 U4268 ( .IN1(WX491), .IN2(n4769), .QN(n3330) );
  XNOR2X1 U4269 ( .IN1(n3296), .IN2(n2586), .Q(DATA_9_27) );
  NAND2X0 U4270 ( .IN1(WX493), .IN2(n4768), .QN(n3296) );
  XNOR2X1 U4271 ( .IN1(n3294), .IN2(n2583), .Q(DATA_9_26) );
  NAND2X0 U4272 ( .IN1(WX495), .IN2(n4769), .QN(n3294) );
  XNOR2X1 U4273 ( .IN1(n3292), .IN2(n2580), .Q(DATA_9_25) );
  NAND2X0 U4274 ( .IN1(WX497), .IN2(n4769), .QN(n3292) );
  XNOR2X1 U4275 ( .IN1(n3290), .IN2(n2577), .Q(DATA_9_24) );
  NAND2X0 U4276 ( .IN1(WX499), .IN2(n4768), .QN(n3290) );
  XNOR2X1 U4277 ( .IN1(n3288), .IN2(n2574), .Q(DATA_9_23) );
  NAND2X0 U4278 ( .IN1(WX501), .IN2(n4768), .QN(n3288) );
  XNOR2X1 U4279 ( .IN1(n3286), .IN2(n2571), .Q(DATA_9_22) );
  NAND2X0 U4280 ( .IN1(WX503), .IN2(n4768), .QN(n3286) );
  XNOR2X1 U4281 ( .IN1(n3284), .IN2(n2568), .Q(DATA_9_21) );
  NAND2X0 U4282 ( .IN1(WX505), .IN2(n4768), .QN(n3284) );
  XNOR2X1 U4283 ( .IN1(n3282), .IN2(n2565), .Q(DATA_9_20) );
  NAND2X0 U4284 ( .IN1(WX507), .IN2(n4768), .QN(n3282) );
  XNOR2X1 U4285 ( .IN1(n3149), .IN2(n2511), .Q(DATA_9_2) );
  NAND2X0 U4286 ( .IN1(WX543), .IN2(n4766), .QN(n3149) );
  XNOR2X1 U4287 ( .IN1(n3280), .IN2(n2562), .Q(DATA_9_19) );
  NAND2X0 U4288 ( .IN1(WX509), .IN2(n4768), .QN(n3280) );
  XNOR2X1 U4289 ( .IN1(n3255), .IN2(n2559), .Q(DATA_9_18) );
  NAND2X0 U4290 ( .IN1(WX511), .IN2(n4768), .QN(n3255) );
  XNOR2X1 U4291 ( .IN1(n3211), .IN2(n2556), .Q(DATA_9_17) );
  NAND2X0 U4292 ( .IN1(WX513), .IN2(n4768), .QN(n3211) );
  XNOR2X1 U4293 ( .IN1(n3209), .IN2(n2553), .Q(DATA_9_16) );
  NAND2X0 U4294 ( .IN1(WX515), .IN2(n4767), .QN(n3209) );
  XNOR2X1 U4295 ( .IN1(n3207), .IN2(n2550), .Q(DATA_9_15) );
  NAND2X0 U4296 ( .IN1(WX517), .IN2(n4767), .QN(n3207) );
  XNOR2X1 U4297 ( .IN1(n3205), .IN2(n2547), .Q(DATA_9_14) );
  NAND2X0 U4298 ( .IN1(test_so1), .IN2(n4767), .QN(n3205) );
  XNOR2X1 U4299 ( .IN1(n3203), .IN2(n2544), .Q(DATA_9_13) );
  NAND2X0 U4300 ( .IN1(WX521), .IN2(n4767), .QN(n3203) );
  XNOR2X1 U4301 ( .IN1(n3201), .IN2(n2541), .Q(DATA_9_12) );
  NAND2X0 U4302 ( .IN1(WX523), .IN2(n4767), .QN(n3201) );
  XNOR2X1 U4303 ( .IN1(n3199), .IN2(n2538), .Q(DATA_9_11) );
  NAND2X0 U4304 ( .IN1(WX525), .IN2(n4767), .QN(n3199) );
  XNOR2X1 U4305 ( .IN1(n3197), .IN2(n2535), .Q(DATA_9_10) );
  NAND2X0 U4306 ( .IN1(WX527), .IN2(n4767), .QN(n3197) );
  XNOR2X1 U4307 ( .IN1(n3147), .IN2(n2508), .Q(DATA_9_1) );
  NAND2X0 U4308 ( .IN1(WX545), .IN2(n4766), .QN(n3147) );
  XNOR2X1 U4309 ( .IN1(n3145), .IN2(n2505), .Q(DATA_9_0) );
  NAND2X0 U4310 ( .IN1(WX547), .IN2(n4767), .QN(n3145) );
  AND3X1 U4311 ( .IN1(RESET), .IN2(n4773), .IN3(n4751), .Q(n2149) );
  INVX0 U4312 ( .IN(n4765), .QN(n4762) );
  INVX0 U4313 ( .IN(TM1), .QN(n4765) );
  INVX0 U4314 ( .IN(TM0), .QN(n4780) );
  XNOR3X1 U4315 ( .IN1(n3466), .IN2(n4775), .IN3(n3467), .Q(n2505) );
  XNOR3X1 U4316 ( .IN1(WX899), .IN2(WX835), .IN3(WX771), .Q(n3466) );
  XNOR3X1 U4317 ( .IN1(n3468), .IN2(n4770), .IN3(n3469), .Q(n2508) );
  XNOR3X1 U4318 ( .IN1(WX897), .IN2(WX833), .IN3(WX769), .Q(n3468) );
  XNOR3X1 U4319 ( .IN1(n3470), .IN2(n4770), .IN3(n3471), .Q(n2511) );
  XNOR3X1 U4320 ( .IN1(WX895), .IN2(test_so7), .IN3(WX767), .Q(n3470) );
  XNOR3X1 U4321 ( .IN1(n3472), .IN2(n4771), .IN3(n3473), .Q(n2514) );
  XNOR3X1 U4322 ( .IN1(WX893), .IN2(WX829), .IN3(WX765), .Q(n3472) );
  XNOR3X1 U4323 ( .IN1(n3474), .IN2(n4771), .IN3(n3475), .Q(n2517) );
  XNOR3X1 U4324 ( .IN1(WX891), .IN2(WX827), .IN3(WX763), .Q(n3474) );
  XNOR3X1 U4325 ( .IN1(n3476), .IN2(n4772), .IN3(n3477), .Q(n2520) );
  XNOR3X1 U4326 ( .IN1(WX889), .IN2(WX825), .IN3(WX761), .Q(n3476) );
  XNOR3X1 U4327 ( .IN1(n3478), .IN2(n4772), .IN3(n3479), .Q(n2523) );
  XNOR3X1 U4328 ( .IN1(WX887), .IN2(WX823), .IN3(test_so5), .Q(n3478) );
  XNOR3X1 U4329 ( .IN1(n3480), .IN2(n4773), .IN3(n3481), .Q(n2526) );
  XNOR3X1 U4330 ( .IN1(WX885), .IN2(WX821), .IN3(WX757), .Q(n3480) );
  XNOR3X1 U4331 ( .IN1(n3482), .IN2(n4773), .IN3(n3483), .Q(n2529) );
  XNOR3X1 U4332 ( .IN1(WX883), .IN2(WX819), .IN3(WX755), .Q(n3482) );
  XNOR3X1 U4333 ( .IN1(n3484), .IN2(n4774), .IN3(n3485), .Q(n2532) );
  XNOR3X1 U4334 ( .IN1(WX881), .IN2(WX817), .IN3(WX753), .Q(n3484) );
  XNOR3X1 U4335 ( .IN1(n3486), .IN2(n4774), .IN3(n3487), .Q(n2535) );
  XNOR3X1 U4336 ( .IN1(WX879), .IN2(WX815), .IN3(WX751), .Q(n3486) );
  XNOR3X1 U4337 ( .IN1(n3488), .IN2(n4775), .IN3(n3489), .Q(n2538) );
  XNOR3X1 U4338 ( .IN1(WX877), .IN2(WX813), .IN3(WX749), .Q(n3488) );
  XNOR3X1 U4339 ( .IN1(n3490), .IN2(n4776), .IN3(n3491), .Q(n2541) );
  XNOR3X1 U4340 ( .IN1(WX875), .IN2(WX811), .IN3(WX747), .Q(n3490) );
  XNOR3X1 U4341 ( .IN1(n3492), .IN2(n4776), .IN3(n3493), .Q(n2544) );
  XNOR3X1 U4342 ( .IN1(WX873), .IN2(WX809), .IN3(WX745), .Q(n3492) );
  XNOR3X1 U4343 ( .IN1(n3494), .IN2(n4777), .IN3(n3495), .Q(n2547) );
  XNOR3X1 U4344 ( .IN1(WX871), .IN2(WX807), .IN3(WX743), .Q(n3494) );
  XNOR3X1 U4345 ( .IN1(n3496), .IN2(n4777), .IN3(n3497), .Q(n2550) );
  XNOR3X1 U4346 ( .IN1(WX869), .IN2(WX805), .IN3(WX741), .Q(n3496) );
  XNOR3X1 U4347 ( .IN1(n3498), .IN2(n4758), .IN3(n3499), .Q(n2553) );
  XNOR3X1 U4348 ( .IN1(test_so8), .IN2(WX803), .IN3(WX739), .Q(n3498) );
  XNOR3X1 U4349 ( .IN1(n3500), .IN2(n4753), .IN3(n3501), .Q(n2556) );
  XNOR3X1 U4350 ( .IN1(WX865), .IN2(WX801), .IN3(WX737), .Q(n3500) );
  XNOR3X1 U4351 ( .IN1(n3502), .IN2(n4752), .IN3(n3503), .Q(n2559) );
  XNOR3X1 U4352 ( .IN1(WX863), .IN2(WX799), .IN3(WX735), .Q(n3502) );
  XNOR3X1 U4353 ( .IN1(n3504), .IN2(n4753), .IN3(n3505), .Q(n2562) );
  XNOR3X1 U4354 ( .IN1(WX861), .IN2(WX797), .IN3(WX733), .Q(n3504) );
  XNOR3X1 U4355 ( .IN1(n3506), .IN2(n4754), .IN3(n3507), .Q(n2565) );
  XNOR3X1 U4356 ( .IN1(WX859), .IN2(test_so6), .IN3(WX731), .Q(n3506) );
  XNOR3X1 U4357 ( .IN1(n3508), .IN2(n4754), .IN3(n3509), .Q(n2568) );
  XNOR3X1 U4358 ( .IN1(WX857), .IN2(WX793), .IN3(WX729), .Q(n3508) );
  XNOR3X1 U4359 ( .IN1(n3510), .IN2(n4755), .IN3(n3511), .Q(n2571) );
  XNOR3X1 U4360 ( .IN1(WX855), .IN2(WX791), .IN3(WX727), .Q(n3510) );
  XNOR3X1 U4361 ( .IN1(n3512), .IN2(n4755), .IN3(n3513), .Q(n2574) );
  XNOR3X1 U4362 ( .IN1(WX853), .IN2(WX789), .IN3(WX725), .Q(n3512) );
  XNOR3X1 U4363 ( .IN1(n3514), .IN2(n4756), .IN3(n3515), .Q(n2577) );
  XNOR3X1 U4364 ( .IN1(WX851), .IN2(WX787), .IN3(test_so4), .Q(n3514) );
  XNOR3X1 U4365 ( .IN1(n3516), .IN2(n4756), .IN3(n3517), .Q(n2580) );
  XNOR3X1 U4366 ( .IN1(WX849), .IN2(WX785), .IN3(WX721), .Q(n3516) );
  XNOR3X1 U4367 ( .IN1(n3518), .IN2(n4757), .IN3(n3519), .Q(n2583) );
  XNOR3X1 U4368 ( .IN1(WX847), .IN2(WX783), .IN3(WX719), .Q(n3518) );
  XNOR3X1 U4369 ( .IN1(n3520), .IN2(n4757), .IN3(n3521), .Q(n2586) );
  XNOR3X1 U4370 ( .IN1(WX845), .IN2(WX781), .IN3(WX717), .Q(n3520) );
  XNOR3X1 U4371 ( .IN1(n3522), .IN2(n4758), .IN3(n3523), .Q(n2589) );
  XNOR3X1 U4372 ( .IN1(WX843), .IN2(WX779), .IN3(WX715), .Q(n3522) );
  XNOR3X1 U4373 ( .IN1(n3524), .IN2(n4759), .IN3(n3525), .Q(n2602) );
  XNOR3X1 U4374 ( .IN1(WX841), .IN2(WX777), .IN3(WX713), .Q(n3524) );
  XNOR3X1 U4375 ( .IN1(n3526), .IN2(n4759), .IN3(n3527), .Q(n2615) );
  XNOR3X1 U4376 ( .IN1(WX839), .IN2(WX775), .IN3(WX711), .Q(n3526) );
  XNOR3X1 U4377 ( .IN1(n3528), .IN2(n4760), .IN3(n3529), .Q(n2630) );
  XNOR3X1 U4378 ( .IN1(WX837), .IN2(WX773), .IN3(WX709), .Q(n3528) );
  AO221X1 U4379 ( .IN1(WX10888), .IN2(n4473), .IN3(n4311), .IN4(n2154), .IN5(
        n3213), .Q(WX11050) );
  AO22X1 U4380 ( .IN1(n4171), .IN2(CRC_OUT_1_0), .IN3(DATA_0_0), .IN4(n4040), 
        .Q(n3213) );
  AO221X1 U4381 ( .IN1(WX10886), .IN2(n4473), .IN3(n4311), .IN4(n2157), .IN5(
        n3215), .Q(WX11048) );
  AO22X1 U4382 ( .IN1(n4171), .IN2(CRC_OUT_1_1), .IN3(DATA_0_1), .IN4(n4041), 
        .Q(n3215) );
  AO221X1 U4383 ( .IN1(WX10884), .IN2(n4474), .IN3(n4312), .IN4(n2160), .IN5(
        n3217), .Q(WX11046) );
  AO22X1 U4384 ( .IN1(n4172), .IN2(CRC_OUT_1_2), .IN3(DATA_0_2), .IN4(n4040), 
        .Q(n3217) );
  AO221X1 U4385 ( .IN1(WX10882), .IN2(n4474), .IN3(n4312), .IN4(n2163), .IN5(
        n3219), .Q(WX11044) );
  AO22X1 U4386 ( .IN1(n4172), .IN2(CRC_OUT_1_3), .IN3(DATA_0_3), .IN4(n4040), 
        .Q(n3219) );
  AO221X1 U4387 ( .IN1(WX10880), .IN2(n4474), .IN3(n4312), .IN4(n2166), .IN5(
        n3221), .Q(WX11042) );
  AO22X1 U4388 ( .IN1(n4172), .IN2(CRC_OUT_1_4), .IN3(DATA_0_4), .IN4(n4041), 
        .Q(n3221) );
  AO221X1 U4389 ( .IN1(WX10878), .IN2(n4474), .IN3(n4312), .IN4(n2169), .IN5(
        n3223), .Q(WX11040) );
  AO22X1 U4390 ( .IN1(n4172), .IN2(CRC_OUT_1_5), .IN3(DATA_0_5), .IN4(n4041), 
        .Q(n3223) );
  AO221X1 U4391 ( .IN1(WX10876), .IN2(n4474), .IN3(n4313), .IN4(n2172), .IN5(
        n3225), .Q(WX11038) );
  AO22X1 U4392 ( .IN1(n4173), .IN2(CRC_OUT_1_6), .IN3(DATA_0_6), .IN4(n4039), 
        .Q(n3225) );
  AO221X1 U4393 ( .IN1(WX10874), .IN2(n4475), .IN3(n4313), .IN4(n2175), .IN5(
        n3227), .Q(WX11036) );
  AO22X1 U4394 ( .IN1(n4173), .IN2(CRC_OUT_1_7), .IN3(DATA_0_7), .IN4(n4041), 
        .Q(n3227) );
  AO221X1 U4395 ( .IN1(WX10872), .IN2(n4475), .IN3(n4313), .IN4(n2178), .IN5(
        n3229), .Q(WX11034) );
  AO22X1 U4396 ( .IN1(n4173), .IN2(CRC_OUT_1_8), .IN3(DATA_0_8), .IN4(n4039), 
        .Q(n3229) );
  AO221X1 U4397 ( .IN1(WX10870), .IN2(n4475), .IN3(n4313), .IN4(n2181), .IN5(
        n3231), .Q(WX11032) );
  AO22X1 U4398 ( .IN1(n4173), .IN2(CRC_OUT_1_9), .IN3(DATA_0_9), .IN4(n4039), 
        .Q(n3231) );
  AO221X1 U4399 ( .IN1(WX10868), .IN2(n4475), .IN3(n4314), .IN4(n2184), .IN5(
        n3233), .Q(WX11030) );
  AO22X1 U4400 ( .IN1(n4174), .IN2(CRC_OUT_1_10), .IN3(DATA_0_10), .IN4(n4040), 
        .Q(n3233) );
  AO221X1 U4401 ( .IN1(WX10866), .IN2(n4475), .IN3(n4314), .IN4(n2187), .IN5(
        n3235), .Q(WX11028) );
  AO22X1 U4402 ( .IN1(n4174), .IN2(CRC_OUT_1_11), .IN3(DATA_0_11), .IN4(n4038), 
        .Q(n3235) );
  AO221X1 U4403 ( .IN1(WX10864), .IN2(n4476), .IN3(n4314), .IN4(n2190), .IN5(
        n3237), .Q(WX11026) );
  AO22X1 U4404 ( .IN1(n4174), .IN2(CRC_OUT_1_12), .IN3(DATA_0_12), .IN4(n4038), 
        .Q(n3237) );
  AO221X1 U4405 ( .IN1(WX10862), .IN2(n4476), .IN3(n4314), .IN4(n2193), .IN5(
        n3239), .Q(WX11024) );
  AO22X1 U4406 ( .IN1(n4174), .IN2(CRC_OUT_1_13), .IN3(DATA_0_13), .IN4(n4037), 
        .Q(n3239) );
  AO221X1 U4407 ( .IN1(WX10860), .IN2(n4476), .IN3(n4315), .IN4(n2196), .IN5(
        n3241), .Q(WX11022) );
  AO22X1 U4408 ( .IN1(n4175), .IN2(CRC_OUT_1_14), .IN3(DATA_0_14), .IN4(n4038), 
        .Q(n3241) );
  AO221X1 U4409 ( .IN1(WX10858), .IN2(n4476), .IN3(n4315), .IN4(n2199), .IN5(
        n3243), .Q(WX11020) );
  AO22X1 U4410 ( .IN1(n4175), .IN2(CRC_OUT_1_15), .IN3(DATA_0_15), .IN4(n4037), 
        .Q(n3243) );
  AO221X1 U4411 ( .IN1(WX10856), .IN2(n4476), .IN3(n4315), .IN4(n2202), .IN5(
        n3245), .Q(WX11018) );
  AO22X1 U4412 ( .IN1(n4175), .IN2(CRC_OUT_1_16), .IN3(DATA_0_16), .IN4(n4040), 
        .Q(n3245) );
  AO221X1 U4413 ( .IN1(WX10854), .IN2(n4477), .IN3(n4315), .IN4(n2205), .IN5(
        n3247), .Q(WX11016) );
  AO22X1 U4414 ( .IN1(n4175), .IN2(CRC_OUT_1_17), .IN3(DATA_0_17), .IN4(n4037), 
        .Q(n3247) );
  AO221X1 U4415 ( .IN1(WX10852), .IN2(n4477), .IN3(n4316), .IN4(n2208), .IN5(
        n3249), .Q(WX11014) );
  AO22X1 U4416 ( .IN1(n4176), .IN2(CRC_OUT_1_18), .IN3(DATA_0_18), .IN4(n4037), 
        .Q(n3249) );
  AO221X1 U4417 ( .IN1(WX10850), .IN2(n4477), .IN3(n4316), .IN4(n2211), .IN5(
        n3251), .Q(WX11012) );
  AO22X1 U4418 ( .IN1(n4176), .IN2(CRC_OUT_1_19), .IN3(DATA_0_19), .IN4(n4039), 
        .Q(n3251) );
  AO221X1 U4419 ( .IN1(WX10848), .IN2(n4477), .IN3(n4316), .IN4(n2214), .IN5(
        n3253), .Q(WX11010) );
  AO22X1 U4420 ( .IN1(n4176), .IN2(CRC_OUT_1_20), .IN3(DATA_0_20), .IN4(n4036), 
        .Q(n3253) );
  AO221X1 U4421 ( .IN1(WX10846), .IN2(n4477), .IN3(n4316), .IN4(n2217), .IN5(
        n3257), .Q(WX11008) );
  AO22X1 U4422 ( .IN1(n4176), .IN2(CRC_OUT_1_21), .IN3(DATA_0_21), .IN4(n4041), 
        .Q(n3257) );
  AO221X1 U4423 ( .IN1(WX10844), .IN2(n4478), .IN3(n4317), .IN4(n2220), .IN5(
        n3259), .Q(WX11006) );
  AO22X1 U4424 ( .IN1(n4177), .IN2(CRC_OUT_1_22), .IN3(DATA_0_22), .IN4(n4038), 
        .Q(n3259) );
  AO221X1 U4425 ( .IN1(WX10842), .IN2(n4478), .IN3(n4317), .IN4(n2223), .IN5(
        n3261), .Q(WX11004) );
  AO22X1 U4426 ( .IN1(n4177), .IN2(CRC_OUT_1_23), .IN3(DATA_0_23), .IN4(n4036), 
        .Q(n3261) );
  AO221X1 U4427 ( .IN1(WX10840), .IN2(n4478), .IN3(n4317), .IN4(n2226), .IN5(
        n3263), .Q(WX11002) );
  AO22X1 U4428 ( .IN1(n4177), .IN2(CRC_OUT_1_24), .IN3(DATA_0_24), .IN4(n4036), 
        .Q(n3263) );
  AO221X1 U4429 ( .IN1(WX10838), .IN2(n4478), .IN3(n4317), .IN4(n2229), .IN5(
        n3265), .Q(WX11000) );
  AO22X1 U4430 ( .IN1(n4177), .IN2(CRC_OUT_1_25), .IN3(DATA_0_25), .IN4(n4038), 
        .Q(n3265) );
  AO221X1 U4431 ( .IN1(WX10836), .IN2(n4478), .IN3(n4318), .IN4(n2232), .IN5(
        n3267), .Q(WX10998) );
  AO22X1 U4432 ( .IN1(n4178), .IN2(CRC_OUT_1_26), .IN3(DATA_0_26), .IN4(n4036), 
        .Q(n3267) );
  AO221X1 U4433 ( .IN1(WX10834), .IN2(n4479), .IN3(n4318), .IN4(n2235), .IN5(
        n3269), .Q(WX10996) );
  AO22X1 U4434 ( .IN1(n4178), .IN2(CRC_OUT_1_27), .IN3(DATA_0_27), .IN4(n4036), 
        .Q(n3269) );
  AO221X1 U4435 ( .IN1(WX10832), .IN2(n4479), .IN3(n4318), .IN4(n2238), .IN5(
        n3271), .Q(WX10994) );
  AO22X1 U4436 ( .IN1(n4178), .IN2(CRC_OUT_1_28), .IN3(DATA_0_28), .IN4(n4037), 
        .Q(n3271) );
  AO221X1 U4437 ( .IN1(WX10830), .IN2(n4479), .IN3(n4318), .IN4(n2241), .IN5(
        n3273), .Q(WX10992) );
  AO22X1 U4438 ( .IN1(n4178), .IN2(CRC_OUT_1_29), .IN3(DATA_0_29), .IN4(n4039), 
        .Q(n3273) );
  AO221X1 U4439 ( .IN1(WX10828), .IN2(n4479), .IN3(n4319), .IN4(n2244), .IN5(
        n3275), .Q(WX10990) );
  AO22X1 U4440 ( .IN1(n4179), .IN2(CRC_OUT_1_30), .IN3(DATA_0_30), .IN4(n4035), 
        .Q(n3275) );
  AO221X1 U4441 ( .IN1(WX9595), .IN2(n4424), .IN3(n4284), .IN4(n2150), .IN5(
        n2151), .Q(WX9757) );
  AO22X1 U4442 ( .IN1(n4144), .IN2(CRC_OUT_2_0), .IN3(n4044), .IN4(n2154), .Q(
        n2151) );
  AO221X1 U4443 ( .IN1(WX9593), .IN2(n4424), .IN3(n4337), .IN4(n2155), .IN5(
        n2156), .Q(WX9755) );
  AO22X1 U4444 ( .IN1(n4197), .IN2(CRC_OUT_2_1), .IN3(n4077), .IN4(n2157), .Q(
        n2156) );
  AO221X1 U4445 ( .IN1(WX9591), .IN2(n4424), .IN3(n4319), .IN4(n2158), .IN5(
        n2159), .Q(WX9753) );
  AO22X1 U4446 ( .IN1(n4179), .IN2(CRC_OUT_2_2), .IN3(n4063), .IN4(n2160), .Q(
        n2159) );
  AO221X1 U4447 ( .IN1(WX9589), .IN2(n4424), .IN3(n4319), .IN4(n2161), .IN5(
        n2162), .Q(WX9751) );
  AO22X1 U4448 ( .IN1(n4179), .IN2(CRC_OUT_2_3), .IN3(n4063), .IN4(n2163), .Q(
        n2162) );
  AO221X1 U4449 ( .IN1(WX9587), .IN2(n4424), .IN3(n4320), .IN4(n2164), .IN5(
        n2165), .Q(WX9749) );
  AO22X1 U4450 ( .IN1(n4180), .IN2(CRC_OUT_2_4), .IN3(n4063), .IN4(n2166), .Q(
        n2165) );
  AO221X1 U4451 ( .IN1(WX9585), .IN2(n4425), .IN3(n4320), .IN4(n2167), .IN5(
        n2168), .Q(WX9747) );
  AO22X1 U4452 ( .IN1(n4180), .IN2(CRC_OUT_2_5), .IN3(n4064), .IN4(n2169), .Q(
        n2168) );
  AO221X1 U4453 ( .IN1(WX9583), .IN2(n4425), .IN3(n4320), .IN4(n2170), .IN5(
        n2171), .Q(WX9745) );
  AO22X1 U4454 ( .IN1(n4180), .IN2(CRC_OUT_2_6), .IN3(n4064), .IN4(n2172), .Q(
        n2171) );
  AO221X1 U4455 ( .IN1(WX9581), .IN2(n4425), .IN3(n4320), .IN4(n2173), .IN5(
        n2174), .Q(WX9743) );
  AO22X1 U4456 ( .IN1(n4180), .IN2(CRC_OUT_2_7), .IN3(n4064), .IN4(n2175), .Q(
        n2174) );
  AO221X1 U4457 ( .IN1(WX9579), .IN2(n4425), .IN3(n4321), .IN4(n2176), .IN5(
        n2177), .Q(WX9741) );
  AO22X1 U4458 ( .IN1(n4181), .IN2(CRC_OUT_2_8), .IN3(n4064), .IN4(n2178), .Q(
        n2177) );
  AO221X1 U4459 ( .IN1(WX9577), .IN2(n4425), .IN3(n4321), .IN4(n2179), .IN5(
        n2180), .Q(WX9739) );
  AO22X1 U4460 ( .IN1(n4181), .IN2(CRC_OUT_2_9), .IN3(n4064), .IN4(n2181), .Q(
        n2180) );
  AO221X1 U4461 ( .IN1(WX9575), .IN2(n4426), .IN3(n4321), .IN4(n2182), .IN5(
        n2183), .Q(WX9737) );
  AO22X1 U4462 ( .IN1(n4181), .IN2(CRC_OUT_2_10), .IN3(n4065), .IN4(n2184), 
        .Q(n2183) );
  AO221X1 U4463 ( .IN1(WX9573), .IN2(n4426), .IN3(n4321), .IN4(n2185), .IN5(
        n2186), .Q(WX9735) );
  AO22X1 U4464 ( .IN1(n4181), .IN2(CRC_OUT_2_11), .IN3(n4065), .IN4(n2187), 
        .Q(n2186) );
  AO221X1 U4465 ( .IN1(WX9571), .IN2(n4426), .IN3(n4322), .IN4(n2188), .IN5(
        n2189), .Q(WX9733) );
  AO22X1 U4466 ( .IN1(n4182), .IN2(CRC_OUT_2_12), .IN3(n4065), .IN4(n2190), 
        .Q(n2189) );
  AO221X1 U4467 ( .IN1(WX9569), .IN2(n4426), .IN3(n4322), .IN4(n2191), .IN5(
        n2192), .Q(WX9731) );
  AO22X1 U4468 ( .IN1(n4182), .IN2(CRC_OUT_2_13), .IN3(n4065), .IN4(n2193), 
        .Q(n2192) );
  AO221X1 U4469 ( .IN1(WX9567), .IN2(n4426), .IN3(n4322), .IN4(n2194), .IN5(
        n2195), .Q(WX9729) );
  AO22X1 U4470 ( .IN1(n4182), .IN2(CRC_OUT_2_14), .IN3(n4065), .IN4(n2196), 
        .Q(n2195) );
  AO221X1 U4471 ( .IN1(WX9565), .IN2(n4427), .IN3(n4322), .IN4(n2197), .IN5(
        n2198), .Q(WX9727) );
  AO22X1 U4472 ( .IN1(n4182), .IN2(CRC_OUT_2_15), .IN3(n4066), .IN4(n2199), 
        .Q(n2198) );
  AO221X1 U4473 ( .IN1(WX9563), .IN2(n4427), .IN3(n4323), .IN4(n2200), .IN5(
        n2201), .Q(WX9725) );
  AO22X1 U4474 ( .IN1(n4183), .IN2(CRC_OUT_2_16), .IN3(n4066), .IN4(n2202), 
        .Q(n2201) );
  AO221X1 U4475 ( .IN1(WX9561), .IN2(n4427), .IN3(n4323), .IN4(n2203), .IN5(
        n2204), .Q(WX9723) );
  AO22X1 U4476 ( .IN1(n4183), .IN2(CRC_OUT_2_17), .IN3(n4066), .IN4(n2205), 
        .Q(n2204) );
  AO221X1 U4477 ( .IN1(WX9559), .IN2(n4427), .IN3(n4323), .IN4(n2206), .IN5(
        n2207), .Q(WX9721) );
  AO22X1 U4478 ( .IN1(n4183), .IN2(CRC_OUT_2_18), .IN3(n4066), .IN4(n2208), 
        .Q(n2207) );
  AO221X1 U4479 ( .IN1(WX9557), .IN2(n4427), .IN3(n4323), .IN4(n2209), .IN5(
        n2210), .Q(WX9719) );
  AO22X1 U4480 ( .IN1(n4183), .IN2(CRC_OUT_2_19), .IN3(n4066), .IN4(n2211), 
        .Q(n2210) );
  AO221X1 U4481 ( .IN1(WX9555), .IN2(n4428), .IN3(n4324), .IN4(n2212), .IN5(
        n2213), .Q(WX9717) );
  AO22X1 U4482 ( .IN1(n4184), .IN2(CRC_OUT_2_20), .IN3(n4067), .IN4(n2214), 
        .Q(n2213) );
  AO221X1 U4483 ( .IN1(WX9553), .IN2(n4428), .IN3(n4324), .IN4(n2215), .IN5(
        n2216), .Q(WX9715) );
  AO22X1 U4484 ( .IN1(n4184), .IN2(CRC_OUT_2_21), .IN3(n4067), .IN4(n2217), 
        .Q(n2216) );
  AO221X1 U4485 ( .IN1(WX9551), .IN2(n4428), .IN3(n4324), .IN4(n2218), .IN5(
        n2219), .Q(WX9713) );
  AO22X1 U4486 ( .IN1(n4184), .IN2(CRC_OUT_2_22), .IN3(n4067), .IN4(n2220), 
        .Q(n2219) );
  AO221X1 U4487 ( .IN1(WX9549), .IN2(n4428), .IN3(n4324), .IN4(n2221), .IN5(
        n2222), .Q(WX9711) );
  AO22X1 U4488 ( .IN1(n4184), .IN2(CRC_OUT_2_23), .IN3(n4067), .IN4(n2223), 
        .Q(n2222) );
  AO221X1 U4489 ( .IN1(WX9547), .IN2(n4428), .IN3(n4325), .IN4(n2224), .IN5(
        n2225), .Q(WX9709) );
  AO22X1 U4490 ( .IN1(n4185), .IN2(CRC_OUT_2_24), .IN3(n4067), .IN4(n2226), 
        .Q(n2225) );
  AO221X1 U4491 ( .IN1(WX9545), .IN2(n4429), .IN3(n4325), .IN4(n2227), .IN5(
        n2228), .Q(WX9707) );
  AO22X1 U4492 ( .IN1(n4185), .IN2(CRC_OUT_2_25), .IN3(n4068), .IN4(n2229), 
        .Q(n2228) );
  AO221X1 U4493 ( .IN1(WX9543), .IN2(n4429), .IN3(n4325), .IN4(n2230), .IN5(
        n2231), .Q(WX9705) );
  AO22X1 U4494 ( .IN1(n4185), .IN2(CRC_OUT_2_26), .IN3(n4068), .IN4(n2232), 
        .Q(n2231) );
  AO221X1 U4495 ( .IN1(WX9541), .IN2(n4429), .IN3(n4325), .IN4(n2233), .IN5(
        n2234), .Q(WX9703) );
  AO22X1 U4496 ( .IN1(n4185), .IN2(CRC_OUT_2_27), .IN3(n4068), .IN4(n2235), 
        .Q(n2234) );
  AO221X1 U4497 ( .IN1(WX9539), .IN2(n4429), .IN3(n4326), .IN4(n2236), .IN5(
        n2237), .Q(WX9701) );
  AO22X1 U4498 ( .IN1(n4186), .IN2(CRC_OUT_2_28), .IN3(n4068), .IN4(n2238), 
        .Q(n2237) );
  AO221X1 U4499 ( .IN1(WX9537), .IN2(n4429), .IN3(n4326), .IN4(n2239), .IN5(
        n2240), .Q(WX9699) );
  AO22X1 U4500 ( .IN1(n4186), .IN2(CRC_OUT_2_29), .IN3(n4068), .IN4(n2241), 
        .Q(n2240) );
  AO221X1 U4501 ( .IN1(WX9535), .IN2(n4430), .IN3(n4326), .IN4(n2242), .IN5(
        n2243), .Q(WX9697) );
  AO22X1 U4502 ( .IN1(n4186), .IN2(CRC_OUT_2_30), .IN3(n4069), .IN4(n2244), 
        .Q(n2243) );
  AO221X1 U4503 ( .IN1(WX9536), .IN2(n2245), .IN3(n4035), .IN4(n2246), .IN5(
        n2247), .Q(WX9695) );
  AO22X1 U4504 ( .IN1(n4355), .IN2(n2248), .IN3(n4215), .IN4(CRC_OUT_2_31), 
        .Q(n2247) );
  AO221X1 U4505 ( .IN1(WX8302), .IN2(n4430), .IN3(n4326), .IN4(n2281), .IN5(
        n2282), .Q(WX8464) );
  AO22X1 U4506 ( .IN1(n4186), .IN2(CRC_OUT_3_0), .IN3(n4069), .IN4(n2150), .Q(
        n2282) );
  AO221X1 U4507 ( .IN1(WX8300), .IN2(n4430), .IN3(n4327), .IN4(n2284), .IN5(
        n2285), .Q(WX8462) );
  AO22X1 U4508 ( .IN1(n4187), .IN2(CRC_OUT_3_1), .IN3(n4069), .IN4(n2155), .Q(
        n2285) );
  AO221X1 U4509 ( .IN1(WX8298), .IN2(n4430), .IN3(n4327), .IN4(n2287), .IN5(
        n2288), .Q(WX8460) );
  AO22X1 U4510 ( .IN1(n4187), .IN2(CRC_OUT_3_2), .IN3(n4069), .IN4(n2158), .Q(
        n2288) );
  AO221X1 U4511 ( .IN1(WX8296), .IN2(n4430), .IN3(n4327), .IN4(n2290), .IN5(
        n2291), .Q(WX8458) );
  AO22X1 U4512 ( .IN1(n4187), .IN2(CRC_OUT_3_3), .IN3(n4069), .IN4(n2161), .Q(
        n2291) );
  AO221X1 U4513 ( .IN1(WX8294), .IN2(n4431), .IN3(n4327), .IN4(n2293), .IN5(
        n2294), .Q(WX8456) );
  AO22X1 U4514 ( .IN1(n4187), .IN2(CRC_OUT_3_4), .IN3(n4070), .IN4(n2164), .Q(
        n2294) );
  AO221X1 U4515 ( .IN1(WX8292), .IN2(n4431), .IN3(n4328), .IN4(n2296), .IN5(
        n2297), .Q(WX8454) );
  AO22X1 U4516 ( .IN1(n4188), .IN2(CRC_OUT_3_5), .IN3(n4070), .IN4(n2167), .Q(
        n2297) );
  AO221X1 U4517 ( .IN1(WX8290), .IN2(n4431), .IN3(n4328), .IN4(n2299), .IN5(
        n2300), .Q(WX8452) );
  AO22X1 U4518 ( .IN1(n4188), .IN2(CRC_OUT_3_6), .IN3(n4070), .IN4(n2170), .Q(
        n2300) );
  AO221X1 U4519 ( .IN1(WX8288), .IN2(n4431), .IN3(n4328), .IN4(n2302), .IN5(
        n2303), .Q(WX8450) );
  AO22X1 U4520 ( .IN1(n4188), .IN2(CRC_OUT_3_7), .IN3(n4070), .IN4(n2173), .Q(
        n2303) );
  AO221X1 U4521 ( .IN1(WX8286), .IN2(n4431), .IN3(n4328), .IN4(n2305), .IN5(
        n2306), .Q(WX8448) );
  AO22X1 U4522 ( .IN1(n4188), .IN2(CRC_OUT_3_8), .IN3(n4070), .IN4(n2176), .Q(
        n2306) );
  AO221X1 U4523 ( .IN1(WX8284), .IN2(n4432), .IN3(n4329), .IN4(n2308), .IN5(
        n2309), .Q(WX8446) );
  AO22X1 U4524 ( .IN1(n4189), .IN2(CRC_OUT_3_9), .IN3(n4071), .IN4(n2179), .Q(
        n2309) );
  AO221X1 U4525 ( .IN1(WX8282), .IN2(n4432), .IN3(n4329), .IN4(n2311), .IN5(
        n2312), .Q(WX8444) );
  AO22X1 U4526 ( .IN1(n4189), .IN2(CRC_OUT_3_10), .IN3(n4071), .IN4(n2182), 
        .Q(n2312) );
  AO221X1 U4527 ( .IN1(WX8280), .IN2(n4432), .IN3(n4329), .IN4(n2314), .IN5(
        n2315), .Q(WX8442) );
  AO22X1 U4528 ( .IN1(n4189), .IN2(CRC_OUT_3_11), .IN3(n4071), .IN4(n2185), 
        .Q(n2315) );
  AO221X1 U4529 ( .IN1(WX8278), .IN2(n4432), .IN3(n4329), .IN4(n2317), .IN5(
        n2318), .Q(WX8440) );
  AO22X1 U4530 ( .IN1(n4189), .IN2(CRC_OUT_3_12), .IN3(n4071), .IN4(n2188), 
        .Q(n2318) );
  AO221X1 U4531 ( .IN1(WX8276), .IN2(n4432), .IN3(n4330), .IN4(n2320), .IN5(
        n2321), .Q(WX8438) );
  AO22X1 U4532 ( .IN1(n4190), .IN2(CRC_OUT_3_13), .IN3(n4071), .IN4(n2191), 
        .Q(n2321) );
  AO221X1 U4533 ( .IN1(WX8274), .IN2(n4433), .IN3(n4330), .IN4(n2323), .IN5(
        n2324), .Q(WX8436) );
  AO22X1 U4534 ( .IN1(n4190), .IN2(CRC_OUT_3_14), .IN3(n4072), .IN4(n2194), 
        .Q(n2324) );
  AO221X1 U4535 ( .IN1(WX8272), .IN2(n4433), .IN3(n4330), .IN4(n2326), .IN5(
        n2327), .Q(WX8434) );
  AO22X1 U4536 ( .IN1(n4190), .IN2(CRC_OUT_3_15), .IN3(n4072), .IN4(n2197), 
        .Q(n2327) );
  AO221X1 U4537 ( .IN1(WX8270), .IN2(n4433), .IN3(n4330), .IN4(n2329), .IN5(
        n2330), .Q(WX8432) );
  AO22X1 U4538 ( .IN1(n4190), .IN2(CRC_OUT_3_16), .IN3(n4072), .IN4(n2200), 
        .Q(n2330) );
  AO221X1 U4539 ( .IN1(WX8268), .IN2(n4433), .IN3(n4331), .IN4(n2332), .IN5(
        n2333), .Q(WX8430) );
  AO22X1 U4540 ( .IN1(n4191), .IN2(CRC_OUT_3_17), .IN3(n4072), .IN4(n2203), 
        .Q(n2333) );
  AO221X1 U4541 ( .IN1(WX8266), .IN2(n4433), .IN3(n4331), .IN4(n2335), .IN5(
        n2336), .Q(WX8428) );
  AO22X1 U4542 ( .IN1(n4191), .IN2(CRC_OUT_3_18), .IN3(n4072), .IN4(n2206), 
        .Q(n2336) );
  AO221X1 U4543 ( .IN1(WX8264), .IN2(n4434), .IN3(n4331), .IN4(n2338), .IN5(
        n2339), .Q(WX8426) );
  AO22X1 U4544 ( .IN1(n4191), .IN2(CRC_OUT_3_19), .IN3(n4073), .IN4(n2209), 
        .Q(n2339) );
  AO221X1 U4545 ( .IN1(WX8262), .IN2(n4434), .IN3(n4331), .IN4(n2341), .IN5(
        n2342), .Q(WX8424) );
  AO22X1 U4546 ( .IN1(n4191), .IN2(CRC_OUT_3_20), .IN3(n4073), .IN4(n2212), 
        .Q(n2342) );
  AO221X1 U4547 ( .IN1(WX8260), .IN2(n4434), .IN3(n4332), .IN4(n2344), .IN5(
        n2345), .Q(WX8422) );
  AO22X1 U4548 ( .IN1(n4192), .IN2(CRC_OUT_3_21), .IN3(n4073), .IN4(n2215), 
        .Q(n2345) );
  AO221X1 U4549 ( .IN1(WX8258), .IN2(n4434), .IN3(n4332), .IN4(n2347), .IN5(
        n2348), .Q(WX8420) );
  AO22X1 U4550 ( .IN1(n4192), .IN2(CRC_OUT_3_22), .IN3(n4073), .IN4(n2218), 
        .Q(n2348) );
  AO221X1 U4551 ( .IN1(WX8256), .IN2(n4434), .IN3(n4332), .IN4(n2350), .IN5(
        n2351), .Q(WX8418) );
  AO22X1 U4552 ( .IN1(n4192), .IN2(CRC_OUT_3_23), .IN3(n4073), .IN4(n2221), 
        .Q(n2351) );
  AO221X1 U4553 ( .IN1(WX8254), .IN2(n4435), .IN3(n4332), .IN4(n2353), .IN5(
        n2354), .Q(WX8416) );
  AO22X1 U4554 ( .IN1(n4192), .IN2(CRC_OUT_3_24), .IN3(n4074), .IN4(n2224), 
        .Q(n2354) );
  AO221X1 U4555 ( .IN1(WX8252), .IN2(n4435), .IN3(n4333), .IN4(n2356), .IN5(
        n2357), .Q(WX8414) );
  AO22X1 U4556 ( .IN1(n4193), .IN2(CRC_OUT_3_25), .IN3(n4074), .IN4(n2227), 
        .Q(n2357) );
  AO221X1 U4557 ( .IN1(WX8250), .IN2(n4435), .IN3(n4333), .IN4(n2359), .IN5(
        n2360), .Q(WX8412) );
  AO22X1 U4558 ( .IN1(n4193), .IN2(CRC_OUT_3_26), .IN3(n4074), .IN4(n2230), 
        .Q(n2360) );
  AO221X1 U4559 ( .IN1(WX8248), .IN2(n4435), .IN3(n4333), .IN4(n2362), .IN5(
        n2363), .Q(WX8410) );
  AO22X1 U4560 ( .IN1(n4193), .IN2(CRC_OUT_3_27), .IN3(n4074), .IN4(n2233), 
        .Q(n2363) );
  AO221X1 U4561 ( .IN1(WX8246), .IN2(n4435), .IN3(n4333), .IN4(n2365), .IN5(
        n2366), .Q(WX8408) );
  AO22X1 U4562 ( .IN1(n4193), .IN2(CRC_OUT_3_28), .IN3(n4074), .IN4(n2236), 
        .Q(n2366) );
  AO221X1 U4563 ( .IN1(WX8244), .IN2(n4436), .IN3(n4334), .IN4(n2368), .IN5(
        n2369), .Q(WX8406) );
  AO22X1 U4564 ( .IN1(n4194), .IN2(CRC_OUT_3_29), .IN3(n4075), .IN4(n2239), 
        .Q(n2369) );
  AO221X1 U4565 ( .IN1(WX8242), .IN2(n4436), .IN3(n4334), .IN4(n2371), .IN5(
        n2372), .Q(WX8404) );
  AO22X1 U4566 ( .IN1(n4194), .IN2(CRC_OUT_3_30), .IN3(n4075), .IN4(n2242), 
        .Q(n2372) );
  AO221X1 U4567 ( .IN1(WX8243), .IN2(n2245), .IN3(n4034), .IN4(n2248), .IN5(
        n2374), .Q(WX8402) );
  AO22X1 U4568 ( .IN1(n4353), .IN2(n2375), .IN3(n4213), .IN4(CRC_OUT_3_31), 
        .Q(n2374) );
  AO221X1 U4569 ( .IN1(WX7009), .IN2(n4436), .IN3(n4334), .IN4(n2409), .IN5(
        n2410), .Q(WX7171) );
  AO22X1 U4570 ( .IN1(n4194), .IN2(CRC_OUT_4_0), .IN3(n4075), .IN4(n2281), .Q(
        n2410) );
  AO221X1 U4571 ( .IN1(WX7007), .IN2(n4436), .IN3(n4334), .IN4(n2412), .IN5(
        n2413), .Q(WX7169) );
  AO22X1 U4572 ( .IN1(n4194), .IN2(CRC_OUT_4_1), .IN3(n4075), .IN4(n2284), .Q(
        n2413) );
  AO221X1 U4573 ( .IN1(WX7005), .IN2(n4436), .IN3(n4335), .IN4(n2415), .IN5(
        n2416), .Q(WX7167) );
  AO22X1 U4574 ( .IN1(n4195), .IN2(CRC_OUT_4_2), .IN3(n4075), .IN4(n2287), .Q(
        n2416) );
  AO221X1 U4575 ( .IN1(WX7003), .IN2(n4437), .IN3(n4335), .IN4(n2418), .IN5(
        n2419), .Q(WX7165) );
  AO22X1 U4576 ( .IN1(n4195), .IN2(CRC_OUT_4_3), .IN3(n4076), .IN4(n2290), .Q(
        n2419) );
  AO221X1 U4577 ( .IN1(WX7001), .IN2(n4437), .IN3(n4335), .IN4(n2421), .IN5(
        n2422), .Q(WX7163) );
  AO22X1 U4578 ( .IN1(n4195), .IN2(CRC_OUT_4_4), .IN3(n4076), .IN4(n2293), .Q(
        n2422) );
  AO221X1 U4579 ( .IN1(WX6999), .IN2(n4437), .IN3(n4335), .IN4(n2424), .IN5(
        n2425), .Q(WX7161) );
  AO22X1 U4580 ( .IN1(n4195), .IN2(CRC_OUT_4_5), .IN3(n4076), .IN4(n2296), .Q(
        n2425) );
  AO221X1 U4581 ( .IN1(WX6997), .IN2(n4437), .IN3(n4336), .IN4(n2427), .IN5(
        n2428), .Q(WX7159) );
  AO22X1 U4582 ( .IN1(n4196), .IN2(CRC_OUT_4_6), .IN3(n4076), .IN4(n2299), .Q(
        n2428) );
  AO221X1 U4583 ( .IN1(WX6995), .IN2(n4437), .IN3(n4336), .IN4(n2430), .IN5(
        n2431), .Q(WX7157) );
  AO22X1 U4584 ( .IN1(n4196), .IN2(CRC_OUT_4_7), .IN3(n4076), .IN4(n2302), .Q(
        n2431) );
  AO221X1 U4585 ( .IN1(WX6993), .IN2(n4438), .IN3(n4336), .IN4(n2433), .IN5(
        n2434), .Q(WX7155) );
  AO22X1 U4586 ( .IN1(n4196), .IN2(CRC_OUT_4_8), .IN3(n4077), .IN4(n2305), .Q(
        n2434) );
  AO221X1 U4587 ( .IN1(WX6991), .IN2(n4438), .IN3(n4336), .IN4(n2436), .IN5(
        n2437), .Q(WX7153) );
  AO22X1 U4588 ( .IN1(n4196), .IN2(CRC_OUT_4_9), .IN3(n4077), .IN4(n2308), .Q(
        n2437) );
  AO221X1 U4589 ( .IN1(WX6989), .IN2(n4438), .IN3(n4337), .IN4(n2439), .IN5(
        n2440), .Q(WX7151) );
  AO22X1 U4590 ( .IN1(n4197), .IN2(CRC_OUT_4_10), .IN3(n4077), .IN4(n2311), 
        .Q(n2440) );
  AO221X1 U4591 ( .IN1(WX6987), .IN2(n4438), .IN3(n4337), .IN4(n2442), .IN5(
        n2443), .Q(WX7149) );
  AO22X1 U4592 ( .IN1(n4197), .IN2(CRC_OUT_4_11), .IN3(n4077), .IN4(n2314), 
        .Q(n2443) );
  AO221X1 U4593 ( .IN1(WX6985), .IN2(n4438), .IN3(n4338), .IN4(n2445), .IN5(
        n2446), .Q(WX7147) );
  AO22X1 U4594 ( .IN1(n4198), .IN2(CRC_OUT_4_12), .IN3(n4078), .IN4(n2317), 
        .Q(n2446) );
  AO221X1 U4595 ( .IN1(WX6983), .IN2(n4439), .IN3(n4338), .IN4(n2448), .IN5(
        n2449), .Q(WX7145) );
  AO22X1 U4596 ( .IN1(n4198), .IN2(CRC_OUT_4_13), .IN3(n4078), .IN4(n2320), 
        .Q(n2449) );
  AO221X1 U4597 ( .IN1(WX6981), .IN2(n4439), .IN3(n4338), .IN4(n2451), .IN5(
        n2452), .Q(WX7143) );
  AO22X1 U4598 ( .IN1(n4198), .IN2(CRC_OUT_4_14), .IN3(n4078), .IN4(n2323), 
        .Q(n2452) );
  AO221X1 U4599 ( .IN1(WX6979), .IN2(n4439), .IN3(n4338), .IN4(n2454), .IN5(
        n2455), .Q(WX7141) );
  AO22X1 U4600 ( .IN1(n4198), .IN2(CRC_OUT_4_15), .IN3(n4078), .IN4(n2326), 
        .Q(n2455) );
  AO221X1 U4601 ( .IN1(WX6977), .IN2(n4439), .IN3(n4339), .IN4(n2457), .IN5(
        n2458), .Q(WX7139) );
  AO22X1 U4602 ( .IN1(n4199), .IN2(CRC_OUT_4_16), .IN3(n4078), .IN4(n2329), 
        .Q(n2458) );
  AO221X1 U4603 ( .IN1(WX6975), .IN2(n4439), .IN3(n4337), .IN4(n2460), .IN5(
        n2461), .Q(WX7137) );
  AO22X1 U4604 ( .IN1(n4197), .IN2(CRC_OUT_4_17), .IN3(n4079), .IN4(n2332), 
        .Q(n2461) );
  AO221X1 U4605 ( .IN1(WX6973), .IN2(n4440), .IN3(n4339), .IN4(n2463), .IN5(
        n2464), .Q(WX7135) );
  AO22X1 U4606 ( .IN1(n4199), .IN2(CRC_OUT_4_18), .IN3(n4079), .IN4(n2335), 
        .Q(n2464) );
  AO221X1 U4607 ( .IN1(WX6971), .IN2(n4440), .IN3(n4339), .IN4(n2466), .IN5(
        n2467), .Q(WX7133) );
  AO22X1 U4608 ( .IN1(n4199), .IN2(CRC_OUT_4_19), .IN3(n4079), .IN4(n2338), 
        .Q(n2467) );
  AO221X1 U4609 ( .IN1(WX6969), .IN2(n4440), .IN3(n4340), .IN4(n2469), .IN5(
        n2470), .Q(WX7131) );
  AO22X1 U4610 ( .IN1(n4200), .IN2(CRC_OUT_4_20), .IN3(n4079), .IN4(n2341), 
        .Q(n2470) );
  AO221X1 U4611 ( .IN1(WX6967), .IN2(n4440), .IN3(n4339), .IN4(n2472), .IN5(
        n2473), .Q(WX7129) );
  AO22X1 U4612 ( .IN1(n4199), .IN2(CRC_OUT_4_21), .IN3(n4079), .IN4(n2344), 
        .Q(n2473) );
  AO221X1 U4613 ( .IN1(WX6965), .IN2(n4440), .IN3(n4340), .IN4(n2475), .IN5(
        n2476), .Q(WX7127) );
  AO22X1 U4614 ( .IN1(n4200), .IN2(CRC_OUT_4_22), .IN3(n4080), .IN4(n2347), 
        .Q(n2476) );
  AO221X1 U4615 ( .IN1(WX6963), .IN2(n4441), .IN3(n4340), .IN4(n2478), .IN5(
        n2479), .Q(WX7125) );
  AO22X1 U4616 ( .IN1(n4200), .IN2(CRC_OUT_4_23), .IN3(n4080), .IN4(n2350), 
        .Q(n2479) );
  AO221X1 U4617 ( .IN1(WX6961), .IN2(n4441), .IN3(n4341), .IN4(n2481), .IN5(
        n2482), .Q(WX7123) );
  AO22X1 U4618 ( .IN1(n4201), .IN2(CRC_OUT_4_24), .IN3(n4080), .IN4(n2353), 
        .Q(n2482) );
  AO221X1 U4619 ( .IN1(WX6959), .IN2(n4441), .IN3(n4341), .IN4(n2484), .IN5(
        n2485), .Q(WX7121) );
  AO22X1 U4620 ( .IN1(n4201), .IN2(CRC_OUT_4_25), .IN3(n4080), .IN4(n2356), 
        .Q(n2485) );
  AO221X1 U4621 ( .IN1(WX6957), .IN2(n4441), .IN3(n4341), .IN4(n2487), .IN5(
        n2488), .Q(WX7119) );
  AO22X1 U4622 ( .IN1(n4201), .IN2(CRC_OUT_4_26), .IN3(n4080), .IN4(n2359), 
        .Q(n2488) );
  AO221X1 U4623 ( .IN1(WX6955), .IN2(n4441), .IN3(n4340), .IN4(n2490), .IN5(
        n2491), .Q(WX7117) );
  AO22X1 U4624 ( .IN1(n4200), .IN2(CRC_OUT_4_27), .IN3(n4081), .IN4(n2362), 
        .Q(n2491) );
  AO221X1 U4625 ( .IN1(WX6953), .IN2(n4442), .IN3(n4342), .IN4(n2493), .IN5(
        n2494), .Q(WX7115) );
  AO22X1 U4626 ( .IN1(n4202), .IN2(CRC_OUT_4_28), .IN3(n4081), .IN4(n2365), 
        .Q(n2494) );
  AO221X1 U4627 ( .IN1(WX6951), .IN2(n4442), .IN3(n4342), .IN4(n2496), .IN5(
        n2497), .Q(WX7113) );
  AO22X1 U4628 ( .IN1(n4202), .IN2(CRC_OUT_4_29), .IN3(n4081), .IN4(n2368), 
        .Q(n2497) );
  AO221X1 U4629 ( .IN1(WX6949), .IN2(n4442), .IN3(n4342), .IN4(n2499), .IN5(
        n2500), .Q(WX7111) );
  AO22X1 U4630 ( .IN1(n4202), .IN2(CRC_OUT_4_30), .IN3(n4081), .IN4(n2371), 
        .Q(n2500) );
  AO221X1 U4631 ( .IN1(WX6950), .IN2(n2245), .IN3(n4035), .IN4(n2375), .IN5(
        n2502), .Q(WX7109) );
  AO22X1 U4632 ( .IN1(n4354), .IN2(n2503), .IN3(n4214), .IN4(CRC_OUT_4_31), 
        .Q(n2502) );
  AO221X1 U4633 ( .IN1(WX5716), .IN2(n4448), .IN3(n4351), .IN4(n2633), .IN5(
        n2634), .Q(WX5878) );
  AO22X1 U4634 ( .IN1(n4211), .IN2(CRC_OUT_5_0), .IN3(n4088), .IN4(n2409), .Q(
        n2634) );
  AO221X1 U4635 ( .IN1(WX5714), .IN2(n4449), .IN3(n4349), .IN4(n2636), .IN5(
        n2637), .Q(WX5876) );
  AO22X1 U4636 ( .IN1(n4209), .IN2(CRC_OUT_5_1), .IN3(n4088), .IN4(n2412), .Q(
        n2637) );
  AO221X1 U4637 ( .IN1(WX5712), .IN2(n4449), .IN3(n4352), .IN4(n2639), .IN5(
        n2640), .Q(WX5874) );
  AO22X1 U4638 ( .IN1(n4212), .IN2(CRC_OUT_5_2), .IN3(n4088), .IN4(n2415), .Q(
        n2640) );
  AO221X1 U4639 ( .IN1(WX5710), .IN2(n4449), .IN3(n4350), .IN4(n2642), .IN5(
        n2643), .Q(WX5872) );
  AO22X1 U4640 ( .IN1(n4210), .IN2(CRC_OUT_5_3), .IN3(n4088), .IN4(n2418), .Q(
        n2643) );
  AO221X1 U4641 ( .IN1(WX5708), .IN2(n4449), .IN3(n4352), .IN4(n2645), .IN5(
        n2646), .Q(WX5870) );
  AO22X1 U4642 ( .IN1(n4212), .IN2(CRC_OUT_5_4), .IN3(n4088), .IN4(n2421), .Q(
        n2646) );
  AO221X1 U4643 ( .IN1(WX5706), .IN2(n4449), .IN3(n4351), .IN4(n2648), .IN5(
        n2649), .Q(WX5868) );
  AO22X1 U4644 ( .IN1(n4211), .IN2(CRC_OUT_5_5), .IN3(n4089), .IN4(n2424), .Q(
        n2649) );
  AO221X1 U4645 ( .IN1(WX5704), .IN2(n4450), .IN3(n4352), .IN4(n2651), .IN5(
        n2652), .Q(WX5866) );
  AO22X1 U4646 ( .IN1(n4212), .IN2(CRC_OUT_5_6), .IN3(n4089), .IN4(n2427), .Q(
        n2652) );
  AO221X1 U4647 ( .IN1(WX5702), .IN2(n4450), .IN3(n4350), .IN4(n2654), .IN5(
        n2655), .Q(WX5864) );
  AO22X1 U4648 ( .IN1(n4210), .IN2(CRC_OUT_5_7), .IN3(n4089), .IN4(n2430), .Q(
        n2655) );
  AO221X1 U4649 ( .IN1(WX5700), .IN2(n4450), .IN3(n4353), .IN4(n2657), .IN5(
        n2658), .Q(WX5862) );
  AO22X1 U4650 ( .IN1(n4213), .IN2(CRC_OUT_5_8), .IN3(n4089), .IN4(n2433), .Q(
        n2658) );
  AO221X1 U4651 ( .IN1(WX5698), .IN2(n4450), .IN3(n4351), .IN4(n2660), .IN5(
        n2661), .Q(WX5860) );
  AO22X1 U4652 ( .IN1(n4211), .IN2(CRC_OUT_5_9), .IN3(n4089), .IN4(n2436), .Q(
        n2661) );
  AO221X1 U4653 ( .IN1(WX5696), .IN2(n4450), .IN3(n4353), .IN4(n2663), .IN5(
        n2664), .Q(WX5858) );
  AO22X1 U4654 ( .IN1(n4213), .IN2(CRC_OUT_5_10), .IN3(n4090), .IN4(n2439), 
        .Q(n2664) );
  AO221X1 U4655 ( .IN1(WX5694), .IN2(n4451), .IN3(n4352), .IN4(n2666), .IN5(
        n2667), .Q(WX5856) );
  AO22X1 U4656 ( .IN1(n4212), .IN2(CRC_OUT_5_11), .IN3(n4090), .IN4(n2442), 
        .Q(n2667) );
  AO221X1 U4657 ( .IN1(WX5692), .IN2(n4451), .IN3(n4353), .IN4(n2669), .IN5(
        n2670), .Q(WX5854) );
  AO22X1 U4658 ( .IN1(n4213), .IN2(CRC_OUT_5_12), .IN3(n4090), .IN4(n2445), 
        .Q(n2670) );
  AO221X1 U4659 ( .IN1(WX5690), .IN2(n4451), .IN3(n4351), .IN4(n2672), .IN5(
        n2673), .Q(WX5852) );
  AO22X1 U4660 ( .IN1(n4211), .IN2(CRC_OUT_5_13), .IN3(n4090), .IN4(n2448), 
        .Q(n2673) );
  AO221X1 U4661 ( .IN1(WX5688), .IN2(n4451), .IN3(n4301), .IN4(n2675), .IN5(
        n2676), .Q(WX5850) );
  AO22X1 U4662 ( .IN1(n4161), .IN2(CRC_OUT_5_14), .IN3(n4090), .IN4(n2451), 
        .Q(n2676) );
  AO221X1 U4663 ( .IN1(WX5686), .IN2(n4451), .IN3(n4284), .IN4(n2678), .IN5(
        n2679), .Q(WX5848) );
  AO22X1 U4664 ( .IN1(n4144), .IN2(CRC_OUT_5_15), .IN3(n4091), .IN4(n2454), 
        .Q(n2679) );
  AO221X1 U4665 ( .IN1(WX5684), .IN2(n4452), .IN3(n4284), .IN4(n2681), .IN5(
        n2682), .Q(WX5846) );
  AO22X1 U4666 ( .IN1(n4144), .IN2(CRC_OUT_5_16), .IN3(n4091), .IN4(n2457), 
        .Q(n2682) );
  AO221X1 U4667 ( .IN1(WX5682), .IN2(n4452), .IN3(n4284), .IN4(n2684), .IN5(
        n2685), .Q(WX5844) );
  AO22X1 U4668 ( .IN1(n4144), .IN2(CRC_OUT_5_17), .IN3(n4091), .IN4(n2460), 
        .Q(n2685) );
  AO221X1 U4669 ( .IN1(WX5680), .IN2(n4452), .IN3(n4285), .IN4(n2687), .IN5(
        n2688), .Q(WX5842) );
  AO22X1 U4670 ( .IN1(n4145), .IN2(CRC_OUT_5_18), .IN3(n4052), .IN4(n2463), 
        .Q(n2688) );
  AO221X1 U4671 ( .IN1(WX5678), .IN2(n4452), .IN3(n4285), .IN4(n2690), .IN5(
        n2691), .Q(WX5840) );
  AO22X1 U4672 ( .IN1(n4145), .IN2(CRC_OUT_5_19), .IN3(n4045), .IN4(n2466), 
        .Q(n2691) );
  AO221X1 U4673 ( .IN1(WX5676), .IN2(n4452), .IN3(n4285), .IN4(n2693), .IN5(
        n2694), .Q(WX5838) );
  AO22X1 U4674 ( .IN1(n4145), .IN2(CRC_OUT_5_20), .IN3(n4042), .IN4(n2469), 
        .Q(n2694) );
  AO221X1 U4675 ( .IN1(WX5674), .IN2(n4453), .IN3(n4285), .IN4(n2696), .IN5(
        n2697), .Q(WX5836) );
  AO22X1 U4676 ( .IN1(n4145), .IN2(CRC_OUT_5_21), .IN3(n4043), .IN4(n2472), 
        .Q(n2697) );
  AO221X1 U4677 ( .IN1(WX5672), .IN2(n4453), .IN3(n4286), .IN4(n2699), .IN5(
        n2700), .Q(WX5834) );
  AO22X1 U4678 ( .IN1(n4146), .IN2(CRC_OUT_5_22), .IN3(n4042), .IN4(n2475), 
        .Q(n2700) );
  AO221X1 U4679 ( .IN1(WX5670), .IN2(n4453), .IN3(n4286), .IN4(n2702), .IN5(
        n2703), .Q(WX5832) );
  AO22X1 U4680 ( .IN1(n4146), .IN2(CRC_OUT_5_23), .IN3(n4042), .IN4(n2478), 
        .Q(n2703) );
  AO221X1 U4681 ( .IN1(WX5668), .IN2(n4453), .IN3(n4286), .IN4(n2705), .IN5(
        n2706), .Q(WX5830) );
  AO22X1 U4682 ( .IN1(n4146), .IN2(CRC_OUT_5_24), .IN3(n4043), .IN4(n2481), 
        .Q(n2706) );
  AO221X1 U4683 ( .IN1(WX5666), .IN2(n4453), .IN3(n4286), .IN4(n2708), .IN5(
        n2709), .Q(WX5828) );
  AO22X1 U4684 ( .IN1(n4146), .IN2(CRC_OUT_5_25), .IN3(n4042), .IN4(n2484), 
        .Q(n2709) );
  AO221X1 U4685 ( .IN1(WX5664), .IN2(n4454), .IN3(n4287), .IN4(n2711), .IN5(
        n2712), .Q(WX5826) );
  AO22X1 U4686 ( .IN1(n4147), .IN2(CRC_OUT_5_26), .IN3(n4042), .IN4(n2487), 
        .Q(n2712) );
  AO221X1 U4687 ( .IN1(WX5662), .IN2(n4454), .IN3(n4287), .IN4(n2714), .IN5(
        n2715), .Q(WX5824) );
  AO22X1 U4688 ( .IN1(n4147), .IN2(CRC_OUT_5_27), .IN3(n4047), .IN4(n2490), 
        .Q(n2715) );
  AO221X1 U4689 ( .IN1(WX5660), .IN2(n4454), .IN3(n4287), .IN4(n2717), .IN5(
        n2718), .Q(WX5822) );
  AO22X1 U4690 ( .IN1(n4147), .IN2(CRC_OUT_5_28), .IN3(n4043), .IN4(n2493), 
        .Q(n2718) );
  AO221X1 U4691 ( .IN1(WX5658), .IN2(n4454), .IN3(n4287), .IN4(n2720), .IN5(
        n2721), .Q(WX5820) );
  AO22X1 U4692 ( .IN1(n4147), .IN2(CRC_OUT_5_29), .IN3(n4043), .IN4(n2496), 
        .Q(n2721) );
  AO221X1 U4693 ( .IN1(WX5656), .IN2(n4454), .IN3(n4288), .IN4(n2723), .IN5(
        n2724), .Q(WX5818) );
  AO22X1 U4694 ( .IN1(n4148), .IN2(CRC_OUT_5_30), .IN3(n4044), .IN4(n2499), 
        .Q(n2724) );
  AO221X1 U4695 ( .IN1(WX5657), .IN2(n2245), .IN3(n4035), .IN4(n2503), .IN5(
        n2726), .Q(WX5816) );
  AO22X1 U4696 ( .IN1(n4354), .IN2(n2727), .IN3(n4214), .IN4(CRC_OUT_5_31), 
        .Q(n2726) );
  AO221X1 U4697 ( .IN1(WX4423), .IN2(n4455), .IN3(n4288), .IN4(n2761), .IN5(
        n2762), .Q(WX4585) );
  AO22X1 U4698 ( .IN1(n4148), .IN2(CRC_OUT_6_0), .IN3(n4043), .IN4(n2633), .Q(
        n2762) );
  AO221X1 U4699 ( .IN1(WX4421), .IN2(n4455), .IN3(n4288), .IN4(n2764), .IN5(
        n2765), .Q(WX4583) );
  AO22X1 U4700 ( .IN1(n4148), .IN2(CRC_OUT_6_1), .IN3(n4045), .IN4(n2636), .Q(
        n2765) );
  AO221X1 U4701 ( .IN1(WX4419), .IN2(n4455), .IN3(n4288), .IN4(n2767), .IN5(
        n2768), .Q(WX4581) );
  AO22X1 U4702 ( .IN1(n4148), .IN2(CRC_OUT_6_2), .IN3(n4044), .IN4(n2639), .Q(
        n2768) );
  AO221X1 U4703 ( .IN1(WX4417), .IN2(n4455), .IN3(n4289), .IN4(n2770), .IN5(
        n2771), .Q(WX4579) );
  AO22X1 U4704 ( .IN1(n4149), .IN2(CRC_OUT_6_3), .IN3(n4049), .IN4(n2642), .Q(
        n2771) );
  AO221X1 U4705 ( .IN1(WX4415), .IN2(n4455), .IN3(n4289), .IN4(n2773), .IN5(
        n2774), .Q(WX4577) );
  AO22X1 U4706 ( .IN1(n4149), .IN2(CRC_OUT_6_4), .IN3(n4044), .IN4(n2645), .Q(
        n2774) );
  AO221X1 U4707 ( .IN1(WX4413), .IN2(n4456), .IN3(n4289), .IN4(n2776), .IN5(
        n2777), .Q(WX4575) );
  AO22X1 U4708 ( .IN1(n4149), .IN2(CRC_OUT_6_5), .IN3(n4044), .IN4(n2648), .Q(
        n2777) );
  AO221X1 U4709 ( .IN1(WX4411), .IN2(n4456), .IN3(n4289), .IN4(n2779), .IN5(
        n2780), .Q(WX4573) );
  AO22X1 U4710 ( .IN1(n4149), .IN2(CRC_OUT_6_6), .IN3(n4045), .IN4(n2651), .Q(
        n2780) );
  AO221X1 U4711 ( .IN1(WX4409), .IN2(n4456), .IN3(n4290), .IN4(n2782), .IN5(
        n2783), .Q(WX4571) );
  AO22X1 U4712 ( .IN1(n4150), .IN2(CRC_OUT_6_7), .IN3(n4045), .IN4(n2654), .Q(
        n2783) );
  AO221X1 U4713 ( .IN1(WX4407), .IN2(n4456), .IN3(n4290), .IN4(n2785), .IN5(
        n2786), .Q(WX4569) );
  AO22X1 U4714 ( .IN1(n4150), .IN2(CRC_OUT_6_8), .IN3(n4045), .IN4(n2657), .Q(
        n2786) );
  AO221X1 U4715 ( .IN1(WX4405), .IN2(n4456), .IN3(n4290), .IN4(n2788), .IN5(
        n2789), .Q(WX4567) );
  AO22X1 U4716 ( .IN1(n4150), .IN2(CRC_OUT_6_9), .IN3(n4046), .IN4(n2660), .Q(
        n2789) );
  AO221X1 U4717 ( .IN1(WX4403), .IN2(n4457), .IN3(n4290), .IN4(n2791), .IN5(
        n2792), .Q(WX4565) );
  AO22X1 U4718 ( .IN1(n4150), .IN2(CRC_OUT_6_10), .IN3(n4050), .IN4(n2663), 
        .Q(n2792) );
  AO221X1 U4719 ( .IN1(WX4401), .IN2(n4457), .IN3(n4291), .IN4(n2794), .IN5(
        n2795), .Q(WX4563) );
  AO22X1 U4720 ( .IN1(n4151), .IN2(CRC_OUT_6_11), .IN3(n4046), .IN4(n2666), 
        .Q(n2795) );
  AO221X1 U4721 ( .IN1(WX4399), .IN2(n4457), .IN3(n4291), .IN4(n2797), .IN5(
        n2798), .Q(WX4561) );
  AO22X1 U4722 ( .IN1(n4151), .IN2(CRC_OUT_6_12), .IN3(n4046), .IN4(n2669), 
        .Q(n2798) );
  AO221X1 U4723 ( .IN1(WX4397), .IN2(n4457), .IN3(n4291), .IN4(n2800), .IN5(
        n2801), .Q(WX4559) );
  AO22X1 U4724 ( .IN1(n4151), .IN2(CRC_OUT_6_13), .IN3(n4046), .IN4(n2672), 
        .Q(n2801) );
  AO221X1 U4725 ( .IN1(WX4395), .IN2(n4457), .IN3(n4291), .IN4(n2803), .IN5(
        n2804), .Q(WX4557) );
  AO22X1 U4726 ( .IN1(n4151), .IN2(CRC_OUT_6_14), .IN3(n4046), .IN4(n2675), 
        .Q(n2804) );
  AO221X1 U4727 ( .IN1(WX4393), .IN2(n4458), .IN3(n4292), .IN4(n2806), .IN5(
        n2807), .Q(WX4555) );
  AO22X1 U4728 ( .IN1(n4152), .IN2(CRC_OUT_6_15), .IN3(n4047), .IN4(n2678), 
        .Q(n2807) );
  AO221X1 U4729 ( .IN1(WX4391), .IN2(n4458), .IN3(n4292), .IN4(n2809), .IN5(
        n2810), .Q(WX4553) );
  AO22X1 U4730 ( .IN1(n4152), .IN2(CRC_OUT_6_16), .IN3(n4047), .IN4(n2681), 
        .Q(n2810) );
  AO221X1 U4731 ( .IN1(WX4389), .IN2(n4458), .IN3(n4292), .IN4(n2812), .IN5(
        n2813), .Q(WX4551) );
  AO22X1 U4732 ( .IN1(n4152), .IN2(CRC_OUT_6_17), .IN3(n4047), .IN4(n2684), 
        .Q(n2813) );
  AO221X1 U4733 ( .IN1(WX4387), .IN2(n4458), .IN3(n4292), .IN4(n2815), .IN5(
        n2816), .Q(WX4549) );
  AO22X1 U4734 ( .IN1(n4152), .IN2(CRC_OUT_6_18), .IN3(n4047), .IN4(n2687), 
        .Q(n2816) );
  AO221X1 U4735 ( .IN1(WX4385), .IN2(n4458), .IN3(n4293), .IN4(n2818), .IN5(
        n2819), .Q(WX4547) );
  AO22X1 U4736 ( .IN1(n4153), .IN2(CRC_OUT_6_19), .IN3(n4048), .IN4(n2690), 
        .Q(n2819) );
  AO221X1 U4737 ( .IN1(WX4383), .IN2(n4459), .IN3(n4293), .IN4(n2821), .IN5(
        n2822), .Q(WX4545) );
  AO22X1 U4738 ( .IN1(n4153), .IN2(CRC_OUT_6_20), .IN3(n4048), .IN4(n2693), 
        .Q(n2822) );
  AO221X1 U4739 ( .IN1(WX4381), .IN2(n4459), .IN3(n4293), .IN4(n2824), .IN5(
        n2825), .Q(WX4543) );
  AO22X1 U4740 ( .IN1(n4153), .IN2(CRC_OUT_6_21), .IN3(n4048), .IN4(n2696), 
        .Q(n2825) );
  AO221X1 U4741 ( .IN1(WX4379), .IN2(n4459), .IN3(n4293), .IN4(n2827), .IN5(
        n2828), .Q(WX4541) );
  AO22X1 U4742 ( .IN1(n4153), .IN2(CRC_OUT_6_22), .IN3(n4048), .IN4(n2699), 
        .Q(n2828) );
  AO221X1 U4743 ( .IN1(WX4377), .IN2(n4459), .IN3(n4294), .IN4(n2830), .IN5(
        n2831), .Q(WX4539) );
  AO22X1 U4744 ( .IN1(n4154), .IN2(CRC_OUT_6_23), .IN3(n4048), .IN4(n2702), 
        .Q(n2831) );
  AO221X1 U4745 ( .IN1(WX4375), .IN2(n4459), .IN3(n4294), .IN4(n2833), .IN5(
        n2834), .Q(WX4537) );
  AO22X1 U4746 ( .IN1(n4154), .IN2(CRC_OUT_6_24), .IN3(n4049), .IN4(n2705), 
        .Q(n2834) );
  AO221X1 U4747 ( .IN1(WX4373), .IN2(n4460), .IN3(n4294), .IN4(n2836), .IN5(
        n2837), .Q(WX4535) );
  AO22X1 U4748 ( .IN1(n4154), .IN2(CRC_OUT_6_25), .IN3(n4049), .IN4(n2708), 
        .Q(n2837) );
  AO221X1 U4749 ( .IN1(WX4371), .IN2(n4460), .IN3(n4294), .IN4(n2839), .IN5(
        n2840), .Q(WX4533) );
  AO22X1 U4750 ( .IN1(n4154), .IN2(CRC_OUT_6_26), .IN3(n4049), .IN4(n2711), 
        .Q(n2840) );
  AO221X1 U4751 ( .IN1(WX4369), .IN2(n4460), .IN3(n4295), .IN4(n2842), .IN5(
        n2843), .Q(WX4531) );
  AO22X1 U4752 ( .IN1(n4155), .IN2(CRC_OUT_6_27), .IN3(n4049), .IN4(n2714), 
        .Q(n2843) );
  AO221X1 U4753 ( .IN1(WX4367), .IN2(n4460), .IN3(n4295), .IN4(n2845), .IN5(
        n2846), .Q(WX4529) );
  AO22X1 U4754 ( .IN1(n4155), .IN2(CRC_OUT_6_28), .IN3(n4050), .IN4(n2717), 
        .Q(n2846) );
  AO221X1 U4755 ( .IN1(WX4365), .IN2(n4460), .IN3(n4295), .IN4(n2848), .IN5(
        n2849), .Q(WX4527) );
  AO22X1 U4756 ( .IN1(n4155), .IN2(CRC_OUT_6_29), .IN3(n4050), .IN4(n2720), 
        .Q(n2849) );
  AO221X1 U4757 ( .IN1(WX4363), .IN2(n4461), .IN3(n4295), .IN4(n2851), .IN5(
        n2852), .Q(WX4525) );
  AO22X1 U4758 ( .IN1(n4155), .IN2(CRC_OUT_6_30), .IN3(n4050), .IN4(n2723), 
        .Q(n2852) );
  AO221X1 U4759 ( .IN1(WX4364), .IN2(n2245), .IN3(n4034), .IN4(n2727), .IN5(
        n2854), .Q(WX4523) );
  AO22X1 U4760 ( .IN1(n4354), .IN2(n2855), .IN3(n4214), .IN4(CRC_OUT_6_31), 
        .Q(n2854) );
  AO221X1 U4761 ( .IN1(WX3130), .IN2(n4461), .IN3(n4296), .IN4(n2889), .IN5(
        n2890), .Q(WX3292) );
  AO22X1 U4762 ( .IN1(n4156), .IN2(CRC_OUT_7_0), .IN3(n4050), .IN4(n2761), .Q(
        n2890) );
  AO221X1 U4763 ( .IN1(WX3128), .IN2(n4461), .IN3(n4296), .IN4(n2892), .IN5(
        n2893), .Q(WX3290) );
  AO22X1 U4764 ( .IN1(n4156), .IN2(CRC_OUT_7_1), .IN3(n4051), .IN4(n2764), .Q(
        n2893) );
  AO221X1 U4765 ( .IN1(WX3126), .IN2(n4461), .IN3(n4296), .IN4(n2895), .IN5(
        n2896), .Q(WX3288) );
  AO22X1 U4766 ( .IN1(n4156), .IN2(CRC_OUT_7_2), .IN3(n4051), .IN4(n2767), .Q(
        n2896) );
  AO221X1 U4767 ( .IN1(WX3124), .IN2(n4461), .IN3(n4296), .IN4(n2898), .IN5(
        n2899), .Q(WX3286) );
  AO22X1 U4768 ( .IN1(n4156), .IN2(CRC_OUT_7_3), .IN3(n4051), .IN4(n2770), .Q(
        n2899) );
  AO221X1 U4769 ( .IN1(WX3122), .IN2(n4462), .IN3(n4297), .IN4(n2901), .IN5(
        n2902), .Q(WX3284) );
  AO22X1 U4770 ( .IN1(n4157), .IN2(CRC_OUT_7_4), .IN3(n4051), .IN4(n2773), .Q(
        n2902) );
  AO221X1 U4771 ( .IN1(WX3120), .IN2(n4462), .IN3(n4297), .IN4(n2904), .IN5(
        n2905), .Q(WX3282) );
  AO22X1 U4772 ( .IN1(n4157), .IN2(CRC_OUT_7_5), .IN3(n4051), .IN4(n2776), .Q(
        n2905) );
  AO221X1 U4773 ( .IN1(WX3118), .IN2(n4462), .IN3(n4297), .IN4(n2907), .IN5(
        n2908), .Q(WX3280) );
  AO22X1 U4774 ( .IN1(n4157), .IN2(CRC_OUT_7_6), .IN3(n4052), .IN4(n2779), .Q(
        n2908) );
  AO221X1 U4775 ( .IN1(WX3116), .IN2(n4462), .IN3(n4297), .IN4(n2910), .IN5(
        n2911), .Q(WX3278) );
  AO22X1 U4776 ( .IN1(n4157), .IN2(CRC_OUT_7_7), .IN3(n4052), .IN4(n2782), .Q(
        n2911) );
  AO221X1 U4777 ( .IN1(WX3114), .IN2(n4462), .IN3(n4298), .IN4(n2913), .IN5(
        n2914), .Q(WX3276) );
  AO22X1 U4778 ( .IN1(n4158), .IN2(CRC_OUT_7_8), .IN3(n4052), .IN4(n2785), .Q(
        n2914) );
  AO221X1 U4779 ( .IN1(WX3112), .IN2(n4463), .IN3(n4298), .IN4(n2916), .IN5(
        n2917), .Q(WX3274) );
  AO22X1 U4780 ( .IN1(n4158), .IN2(CRC_OUT_7_9), .IN3(n4052), .IN4(n2788), .Q(
        n2917) );
  AO221X1 U4781 ( .IN1(WX3110), .IN2(n4463), .IN3(n4298), .IN4(n2919), .IN5(
        n2920), .Q(WX3272) );
  AO22X1 U4782 ( .IN1(n4158), .IN2(CRC_OUT_7_10), .IN3(n4053), .IN4(n2791), 
        .Q(n2920) );
  AO221X1 U4783 ( .IN1(WX3108), .IN2(n4463), .IN3(n4298), .IN4(n2922), .IN5(
        n2923), .Q(WX3270) );
  AO22X1 U4784 ( .IN1(n4158), .IN2(CRC_OUT_7_11), .IN3(n4053), .IN4(n2794), 
        .Q(n2923) );
  AO221X1 U4785 ( .IN1(WX3106), .IN2(n4463), .IN3(n4299), .IN4(n2925), .IN5(
        n2926), .Q(WX3268) );
  AO22X1 U4786 ( .IN1(n4159), .IN2(CRC_OUT_7_12), .IN3(n4053), .IN4(n2797), 
        .Q(n2926) );
  AO221X1 U4787 ( .IN1(WX3104), .IN2(n4463), .IN3(n4299), .IN4(n2928), .IN5(
        n2929), .Q(WX3266) );
  AO22X1 U4788 ( .IN1(n4159), .IN2(CRC_OUT_7_13), .IN3(n4053), .IN4(n2800), 
        .Q(n2929) );
  AO221X1 U4789 ( .IN1(WX3102), .IN2(n4464), .IN3(n4299), .IN4(n2931), .IN5(
        n2932), .Q(WX3264) );
  AO22X1 U4790 ( .IN1(n4159), .IN2(CRC_OUT_7_14), .IN3(n4053), .IN4(n2803), 
        .Q(n2932) );
  AO221X1 U4791 ( .IN1(WX3100), .IN2(n4464), .IN3(n4299), .IN4(n2934), .IN5(
        n2935), .Q(WX3262) );
  AO22X1 U4792 ( .IN1(n4159), .IN2(CRC_OUT_7_15), .IN3(n4054), .IN4(n2806), 
        .Q(n2935) );
  AO221X1 U4793 ( .IN1(WX3098), .IN2(n4464), .IN3(n4300), .IN4(n2937), .IN5(
        n2938), .Q(WX3260) );
  AO22X1 U4794 ( .IN1(n4160), .IN2(CRC_OUT_7_16), .IN3(n4054), .IN4(n2809), 
        .Q(n2938) );
  AO221X1 U4795 ( .IN1(WX3096), .IN2(n4464), .IN3(n4300), .IN4(n2940), .IN5(
        n2941), .Q(WX3258) );
  AO22X1 U4796 ( .IN1(n4160), .IN2(CRC_OUT_7_17), .IN3(n4054), .IN4(n2812), 
        .Q(n2941) );
  AO221X1 U4797 ( .IN1(WX3094), .IN2(n4464), .IN3(n4300), .IN4(n2943), .IN5(
        n2944), .Q(WX3256) );
  AO22X1 U4798 ( .IN1(n4160), .IN2(CRC_OUT_7_18), .IN3(n4054), .IN4(n2815), 
        .Q(n2944) );
  AO221X1 U4799 ( .IN1(WX3092), .IN2(n4465), .IN3(n4300), .IN4(n2946), .IN5(
        n2947), .Q(WX3254) );
  AO22X1 U4800 ( .IN1(n4160), .IN2(CRC_OUT_7_19), .IN3(n4054), .IN4(n2818), 
        .Q(n2947) );
  AO221X1 U4801 ( .IN1(WX3090), .IN2(n4465), .IN3(n4301), .IN4(n2949), .IN5(
        n2950), .Q(WX3252) );
  AO22X1 U4802 ( .IN1(n4161), .IN2(CRC_OUT_7_20), .IN3(n4055), .IN4(n2821), 
        .Q(n2950) );
  AO221X1 U4803 ( .IN1(WX3088), .IN2(n4465), .IN3(n4301), .IN4(n2952), .IN5(
        n2953), .Q(WX3250) );
  AO22X1 U4804 ( .IN1(n4161), .IN2(CRC_OUT_7_21), .IN3(n4055), .IN4(n2824), 
        .Q(n2953) );
  AO221X1 U4805 ( .IN1(WX3086), .IN2(n4465), .IN3(n4301), .IN4(n2955), .IN5(
        n2956), .Q(WX3248) );
  AO22X1 U4806 ( .IN1(n4161), .IN2(CRC_OUT_7_22), .IN3(n4055), .IN4(n2827), 
        .Q(n2956) );
  AO221X1 U4807 ( .IN1(WX3084), .IN2(n4465), .IN3(n4319), .IN4(n2958), .IN5(
        n2959), .Q(WX3246) );
  AO22X1 U4808 ( .IN1(n4179), .IN2(CRC_OUT_7_23), .IN3(n4063), .IN4(n2830), 
        .Q(n2959) );
  AO221X1 U4809 ( .IN1(WX3082), .IN2(n4466), .IN3(n4302), .IN4(n2961), .IN5(
        n2962), .Q(WX3244) );
  AO22X1 U4810 ( .IN1(n4162), .IN2(CRC_OUT_7_24), .IN3(n4055), .IN4(n2833), 
        .Q(n2962) );
  AO221X1 U4811 ( .IN1(WX3080), .IN2(n4466), .IN3(n4302), .IN4(n2964), .IN5(
        n2965), .Q(WX3242) );
  AO22X1 U4812 ( .IN1(n4162), .IN2(CRC_OUT_7_25), .IN3(n4055), .IN4(n2836), 
        .Q(n2965) );
  AO221X1 U4813 ( .IN1(WX3078), .IN2(n4466), .IN3(n4302), .IN4(n2967), .IN5(
        n2968), .Q(WX3240) );
  AO22X1 U4814 ( .IN1(n4162), .IN2(CRC_OUT_7_26), .IN3(n4056), .IN4(n2839), 
        .Q(n2968) );
  AO221X1 U4815 ( .IN1(WX3076), .IN2(n4466), .IN3(n4302), .IN4(n2970), .IN5(
        n2971), .Q(WX3238) );
  AO22X1 U4816 ( .IN1(n4162), .IN2(CRC_OUT_7_27), .IN3(n4056), .IN4(n2842), 
        .Q(n2971) );
  AO221X1 U4817 ( .IN1(WX3074), .IN2(n4466), .IN3(n4303), .IN4(n2973), .IN5(
        n2974), .Q(WX3236) );
  AO22X1 U4818 ( .IN1(n4163), .IN2(CRC_OUT_7_28), .IN3(n4056), .IN4(n2845), 
        .Q(n2974) );
  AO221X1 U4819 ( .IN1(WX3072), .IN2(n4467), .IN3(n4303), .IN4(n2976), .IN5(
        n2977), .Q(WX3234) );
  AO22X1 U4820 ( .IN1(n4163), .IN2(CRC_OUT_7_29), .IN3(n4056), .IN4(n2848), 
        .Q(n2977) );
  AO221X1 U4821 ( .IN1(WX3070), .IN2(n4467), .IN3(n4303), .IN4(n2979), .IN5(
        n2980), .Q(WX3232) );
  AO22X1 U4822 ( .IN1(n4163), .IN2(CRC_OUT_7_30), .IN3(n4056), .IN4(n2851), 
        .Q(n2980) );
  AO221X1 U4823 ( .IN1(WX3071), .IN2(n2245), .IN3(n4035), .IN4(n2855), .IN5(
        n2982), .Q(WX3230) );
  AO22X1 U4824 ( .IN1(n4354), .IN2(n2983), .IN3(n4214), .IN4(CRC_OUT_7_31), 
        .Q(n2982) );
  AO221X1 U4825 ( .IN1(WX1837), .IN2(n4467), .IN3(n4303), .IN4(n2507), .IN5(
        n3017), .Q(WX1999) );
  AO22X1 U4826 ( .IN1(n4163), .IN2(CRC_OUT_8_0), .IN3(n4057), .IN4(n2889), .Q(
        n3017) );
  AO221X1 U4827 ( .IN1(WX1835), .IN2(n4467), .IN3(n4304), .IN4(n2510), .IN5(
        n3020), .Q(WX1997) );
  AO22X1 U4828 ( .IN1(n4164), .IN2(CRC_OUT_8_1), .IN3(n4057), .IN4(n2892), .Q(
        n3020) );
  AO221X1 U4829 ( .IN1(WX1833), .IN2(n4467), .IN3(n4304), .IN4(n2513), .IN5(
        n3023), .Q(WX1995) );
  AO22X1 U4830 ( .IN1(n4164), .IN2(CRC_OUT_8_2), .IN3(n4057), .IN4(n2895), .Q(
        n3023) );
  AO221X1 U4831 ( .IN1(WX1831), .IN2(n4468), .IN3(n4304), .IN4(n2516), .IN5(
        n3026), .Q(WX1993) );
  AO22X1 U4832 ( .IN1(n4164), .IN2(CRC_OUT_8_3), .IN3(n4057), .IN4(n2898), .Q(
        n3026) );
  AO221X1 U4833 ( .IN1(WX1829), .IN2(n4468), .IN3(n4304), .IN4(n2519), .IN5(
        n3029), .Q(WX1991) );
  AO22X1 U4834 ( .IN1(n4164), .IN2(CRC_OUT_8_4), .IN3(n4057), .IN4(n2901), .Q(
        n3029) );
  AO221X1 U4835 ( .IN1(WX1827), .IN2(n4468), .IN3(n4305), .IN4(n2522), .IN5(
        n3032), .Q(WX1989) );
  AO22X1 U4836 ( .IN1(n4165), .IN2(CRC_OUT_8_5), .IN3(n4058), .IN4(n2904), .Q(
        n3032) );
  AO221X1 U4837 ( .IN1(WX1825), .IN2(n4468), .IN3(n4305), .IN4(n2525), .IN5(
        n3035), .Q(WX1987) );
  AO22X1 U4838 ( .IN1(n4165), .IN2(CRC_OUT_8_6), .IN3(n4058), .IN4(n2907), .Q(
        n3035) );
  AO221X1 U4839 ( .IN1(WX1823), .IN2(n4468), .IN3(n4305), .IN4(n2528), .IN5(
        n3038), .Q(WX1985) );
  AO22X1 U4840 ( .IN1(n4165), .IN2(CRC_OUT_8_7), .IN3(n4058), .IN4(n2910), .Q(
        n3038) );
  AO221X1 U4841 ( .IN1(WX1821), .IN2(n4469), .IN3(n4305), .IN4(n2531), .IN5(
        n3041), .Q(WX1983) );
  AO22X1 U4842 ( .IN1(n4165), .IN2(CRC_OUT_8_8), .IN3(n4058), .IN4(n2913), .Q(
        n3041) );
  AO221X1 U4843 ( .IN1(WX1819), .IN2(n4469), .IN3(n4306), .IN4(n2534), .IN5(
        n3044), .Q(WX1981) );
  AO22X1 U4844 ( .IN1(n4166), .IN2(CRC_OUT_8_9), .IN3(n4058), .IN4(n2916), .Q(
        n3044) );
  AO221X1 U4845 ( .IN1(WX1817), .IN2(n4469), .IN3(n4306), .IN4(n2537), .IN5(
        n3047), .Q(WX1979) );
  AO22X1 U4846 ( .IN1(n4166), .IN2(CRC_OUT_8_10), .IN3(n4059), .IN4(n2919), 
        .Q(n3047) );
  AO221X1 U4847 ( .IN1(WX1815), .IN2(n4469), .IN3(n4306), .IN4(n2540), .IN5(
        n3050), .Q(WX1977) );
  AO22X1 U4848 ( .IN1(n4166), .IN2(CRC_OUT_8_11), .IN3(n4059), .IN4(n2922), 
        .Q(n3050) );
  AO221X1 U4849 ( .IN1(WX1813), .IN2(n4469), .IN3(n4306), .IN4(n2543), .IN5(
        n3053), .Q(WX1975) );
  AO22X1 U4850 ( .IN1(n4166), .IN2(CRC_OUT_8_12), .IN3(n4059), .IN4(n2925), 
        .Q(n3053) );
  AO221X1 U4851 ( .IN1(WX1811), .IN2(n4470), .IN3(n4307), .IN4(n2546), .IN5(
        n3056), .Q(WX1973) );
  AO22X1 U4852 ( .IN1(n4167), .IN2(CRC_OUT_8_13), .IN3(n4059), .IN4(n2928), 
        .Q(n3056) );
  AO221X1 U4853 ( .IN1(WX1809), .IN2(n4470), .IN3(n4307), .IN4(n2549), .IN5(
        n3059), .Q(WX1971) );
  AO22X1 U4854 ( .IN1(n4167), .IN2(CRC_OUT_8_14), .IN3(n4059), .IN4(n2931), 
        .Q(n3059) );
  AO221X1 U4855 ( .IN1(WX1807), .IN2(n4470), .IN3(n4307), .IN4(n2552), .IN5(
        n3062), .Q(WX1969) );
  AO22X1 U4856 ( .IN1(n4167), .IN2(CRC_OUT_8_15), .IN3(n4060), .IN4(n2934), 
        .Q(n3062) );
  AO221X1 U4857 ( .IN1(WX1805), .IN2(n4470), .IN3(n4307), .IN4(n2555), .IN5(
        n3065), .Q(WX1967) );
  AO22X1 U4858 ( .IN1(n4167), .IN2(CRC_OUT_8_16), .IN3(n4060), .IN4(n2937), 
        .Q(n3065) );
  AO221X1 U4859 ( .IN1(WX1803), .IN2(n4470), .IN3(n4308), .IN4(n2558), .IN5(
        n3068), .Q(WX1965) );
  AO22X1 U4860 ( .IN1(n4168), .IN2(CRC_OUT_8_17), .IN3(n4060), .IN4(n2940), 
        .Q(n3068) );
  AO221X1 U4861 ( .IN1(WX1801), .IN2(n4471), .IN3(n4308), .IN4(n2561), .IN5(
        n3071), .Q(WX1963) );
  AO22X1 U4862 ( .IN1(n4168), .IN2(CRC_OUT_8_18), .IN3(n4060), .IN4(n2943), 
        .Q(n3071) );
  AO221X1 U4863 ( .IN1(WX1799), .IN2(n4471), .IN3(n4308), .IN4(n2564), .IN5(
        n3074), .Q(WX1961) );
  AO22X1 U4864 ( .IN1(n4168), .IN2(CRC_OUT_8_19), .IN3(n4060), .IN4(n2946), 
        .Q(n3074) );
  AO221X1 U4865 ( .IN1(WX1797), .IN2(n4471), .IN3(n4308), .IN4(n2567), .IN5(
        n3077), .Q(WX1959) );
  AO22X1 U4866 ( .IN1(n4168), .IN2(CRC_OUT_8_20), .IN3(n4061), .IN4(n2949), 
        .Q(n3077) );
  AO221X1 U4867 ( .IN1(WX1795), .IN2(n4471), .IN3(n4309), .IN4(n2570), .IN5(
        n3080), .Q(WX1957) );
  AO22X1 U4868 ( .IN1(n4169), .IN2(CRC_OUT_8_21), .IN3(n4061), .IN4(n2952), 
        .Q(n3080) );
  AO221X1 U4869 ( .IN1(WX1793), .IN2(n4471), .IN3(n4309), .IN4(n2573), .IN5(
        n3083), .Q(WX1955) );
  AO22X1 U4870 ( .IN1(n4169), .IN2(CRC_OUT_8_22), .IN3(n4061), .IN4(n2955), 
        .Q(n3083) );
  AO221X1 U4871 ( .IN1(WX1791), .IN2(n4472), .IN3(n4309), .IN4(n2576), .IN5(
        n3086), .Q(WX1953) );
  AO22X1 U4872 ( .IN1(n4169), .IN2(CRC_OUT_8_23), .IN3(n4061), .IN4(n2958), 
        .Q(n3086) );
  AO221X1 U4873 ( .IN1(WX1789), .IN2(n4472), .IN3(n4309), .IN4(n2579), .IN5(
        n3089), .Q(WX1951) );
  AO22X1 U4874 ( .IN1(n4169), .IN2(CRC_OUT_8_24), .IN3(n4061), .IN4(n2961), 
        .Q(n3089) );
  AO221X1 U4875 ( .IN1(WX1787), .IN2(n4472), .IN3(n4310), .IN4(n2582), .IN5(
        n3092), .Q(WX1949) );
  AO22X1 U4876 ( .IN1(n4170), .IN2(CRC_OUT_8_25), .IN3(n4062), .IN4(n2964), 
        .Q(n3092) );
  AO221X1 U4877 ( .IN1(WX1785), .IN2(n4472), .IN3(n4310), .IN4(n2585), .IN5(
        n3095), .Q(WX1947) );
  AO22X1 U4878 ( .IN1(n4170), .IN2(CRC_OUT_8_26), .IN3(n4062), .IN4(n2967), 
        .Q(n3095) );
  AO221X1 U4879 ( .IN1(WX1783), .IN2(n4472), .IN3(n4310), .IN4(n2588), .IN5(
        n3098), .Q(WX1945) );
  AO22X1 U4880 ( .IN1(n4170), .IN2(CRC_OUT_8_27), .IN3(n4062), .IN4(n2970), 
        .Q(n3098) );
  AO221X1 U4881 ( .IN1(WX1781), .IN2(n4473), .IN3(n4310), .IN4(n2591), .IN5(
        n3101), .Q(WX1943) );
  AO22X1 U4882 ( .IN1(n4170), .IN2(CRC_OUT_8_28), .IN3(n4062), .IN4(n2973), 
        .Q(n3101) );
  AO221X1 U4883 ( .IN1(WX1779), .IN2(n4473), .IN3(n4311), .IN4(n2604), .IN5(
        n3104), .Q(WX1941) );
  AO22X1 U4884 ( .IN1(n4171), .IN2(CRC_OUT_8_29), .IN3(n4062), .IN4(n2976), 
        .Q(n3104) );
  AO221X1 U4885 ( .IN1(WX1777), .IN2(n4473), .IN3(n4311), .IN4(n2617), .IN5(
        n3107), .Q(WX1939) );
  AO22X1 U4886 ( .IN1(n4171), .IN2(CRC_OUT_8_30), .IN3(n4063), .IN4(n2979), 
        .Q(n3107) );
  AO221X1 U4887 ( .IN1(WX1778), .IN2(n2245), .IN3(n4034), .IN4(n2983), .IN5(
        n3110), .Q(WX1937) );
  AO22X1 U4888 ( .IN1(n4355), .IN2(n2628), .IN3(n4215), .IN4(CRC_OUT_8_31), 
        .Q(n3110) );
  AO221X1 U4889 ( .IN1(WX544), .IN2(n4442), .IN3(n4341), .IN4(n2505), .IN5(
        n2506), .Q(WX706) );
  AO22X1 U4890 ( .IN1(n4201), .IN2(CRC_OUT_9_0), .IN3(n4081), .IN4(n2507), .Q(
        n2506) );
  AO221X1 U4891 ( .IN1(WX542), .IN2(n4442), .IN3(n4343), .IN4(n2508), .IN5(
        n2509), .Q(WX704) );
  AO22X1 U4892 ( .IN1(n4203), .IN2(CRC_OUT_9_1), .IN3(n4082), .IN4(n2510), .Q(
        n2509) );
  AO221X1 U4893 ( .IN1(WX540), .IN2(n4443), .IN3(n4343), .IN4(n2511), .IN5(
        n2512), .Q(WX702) );
  AO22X1 U4894 ( .IN1(n4203), .IN2(CRC_OUT_9_2), .IN3(n4082), .IN4(n2513), .Q(
        n2512) );
  AO221X1 U4895 ( .IN1(WX538), .IN2(n4443), .IN3(n4343), .IN4(n2514), .IN5(
        n2515), .Q(WX700) );
  AO22X1 U4896 ( .IN1(n4203), .IN2(CRC_OUT_9_3), .IN3(n4082), .IN4(n2516), .Q(
        n2515) );
  AO221X1 U4897 ( .IN1(WX536), .IN2(n4443), .IN3(n4343), .IN4(n2517), .IN5(
        n2518), .Q(WX698) );
  AO22X1 U4898 ( .IN1(n4203), .IN2(CRC_OUT_9_4), .IN3(n4082), .IN4(n2519), .Q(
        n2518) );
  AO221X1 U4899 ( .IN1(WX534), .IN2(n4443), .IN3(n4344), .IN4(n2520), .IN5(
        n2521), .Q(WX696) );
  AO22X1 U4900 ( .IN1(n4204), .IN2(CRC_OUT_9_5), .IN3(n4082), .IN4(n2522), .Q(
        n2521) );
  AO221X1 U4901 ( .IN1(WX532), .IN2(n4443), .IN3(n4342), .IN4(n2523), .IN5(
        n2524), .Q(WX694) );
  AO22X1 U4902 ( .IN1(n4202), .IN2(CRC_OUT_9_6), .IN3(n4083), .IN4(n2525), .Q(
        n2524) );
  AO221X1 U4903 ( .IN1(WX530), .IN2(n4444), .IN3(n4344), .IN4(n2526), .IN5(
        n2527), .Q(WX692) );
  AO22X1 U4904 ( .IN1(n4204), .IN2(CRC_OUT_9_7), .IN3(n4083), .IN4(n2528), .Q(
        n2527) );
  AO221X1 U4905 ( .IN1(WX528), .IN2(n4444), .IN3(n4344), .IN4(n2529), .IN5(
        n2530), .Q(WX690) );
  AO22X1 U4906 ( .IN1(n4204), .IN2(CRC_OUT_9_8), .IN3(n4083), .IN4(n2531), .Q(
        n2530) );
  AO221X1 U4907 ( .IN1(WX526), .IN2(n4444), .IN3(n4345), .IN4(n2532), .IN5(
        n2533), .Q(WX688) );
  AO22X1 U4908 ( .IN1(n4205), .IN2(CRC_OUT_9_9), .IN3(n4083), .IN4(n2534), .Q(
        n2533) );
  AO221X1 U4909 ( .IN1(WX524), .IN2(n4444), .IN3(n4345), .IN4(n2535), .IN5(
        n2536), .Q(WX686) );
  AO22X1 U4910 ( .IN1(n4205), .IN2(CRC_OUT_9_10), .IN3(n4083), .IN4(n2537), 
        .Q(n2536) );
  AO221X1 U4911 ( .IN1(WX522), .IN2(n4444), .IN3(n4345), .IN4(n2538), .IN5(
        n2539), .Q(WX684) );
  AO22X1 U4912 ( .IN1(n4205), .IN2(CRC_OUT_9_11), .IN3(n4084), .IN4(n2540), 
        .Q(n2539) );
  AO221X1 U4913 ( .IN1(WX520), .IN2(n4445), .IN3(n4344), .IN4(n2541), .IN5(
        n2542), .Q(WX682) );
  AO22X1 U4914 ( .IN1(n4204), .IN2(CRC_OUT_9_12), .IN3(n4084), .IN4(n2543), 
        .Q(n2542) );
  AO221X1 U4915 ( .IN1(WX518), .IN2(n4445), .IN3(n4346), .IN4(n2544), .IN5(
        n2545), .Q(WX680) );
  AO22X1 U4916 ( .IN1(n4206), .IN2(CRC_OUT_9_13), .IN3(n4084), .IN4(n2546), 
        .Q(n2545) );
  AO221X1 U4917 ( .IN1(WX516), .IN2(n4445), .IN3(n4346), .IN4(n2547), .IN5(
        n2548), .Q(WX678) );
  AO22X1 U4918 ( .IN1(n4206), .IN2(CRC_OUT_9_14), .IN3(n4084), .IN4(n2549), 
        .Q(n2548) );
  AO221X1 U4919 ( .IN1(WX514), .IN2(n4445), .IN3(n4346), .IN4(n2550), .IN5(
        n2551), .Q(WX676) );
  AO22X1 U4920 ( .IN1(n4206), .IN2(CRC_OUT_9_15), .IN3(n4084), .IN4(n2552), 
        .Q(n2551) );
  AO221X1 U4921 ( .IN1(WX512), .IN2(n4445), .IN3(n4347), .IN4(n2553), .IN5(
        n2554), .Q(WX674) );
  AO22X1 U4922 ( .IN1(n4207), .IN2(CRC_OUT_9_16), .IN3(n4085), .IN4(n2555), 
        .Q(n2554) );
  AO221X1 U4923 ( .IN1(WX510), .IN2(n4446), .IN3(n4347), .IN4(n2556), .IN5(
        n2557), .Q(WX672) );
  AO22X1 U4924 ( .IN1(n4207), .IN2(CRC_OUT_9_17), .IN3(n4085), .IN4(n2558), 
        .Q(n2557) );
  AO221X1 U4925 ( .IN1(WX508), .IN2(n4446), .IN3(n4347), .IN4(n2559), .IN5(
        n2560), .Q(WX670) );
  AO22X1 U4926 ( .IN1(n4207), .IN2(CRC_OUT_9_18), .IN3(n4085), .IN4(n2561), 
        .Q(n2560) );
  AO221X1 U4927 ( .IN1(WX506), .IN2(n4446), .IN3(n4348), .IN4(n2562), .IN5(
        n2563), .Q(WX668) );
  AO22X1 U4928 ( .IN1(n4208), .IN2(CRC_OUT_9_19), .IN3(n4085), .IN4(n2564), 
        .Q(n2563) );
  AO221X1 U4929 ( .IN1(WX504), .IN2(n4446), .IN3(n4347), .IN4(n2565), .IN5(
        n2566), .Q(WX666) );
  AO22X1 U4930 ( .IN1(n4207), .IN2(CRC_OUT_9_20), .IN3(n4085), .IN4(n2567), 
        .Q(n2566) );
  AO221X1 U4931 ( .IN1(WX502), .IN2(n4446), .IN3(n4348), .IN4(n2568), .IN5(
        n2569), .Q(WX664) );
  AO22X1 U4932 ( .IN1(n4208), .IN2(CRC_OUT_9_21), .IN3(n4086), .IN4(n2570), 
        .Q(n2569) );
  AO221X1 U4933 ( .IN1(WX500), .IN2(n4447), .IN3(n4346), .IN4(n2571), .IN5(
        n2572), .Q(WX662) );
  AO22X1 U4934 ( .IN1(n4206), .IN2(CRC_OUT_9_22), .IN3(n4086), .IN4(n2573), 
        .Q(n2572) );
  AO221X1 U4935 ( .IN1(WX498), .IN2(n4447), .IN3(n4349), .IN4(n2574), .IN5(
        n2575), .Q(WX660) );
  AO22X1 U4936 ( .IN1(n4209), .IN2(CRC_OUT_9_23), .IN3(n4086), .IN4(n2576), 
        .Q(n2575) );
  AO221X1 U4937 ( .IN1(WX496), .IN2(n4447), .IN3(n4348), .IN4(n2577), .IN5(
        n2578), .Q(WX658) );
  AO22X1 U4938 ( .IN1(n4208), .IN2(CRC_OUT_9_24), .IN3(n4086), .IN4(n2579), 
        .Q(n2578) );
  AO221X1 U4939 ( .IN1(WX494), .IN2(n4447), .IN3(n4349), .IN4(n2580), .IN5(
        n2581), .Q(WX656) );
  AO22X1 U4940 ( .IN1(n4209), .IN2(CRC_OUT_9_25), .IN3(n4086), .IN4(n2582), 
        .Q(n2581) );
  AO221X1 U4941 ( .IN1(WX492), .IN2(n4447), .IN3(n4349), .IN4(n2583), .IN5(
        n2584), .Q(WX654) );
  AO22X1 U4942 ( .IN1(n4209), .IN2(CRC_OUT_9_26), .IN3(n4087), .IN4(n2585), 
        .Q(n2584) );
  AO221X1 U4943 ( .IN1(WX490), .IN2(n4448), .IN3(n4350), .IN4(n2586), .IN5(
        n2587), .Q(WX652) );
  AO22X1 U4944 ( .IN1(n4210), .IN2(CRC_OUT_9_27), .IN3(n4087), .IN4(n2588), 
        .Q(n2587) );
  AO221X1 U4945 ( .IN1(WX488), .IN2(n4448), .IN3(n4348), .IN4(n2589), .IN5(
        n2590), .Q(WX650) );
  AO22X1 U4946 ( .IN1(n4208), .IN2(CRC_OUT_9_28), .IN3(n4087), .IN4(n2591), 
        .Q(n2590) );
  AO221X1 U4947 ( .IN1(WX486), .IN2(n4448), .IN3(n4350), .IN4(n2602), .IN5(
        n2603), .Q(WX648) );
  AO22X1 U4948 ( .IN1(n4210), .IN2(CRC_OUT_9_29), .IN3(n4087), .IN4(n2604), 
        .Q(n2603) );
  AO221X1 U4949 ( .IN1(WX484), .IN2(n4448), .IN3(n4345), .IN4(n2615), .IN5(
        n2616), .Q(WX646) );
  AO22X1 U4950 ( .IN1(n4205), .IN2(CRC_OUT_9_30), .IN3(n4087), .IN4(n2617), 
        .Q(n2616) );
  AO221X1 U4951 ( .IN1(WX485), .IN2(n2245), .IN3(n4034), .IN4(n2628), .IN5(
        n2629), .Q(WX644) );
  AO22X1 U4952 ( .IN1(n4355), .IN2(n2630), .IN3(n4215), .IN4(CRC_OUT_9_31), 
        .Q(n2629) );
  AO221X1 U4953 ( .IN1(WX10829), .IN2(n2245), .IN3(DATA_0_31), .IN4(n4034), 
        .IN5(n3277), .Q(WX10988) );
  AO22X1 U4954 ( .IN1(n4355), .IN2(n2246), .IN3(n4215), .IN4(CRC_OUT_1_31), 
        .Q(n3277) );
  INVX0 U4955 ( .IN(RESET), .QN(n1729) );
  XNOR3X1 U4956 ( .IN1(n3279), .IN2(n4751), .IN3(n3338), .Q(n2246) );
  XOR3X1 U4957 ( .IN1(WX11181), .IN2(WX11117), .IN3(WX11053), .Q(n3279) );
  XNOR3X1 U4958 ( .IN1(n2376), .IN2(n4744), .IN3(n3339), .Q(n2248) );
  XOR3X1 U4959 ( .IN1(test_so85), .IN2(WX9824), .IN3(WX9760), .Q(n2376) );
  XNOR3X1 U4960 ( .IN1(n2504), .IN2(n4745), .IN3(n3340), .Q(n2375) );
  XOR3X1 U4961 ( .IN1(WX8595), .IN2(WX8531), .IN3(WX8467), .Q(n2504) );
  XNOR3X1 U4962 ( .IN1(n2728), .IN2(n4746), .IN3(n3341), .Q(n2503) );
  XOR3X1 U4963 ( .IN1(WX7302), .IN2(WX7238), .IN3(WX7174), .Q(n2728) );
  XNOR3X1 U4964 ( .IN1(n2856), .IN2(n4747), .IN3(n3342), .Q(n2727) );
  XOR3X1 U4965 ( .IN1(WX6009), .IN2(WX5945), .IN3(WX5881), .Q(n2856) );
  XNOR3X1 U4966 ( .IN1(n2984), .IN2(n4749), .IN3(n3343), .Q(n2855) );
  XOR3X1 U4967 ( .IN1(WX4716), .IN2(WX4652), .IN3(WX4588), .Q(n2984) );
  XNOR3X1 U4968 ( .IN1(n3112), .IN2(n4750), .IN3(n3344), .Q(n2983) );
  XOR3X1 U4969 ( .IN1(WX3423), .IN2(WX3359), .IN3(WX3295), .Q(n3112) );
  XNOR3X1 U4970 ( .IN1(n3111), .IN2(n4750), .IN3(n3345), .Q(n2628) );
  XOR3X1 U4971 ( .IN1(WX2130), .IN2(WX2066), .IN3(WX2002), .Q(n3111) );
  XNOR3X1 U4972 ( .IN1(n3246), .IN2(n4762), .IN3(n3346), .Q(n2202) );
  XOR3X1 U4973 ( .IN1(WX11211), .IN2(WX11147), .IN3(WX11083), .Q(n3246) );
  XNOR3X1 U4974 ( .IN1(n3248), .IN2(n4763), .IN3(n3347), .Q(n2205) );
  XOR3X1 U4975 ( .IN1(WX11209), .IN2(WX11145), .IN3(WX11081), .Q(n3248) );
  XNOR3X1 U4976 ( .IN1(n3250), .IN2(n4762), .IN3(n3348), .Q(n2208) );
  XOR3X1 U4977 ( .IN1(WX11207), .IN2(WX11143), .IN3(WX11079), .Q(n3250) );
  XNOR3X1 U4978 ( .IN1(n3252), .IN2(n4763), .IN3(n3349), .Q(n2211) );
  XOR3X1 U4979 ( .IN1(test_so97), .IN2(WX11141), .IN3(WX11077), .Q(n3252) );
  XNOR3X1 U4980 ( .IN1(n3254), .IN2(n4751), .IN3(n3350), .Q(n2214) );
  XOR3X1 U4981 ( .IN1(WX11203), .IN2(WX11139), .IN3(WX11075), .Q(n3254) );
  XNOR3X1 U4982 ( .IN1(n3258), .IN2(n4751), .IN3(n3351), .Q(n2217) );
  XOR3X1 U4983 ( .IN1(WX11201), .IN2(test_so95), .IN3(WX11073), .Q(n3258) );
  XNOR3X1 U4984 ( .IN1(n3260), .IN2(n4751), .IN3(n3352), .Q(n2220) );
  XOR3X1 U4985 ( .IN1(WX11199), .IN2(WX11135), .IN3(WX11071), .Q(n3260) );
  XNOR3X1 U4986 ( .IN1(n3262), .IN2(n4751), .IN3(n3353), .Q(n2223) );
  XOR3X1 U4987 ( .IN1(WX11197), .IN2(WX11133), .IN3(test_so93), .Q(n3262) );
  XNOR3X1 U4988 ( .IN1(n3264), .IN2(n4751), .IN3(n3354), .Q(n2226) );
  XOR3X1 U4989 ( .IN1(WX11195), .IN2(WX11131), .IN3(WX11067), .Q(n3264) );
  XNOR3X1 U4990 ( .IN1(n3266), .IN2(n4751), .IN3(n3355), .Q(n2229) );
  XOR3X1 U4991 ( .IN1(WX11193), .IN2(WX11129), .IN3(WX11065), .Q(n3266) );
  XNOR3X1 U4992 ( .IN1(n3268), .IN2(n4751), .IN3(n3356), .Q(n2232) );
  XOR3X1 U4993 ( .IN1(WX11191), .IN2(WX11127), .IN3(WX11063), .Q(n3268) );
  XNOR3X1 U4994 ( .IN1(n3270), .IN2(n4751), .IN3(n3357), .Q(n2235) );
  XOR3X1 U4995 ( .IN1(WX11189), .IN2(WX11125), .IN3(WX11061), .Q(n3270) );
  XNOR3X1 U4996 ( .IN1(n3272), .IN2(n4751), .IN3(n3358), .Q(n2238) );
  XOR3X1 U4997 ( .IN1(WX11187), .IN2(WX11123), .IN3(WX11059), .Q(n3272) );
  XNOR3X1 U4998 ( .IN1(n3274), .IN2(n4751), .IN3(n3359), .Q(n2241) );
  XOR3X1 U4999 ( .IN1(WX11185), .IN2(WX11121), .IN3(WX11057), .Q(n3274) );
  XNOR3X1 U5000 ( .IN1(n3276), .IN2(n4751), .IN3(n3360), .Q(n2244) );
  XOR3X1 U5001 ( .IN1(WX11183), .IN2(WX11119), .IN3(WX11055), .Q(n3276) );
  XNOR3X1 U5002 ( .IN1(n2331), .IN2(n4748), .IN3(n3361), .Q(n2200) );
  XOR3X1 U5003 ( .IN1(WX9918), .IN2(test_so84), .IN3(WX9790), .Q(n2331) );
  XNOR3X1 U5004 ( .IN1(n2334), .IN2(n4743), .IN3(n3362), .Q(n2203) );
  XOR3X1 U5005 ( .IN1(WX9916), .IN2(WX9852), .IN3(WX9788), .Q(n2334) );
  XNOR3X1 U5006 ( .IN1(n2337), .IN2(n4743), .IN3(n3363), .Q(n2206) );
  XOR3X1 U5007 ( .IN1(WX9914), .IN2(WX9850), .IN3(test_so82), .Q(n2337) );
  XNOR3X1 U5008 ( .IN1(n2340), .IN2(n4743), .IN3(n3364), .Q(n2209) );
  XOR3X1 U5009 ( .IN1(WX9912), .IN2(WX9848), .IN3(WX9784), .Q(n2340) );
  XNOR3X1 U5010 ( .IN1(n2343), .IN2(n4743), .IN3(n3365), .Q(n2212) );
  XOR3X1 U5011 ( .IN1(WX9910), .IN2(WX9846), .IN3(WX9782), .Q(n2343) );
  XNOR3X1 U5012 ( .IN1(n2346), .IN2(n4743), .IN3(n3366), .Q(n2215) );
  XOR3X1 U5013 ( .IN1(WX9908), .IN2(WX9844), .IN3(WX9780), .Q(n2346) );
  XNOR3X1 U5014 ( .IN1(n2349), .IN2(n4743), .IN3(n3367), .Q(n2218) );
  XOR3X1 U5015 ( .IN1(WX9906), .IN2(WX9842), .IN3(WX9778), .Q(n2349) );
  XNOR3X1 U5016 ( .IN1(n2352), .IN2(n4743), .IN3(n3368), .Q(n2221) );
  XOR3X1 U5017 ( .IN1(WX9904), .IN2(WX9840), .IN3(WX9776), .Q(n2352) );
  XNOR3X1 U5018 ( .IN1(n2355), .IN2(n4743), .IN3(n3369), .Q(n2224) );
  XOR3X1 U5019 ( .IN1(WX9902), .IN2(WX9838), .IN3(WX9774), .Q(n2355) );
  XNOR3X1 U5020 ( .IN1(n2358), .IN2(n4743), .IN3(n3370), .Q(n2227) );
  XOR3X1 U5021 ( .IN1(WX9900), .IN2(WX9836), .IN3(WX9772), .Q(n2358) );
  XNOR3X1 U5022 ( .IN1(n2361), .IN2(n4743), .IN3(n3371), .Q(n2230) );
  XOR3X1 U5023 ( .IN1(WX9898), .IN2(WX9834), .IN3(WX9770), .Q(n2361) );
  XNOR3X1 U5024 ( .IN1(n2364), .IN2(n4743), .IN3(n3372), .Q(n2233) );
  XOR3X1 U5025 ( .IN1(WX9896), .IN2(WX9832), .IN3(WX9768), .Q(n2364) );
  XNOR3X1 U5026 ( .IN1(n2367), .IN2(n4743), .IN3(n3373), .Q(n2236) );
  XOR3X1 U5027 ( .IN1(WX9894), .IN2(WX9830), .IN3(WX9766), .Q(n2367) );
  XNOR3X1 U5028 ( .IN1(n2370), .IN2(n4744), .IN3(n3374), .Q(n2239) );
  XOR3X1 U5029 ( .IN1(WX9892), .IN2(WX9828), .IN3(WX9764), .Q(n2370) );
  XNOR3X1 U5030 ( .IN1(n2373), .IN2(n4744), .IN3(n3375), .Q(n2242) );
  XOR3X1 U5031 ( .IN1(WX9890), .IN2(WX9826), .IN3(WX9762), .Q(n2373) );
  XNOR3X1 U5032 ( .IN1(n2459), .IN2(n4744), .IN3(n3376), .Q(n2329) );
  XOR3X1 U5033 ( .IN1(WX8625), .IN2(WX8561), .IN3(WX8497), .Q(n2459) );
  XNOR3X1 U5034 ( .IN1(n2462), .IN2(n4744), .IN3(n3377), .Q(n2332) );
  XOR3X1 U5035 ( .IN1(WX8623), .IN2(WX8559), .IN3(WX8495), .Q(n2462) );
  XNOR3X1 U5036 ( .IN1(n2465), .IN2(n4744), .IN3(n3378), .Q(n2335) );
  XOR3X1 U5037 ( .IN1(WX8621), .IN2(WX8557), .IN3(WX8493), .Q(n2465) );
  XNOR3X1 U5038 ( .IN1(n2468), .IN2(n4744), .IN3(n3379), .Q(n2338) );
  XOR3X1 U5039 ( .IN1(WX8619), .IN2(WX8555), .IN3(WX8491), .Q(n2468) );
  XNOR3X1 U5040 ( .IN1(n2471), .IN2(n4744), .IN3(n3380), .Q(n2341) );
  XOR3X1 U5041 ( .IN1(WX8617), .IN2(WX8553), .IN3(WX8489), .Q(n2471) );
  XNOR3X1 U5042 ( .IN1(n2474), .IN2(n4744), .IN3(n3381), .Q(n2344) );
  XOR3X1 U5043 ( .IN1(WX8615), .IN2(WX8551), .IN3(WX8487), .Q(n2474) );
  XNOR3X1 U5044 ( .IN1(n2477), .IN2(n4744), .IN3(n3382), .Q(n2347) );
  XOR3X1 U5045 ( .IN1(WX8613), .IN2(WX8549), .IN3(WX8485), .Q(n2477) );
  XNOR3X1 U5046 ( .IN1(n2480), .IN2(n4744), .IN3(n3383), .Q(n2350) );
  XOR3X1 U5047 ( .IN1(WX8611), .IN2(WX8547), .IN3(WX8483), .Q(n2480) );
  XNOR3X1 U5048 ( .IN1(n2483), .IN2(n4744), .IN3(n3384), .Q(n2353) );
  XOR3X1 U5049 ( .IN1(WX8609), .IN2(WX8545), .IN3(WX8481), .Q(n2483) );
  XNOR3X1 U5050 ( .IN1(n2486), .IN2(n4744), .IN3(n3385), .Q(n2356) );
  XOR3X1 U5051 ( .IN1(WX8607), .IN2(WX8543), .IN3(WX8479), .Q(n2486) );
  XNOR3X1 U5052 ( .IN1(n2489), .IN2(n4745), .IN3(n3386), .Q(n2359) );
  XOR3X1 U5053 ( .IN1(test_so74), .IN2(WX8541), .IN3(WX8477), .Q(n2489) );
  XNOR3X1 U5054 ( .IN1(n2492), .IN2(n4745), .IN3(n3387), .Q(n2362) );
  XOR3X1 U5055 ( .IN1(WX8603), .IN2(WX8539), .IN3(WX8475), .Q(n2492) );
  XNOR3X1 U5056 ( .IN1(n2495), .IN2(n4745), .IN3(n3388), .Q(n2365) );
  XOR3X1 U5057 ( .IN1(WX8601), .IN2(test_so72), .IN3(WX8473), .Q(n2495) );
  XNOR3X1 U5058 ( .IN1(n2498), .IN2(n4745), .IN3(n3389), .Q(n2368) );
  XOR3X1 U5059 ( .IN1(WX8599), .IN2(WX8535), .IN3(WX8471), .Q(n2498) );
  XNOR3X1 U5060 ( .IN1(n2501), .IN2(n4745), .IN3(n3390), .Q(n2371) );
  XOR3X1 U5061 ( .IN1(WX8597), .IN2(WX8533), .IN3(test_so70), .Q(n2501) );
  XNOR3X1 U5062 ( .IN1(n2683), .IN2(n4745), .IN3(n3391), .Q(n2457) );
  XOR3X1 U5063 ( .IN1(WX7332), .IN2(WX7268), .IN3(WX7204), .Q(n2683) );
  XNOR3X1 U5064 ( .IN1(n2686), .IN2(n4745), .IN3(n3392), .Q(n2460) );
  XOR3X1 U5065 ( .IN1(WX7330), .IN2(WX7266), .IN3(WX7202), .Q(n2686) );
  XNOR3X1 U5066 ( .IN1(n2689), .IN2(n4745), .IN3(n3393), .Q(n2463) );
  XOR3X1 U5067 ( .IN1(WX7328), .IN2(WX7264), .IN3(WX7200), .Q(n2689) );
  XNOR3X1 U5068 ( .IN1(n2692), .IN2(n4745), .IN3(n3394), .Q(n2466) );
  XOR3X1 U5069 ( .IN1(WX7326), .IN2(WX7262), .IN3(WX7198), .Q(n2692) );
  XNOR3X1 U5070 ( .IN1(n2695), .IN2(n4745), .IN3(n3395), .Q(n2469) );
  XOR3X1 U5071 ( .IN1(WX7324), .IN2(WX7260), .IN3(WX7196), .Q(n2695) );
  XNOR3X1 U5072 ( .IN1(n2698), .IN2(n4745), .IN3(n3396), .Q(n2472) );
  XOR3X1 U5073 ( .IN1(test_so63), .IN2(WX7258), .IN3(WX7194), .Q(n2698) );
  XNOR3X1 U5074 ( .IN1(n2701), .IN2(n4745), .IN3(n3397), .Q(n2475) );
  XOR3X1 U5075 ( .IN1(WX7320), .IN2(WX7256), .IN3(WX7192), .Q(n2701) );
  XNOR3X1 U5076 ( .IN1(n2704), .IN2(n4746), .IN3(n3398), .Q(n2478) );
  XOR3X1 U5077 ( .IN1(WX7318), .IN2(test_so61), .IN3(WX7190), .Q(n2704) );
  XNOR3X1 U5078 ( .IN1(n2707), .IN2(n4746), .IN3(n3399), .Q(n2481) );
  XOR3X1 U5079 ( .IN1(WX7316), .IN2(WX7252), .IN3(WX7188), .Q(n2707) );
  XNOR3X1 U5080 ( .IN1(n2710), .IN2(n4746), .IN3(n3400), .Q(n2484) );
  XOR3X1 U5081 ( .IN1(WX7314), .IN2(WX7250), .IN3(test_so59), .Q(n2710) );
  XNOR3X1 U5082 ( .IN1(n2713), .IN2(n4746), .IN3(n3401), .Q(n2487) );
  XOR3X1 U5083 ( .IN1(WX7312), .IN2(WX7248), .IN3(WX7184), .Q(n2713) );
  XNOR3X1 U5084 ( .IN1(n2716), .IN2(n4746), .IN3(n3402), .Q(n2490) );
  XOR3X1 U5085 ( .IN1(WX7310), .IN2(WX7246), .IN3(WX7182), .Q(n2716) );
  XNOR3X1 U5086 ( .IN1(n2719), .IN2(n4746), .IN3(n3403), .Q(n2493) );
  XOR3X1 U5087 ( .IN1(WX7308), .IN2(WX7244), .IN3(WX7180), .Q(n2719) );
  XNOR3X1 U5088 ( .IN1(n2722), .IN2(n4746), .IN3(n3404), .Q(n2496) );
  XOR3X1 U5089 ( .IN1(WX7306), .IN2(WX7242), .IN3(WX7178), .Q(n2722) );
  XNOR3X1 U5090 ( .IN1(n2725), .IN2(n4746), .IN3(n3405), .Q(n2499) );
  XOR3X1 U5091 ( .IN1(WX7304), .IN2(WX7240), .IN3(WX7176), .Q(n2725) );
  XNOR3X1 U5092 ( .IN1(n2811), .IN2(n4746), .IN3(n3406), .Q(n2681) );
  XOR3X1 U5093 ( .IN1(test_so52), .IN2(WX5975), .IN3(WX5911), .Q(n2811) );
  XNOR3X1 U5094 ( .IN1(n2814), .IN2(n4746), .IN3(n3407), .Q(n2684) );
  XOR3X1 U5095 ( .IN1(WX6037), .IN2(WX5973), .IN3(WX5909), .Q(n2814) );
  XNOR3X1 U5096 ( .IN1(n2817), .IN2(n4746), .IN3(n3408), .Q(n2687) );
  XOR3X1 U5097 ( .IN1(WX6035), .IN2(test_so50), .IN3(WX5907), .Q(n2817) );
  XNOR3X1 U5098 ( .IN1(n2820), .IN2(n4746), .IN3(n3409), .Q(n2690) );
  XOR3X1 U5099 ( .IN1(WX6033), .IN2(WX5969), .IN3(WX5905), .Q(n2820) );
  XNOR3X1 U5100 ( .IN1(n2823), .IN2(n4747), .IN3(n3410), .Q(n2693) );
  XOR3X1 U5101 ( .IN1(WX6031), .IN2(WX5967), .IN3(test_so48), .Q(n2823) );
  XNOR3X1 U5102 ( .IN1(n2826), .IN2(n4747), .IN3(n3411), .Q(n2696) );
  XOR3X1 U5103 ( .IN1(WX6029), .IN2(WX5965), .IN3(WX5901), .Q(n2826) );
  XNOR3X1 U5104 ( .IN1(n2829), .IN2(n4747), .IN3(n3412), .Q(n2699) );
  XOR3X1 U5105 ( .IN1(WX6027), .IN2(WX5963), .IN3(WX5899), .Q(n2829) );
  XNOR3X1 U5106 ( .IN1(n2832), .IN2(n4747), .IN3(n3413), .Q(n2702) );
  XOR3X1 U5107 ( .IN1(WX6025), .IN2(WX5961), .IN3(WX5897), .Q(n2832) );
  XNOR3X1 U5108 ( .IN1(n2835), .IN2(n4747), .IN3(n3414), .Q(n2705) );
  XOR3X1 U5109 ( .IN1(WX6023), .IN2(WX5959), .IN3(WX5895), .Q(n2835) );
  XNOR3X1 U5110 ( .IN1(n2838), .IN2(n4747), .IN3(n3415), .Q(n2708) );
  XOR3X1 U5111 ( .IN1(WX6021), .IN2(WX5957), .IN3(WX5893), .Q(n2838) );
  XNOR3X1 U5112 ( .IN1(n2841), .IN2(n4747), .IN3(n3416), .Q(n2711) );
  XOR3X1 U5113 ( .IN1(WX6019), .IN2(WX5955), .IN3(WX5891), .Q(n2841) );
  XNOR3X1 U5114 ( .IN1(n2844), .IN2(n4747), .IN3(n3417), .Q(n2714) );
  XOR3X1 U5115 ( .IN1(WX6017), .IN2(WX5953), .IN3(WX5889), .Q(n2844) );
  XNOR3X1 U5116 ( .IN1(n2847), .IN2(n4747), .IN3(n3418), .Q(n2717) );
  XOR3X1 U5117 ( .IN1(WX6015), .IN2(WX5951), .IN3(WX5887), .Q(n2847) );
  XNOR3X1 U5118 ( .IN1(n2850), .IN2(n4747), .IN3(n3419), .Q(n2720) );
  XOR3X1 U5119 ( .IN1(WX6013), .IN2(WX5949), .IN3(WX5885), .Q(n2850) );
  XNOR3X1 U5120 ( .IN1(n2853), .IN2(n4747), .IN3(n3420), .Q(n2723) );
  XOR3X1 U5121 ( .IN1(WX6011), .IN2(WX5947), .IN3(WX5883), .Q(n2853) );
  XNOR3X1 U5122 ( .IN1(n2939), .IN2(n4747), .IN3(n3421), .Q(n2809) );
  XOR3X1 U5123 ( .IN1(WX4746), .IN2(WX4682), .IN3(WX4618), .Q(n2939) );
  XNOR3X1 U5124 ( .IN1(n2942), .IN2(n4748), .IN3(n3422), .Q(n2812) );
  XOR3X1 U5125 ( .IN1(WX4744), .IN2(WX4680), .IN3(WX4616), .Q(n2942) );
  XNOR3X1 U5126 ( .IN1(n2945), .IN2(n4748), .IN3(n3423), .Q(n2815) );
  XOR3X1 U5127 ( .IN1(WX4742), .IN2(WX4678), .IN3(WX4614), .Q(n2945) );
  XNOR3X1 U5128 ( .IN1(n2948), .IN2(n4748), .IN3(n3424), .Q(n2818) );
  XOR3X1 U5129 ( .IN1(WX4740), .IN2(WX4676), .IN3(WX4612), .Q(n2948) );
  XNOR3X1 U5130 ( .IN1(n2951), .IN2(n4748), .IN3(n3425), .Q(n2821) );
  XOR3X1 U5131 ( .IN1(WX4738), .IN2(WX4674), .IN3(WX4610), .Q(n2951) );
  XNOR3X1 U5132 ( .IN1(n2954), .IN2(n4748), .IN3(n3426), .Q(n2824) );
  XOR3X1 U5133 ( .IN1(WX4736), .IN2(WX4672), .IN3(WX4608), .Q(n2954) );
  XNOR3X1 U5134 ( .IN1(n2957), .IN2(n4748), .IN3(n3427), .Q(n2827) );
  XOR3X1 U5135 ( .IN1(WX4734), .IN2(WX4670), .IN3(WX4606), .Q(n2957) );
  XNOR3X1 U5136 ( .IN1(n2960), .IN2(n4748), .IN3(n3428), .Q(n2830) );
  XOR3X1 U5137 ( .IN1(WX4732), .IN2(WX4668), .IN3(WX4604), .Q(n2960) );
  XNOR3X1 U5138 ( .IN1(n2963), .IN2(n4748), .IN3(n3429), .Q(n2833) );
  XOR3X1 U5139 ( .IN1(WX4730), .IN2(WX4666), .IN3(WX4602), .Q(n2963) );
  XNOR3X1 U5140 ( .IN1(n2966), .IN2(n4748), .IN3(n3430), .Q(n2836) );
  XOR3X1 U5141 ( .IN1(WX4728), .IN2(WX4664), .IN3(WX4600), .Q(n2966) );
  XNOR3X1 U5142 ( .IN1(n2969), .IN2(n4748), .IN3(n3431), .Q(n2839) );
  XOR3X1 U5143 ( .IN1(WX4726), .IN2(WX4662), .IN3(WX4598), .Q(n2969) );
  XNOR3X1 U5144 ( .IN1(n2972), .IN2(n4748), .IN3(n3432), .Q(n2842) );
  XOR3X1 U5145 ( .IN1(WX4724), .IN2(WX4660), .IN3(WX4596), .Q(n2972) );
  XNOR3X1 U5146 ( .IN1(n2975), .IN2(n4748), .IN3(n3433), .Q(n2845) );
  XOR3X1 U5147 ( .IN1(test_so40), .IN2(WX4658), .IN3(WX4594), .Q(n2975) );
  XNOR3X1 U5148 ( .IN1(n2978), .IN2(n4749), .IN3(n3434), .Q(n2848) );
  XOR3X1 U5149 ( .IN1(WX4720), .IN2(WX4656), .IN3(WX4592), .Q(n2978) );
  XNOR3X1 U5150 ( .IN1(n2981), .IN2(n4749), .IN3(n3435), .Q(n2851) );
  XOR3X1 U5151 ( .IN1(WX4718), .IN2(test_so38), .IN3(WX4590), .Q(n2981) );
  XNOR3X1 U5152 ( .IN1(n3066), .IN2(n4749), .IN3(n3436), .Q(n2937) );
  XOR3X1 U5153 ( .IN1(WX3453), .IN2(WX3389), .IN3(WX3325), .Q(n3066) );
  XNOR3X1 U5154 ( .IN1(n3069), .IN2(n4749), .IN3(n3437), .Q(n2940) );
  XOR3X1 U5155 ( .IN1(WX3451), .IN2(WX3387), .IN3(WX3323), .Q(n3069) );
  XNOR3X1 U5156 ( .IN1(n3072), .IN2(n4749), .IN3(n3438), .Q(n2943) );
  XOR3X1 U5157 ( .IN1(WX3449), .IN2(WX3385), .IN3(WX3321), .Q(n3072) );
  XNOR3X1 U5158 ( .IN1(n3075), .IN2(n4749), .IN3(n3439), .Q(n2946) );
  XOR3X1 U5159 ( .IN1(WX3447), .IN2(WX3383), .IN3(WX3319), .Q(n3075) );
  XNOR3X1 U5160 ( .IN1(n3078), .IN2(n4749), .IN3(n3440), .Q(n2949) );
  XOR3X1 U5161 ( .IN1(WX3445), .IN2(WX3381), .IN3(WX3317), .Q(n3078) );
  XNOR3X1 U5162 ( .IN1(n3081), .IN2(n4750), .IN3(n3441), .Q(n2952) );
  XOR3X1 U5163 ( .IN1(WX3443), .IN2(WX3379), .IN3(WX3315), .Q(n3081) );
  XNOR3X1 U5164 ( .IN1(n3084), .IN2(n4750), .IN3(n3442), .Q(n2955) );
  XOR3X1 U5165 ( .IN1(WX3441), .IN2(WX3377), .IN3(WX3313), .Q(n3084) );
  XNOR3X1 U5166 ( .IN1(n3087), .IN2(n4750), .IN3(n3443), .Q(n2958) );
  XOR3X1 U5167 ( .IN1(test_so29), .IN2(WX3375), .IN3(WX3311), .Q(n3087) );
  XNOR3X1 U5168 ( .IN1(n3090), .IN2(n4750), .IN3(n3444), .Q(n2961) );
  XOR3X1 U5169 ( .IN1(WX3437), .IN2(WX3373), .IN3(WX3309), .Q(n3090) );
  XNOR3X1 U5170 ( .IN1(n3093), .IN2(n4750), .IN3(n3445), .Q(n2964) );
  XOR3X1 U5171 ( .IN1(WX3435), .IN2(WX3371), .IN3(WX3307), .Q(n3093) );
  XNOR3X1 U5172 ( .IN1(n3096), .IN2(n4750), .IN3(n3446), .Q(n2967) );
  XOR3X1 U5173 ( .IN1(WX3433), .IN2(test_so27), .IN3(WX3305), .Q(n3096) );
  XNOR3X1 U5174 ( .IN1(n3099), .IN2(n4750), .IN3(n3447), .Q(n2970) );
  XOR3X1 U5175 ( .IN1(WX3431), .IN2(WX3367), .IN3(WX3303), .Q(n3099) );
  XNOR3X1 U5176 ( .IN1(n3102), .IN2(n4762), .IN3(n3448), .Q(n2973) );
  XOR3X1 U5177 ( .IN1(WX3429), .IN2(WX3365), .IN3(WX3301), .Q(n3102) );
  XNOR3X1 U5178 ( .IN1(n3105), .IN2(n4763), .IN3(n3449), .Q(n2976) );
  XOR3X1 U5179 ( .IN1(WX3427), .IN2(WX3363), .IN3(WX3299), .Q(n3105) );
  XNOR3X1 U5180 ( .IN1(n3108), .IN2(n4762), .IN3(n3450), .Q(n2979) );
  XOR3X1 U5181 ( .IN1(WX3425), .IN2(WX3361), .IN3(test_so25), .Q(n3108) );
  XNOR3X1 U5182 ( .IN1(n3067), .IN2(n4749), .IN3(n3451), .Q(n2555) );
  XOR3X1 U5183 ( .IN1(WX2160), .IN2(WX2096), .IN3(WX2032), .Q(n3067) );
  XNOR3X1 U5184 ( .IN1(n3070), .IN2(n4749), .IN3(n3452), .Q(n2558) );
  XOR3X1 U5185 ( .IN1(WX2158), .IN2(WX2094), .IN3(WX2030), .Q(n3070) );
  XNOR3X1 U5186 ( .IN1(n3073), .IN2(n4749), .IN3(n3453), .Q(n2561) );
  XOR3X1 U5187 ( .IN1(WX2156), .IN2(WX2092), .IN3(test_so15), .Q(n3073) );
  XNOR3X1 U5188 ( .IN1(n3076), .IN2(n4749), .IN3(n3454), .Q(n2564) );
  XOR3X1 U5189 ( .IN1(WX2154), .IN2(WX2090), .IN3(WX2026), .Q(n3076) );
  XNOR3X1 U5190 ( .IN1(n3079), .IN2(n4749), .IN3(n3455), .Q(n2567) );
  XOR3X1 U5191 ( .IN1(WX2152), .IN2(WX2088), .IN3(WX2024), .Q(n3079) );
  XNOR3X1 U5192 ( .IN1(n3082), .IN2(n4750), .IN3(n3456), .Q(n2570) );
  XOR3X1 U5193 ( .IN1(WX2150), .IN2(WX2086), .IN3(WX2022), .Q(n3082) );
  XNOR3X1 U5194 ( .IN1(n3085), .IN2(n4750), .IN3(n3457), .Q(n2573) );
  XOR3X1 U5195 ( .IN1(WX2148), .IN2(WX2084), .IN3(WX2020), .Q(n3085) );
  XNOR3X1 U5196 ( .IN1(n3088), .IN2(n4750), .IN3(n3458), .Q(n2576) );
  XOR3X1 U5197 ( .IN1(WX2146), .IN2(WX2082), .IN3(WX2018), .Q(n3088) );
  XNOR3X1 U5198 ( .IN1(n3091), .IN2(n4750), .IN3(n3459), .Q(n2579) );
  XOR3X1 U5199 ( .IN1(WX2144), .IN2(WX2080), .IN3(WX2016), .Q(n3091) );
  XNOR3X1 U5200 ( .IN1(n3094), .IN2(n4750), .IN3(n3460), .Q(n2582) );
  XOR3X1 U5201 ( .IN1(WX2142), .IN2(WX2078), .IN3(WX2014), .Q(n3094) );
  XNOR3X1 U5202 ( .IN1(n3097), .IN2(n4750), .IN3(n3461), .Q(n2585) );
  XOR3X1 U5203 ( .IN1(WX2140), .IN2(WX2076), .IN3(WX2012), .Q(n3097) );
  XNOR3X1 U5204 ( .IN1(n3100), .IN2(n4764), .IN3(n3462), .Q(n2588) );
  XOR3X1 U5205 ( .IN1(WX2138), .IN2(WX2074), .IN3(WX2010), .Q(n3100) );
  XNOR3X1 U5206 ( .IN1(n3103), .IN2(n4764), .IN3(n3463), .Q(n2591) );
  XOR3X1 U5207 ( .IN1(test_so18), .IN2(WX2072), .IN3(WX2008), .Q(n3103) );
  XNOR3X1 U5208 ( .IN1(n3106), .IN2(n4750), .IN3(n3464), .Q(n2604) );
  XOR3X1 U5209 ( .IN1(WX2134), .IN2(WX2070), .IN3(WX2006), .Q(n3106) );
  XNOR3X1 U5210 ( .IN1(n3109), .IN2(n4764), .IN3(n3465), .Q(n2617) );
  XOR3X1 U5211 ( .IN1(WX2132), .IN2(WX2068), .IN3(WX2004), .Q(n3109) );
  XOR3X1 U5212 ( .IN1(n3530), .IN2(n3531), .IN3(WX11051), .Q(n2154) );
  XNOR2X1 U5213 ( .IN1(WX11243), .IN2(WX11179), .Q(n3530) );
  XOR3X1 U5214 ( .IN1(n3532), .IN2(n3533), .IN3(WX11049), .Q(n2157) );
  XNOR2X1 U5215 ( .IN1(WX11241), .IN2(WX11177), .Q(n3532) );
  XOR3X1 U5216 ( .IN1(n3534), .IN2(n3535), .IN3(WX11047), .Q(n2160) );
  XNOR2X1 U5217 ( .IN1(test_so98), .IN2(WX11175), .Q(n3534) );
  XOR3X1 U5218 ( .IN1(n3536), .IN2(n3537), .IN3(WX11045), .Q(n2163) );
  XNOR2X1 U5219 ( .IN1(WX11237), .IN2(WX11173), .Q(n3536) );
  XOR3X1 U5220 ( .IN1(n3538), .IN2(n3539), .IN3(WX11043), .Q(n2166) );
  XNOR2X1 U5221 ( .IN1(WX11235), .IN2(test_so96), .Q(n3538) );
  XOR3X1 U5222 ( .IN1(n3540), .IN2(n3541), .IN3(WX11041), .Q(n2169) );
  XNOR2X1 U5223 ( .IN1(WX11233), .IN2(WX11169), .Q(n3540) );
  XOR3X1 U5224 ( .IN1(n3542), .IN2(n3543), .IN3(WX11039), .Q(n2172) );
  XNOR2X1 U5225 ( .IN1(WX11231), .IN2(WX11167), .Q(n3542) );
  XOR3X1 U5226 ( .IN1(n3544), .IN2(n3545), .IN3(WX11037), .Q(n2175) );
  XNOR2X1 U5227 ( .IN1(WX11229), .IN2(WX11165), .Q(n3544) );
  XOR3X1 U5228 ( .IN1(n3546), .IN2(n3547), .IN3(test_so92), .Q(n2178) );
  XNOR2X1 U5229 ( .IN1(WX11227), .IN2(WX11163), .Q(n3546) );
  XOR3X1 U5230 ( .IN1(n3548), .IN2(n3549), .IN3(WX11033), .Q(n2181) );
  XNOR2X1 U5231 ( .IN1(WX11225), .IN2(WX11161), .Q(n3548) );
  XOR3X1 U5232 ( .IN1(n3550), .IN2(n3551), .IN3(WX11031), .Q(n2184) );
  XNOR2X1 U5233 ( .IN1(WX11223), .IN2(WX11159), .Q(n3550) );
  XOR3X1 U5234 ( .IN1(n3552), .IN2(n3553), .IN3(WX11029), .Q(n2187) );
  XNOR2X1 U5235 ( .IN1(WX11221), .IN2(WX11157), .Q(n3552) );
  XOR3X1 U5236 ( .IN1(n3554), .IN2(n3555), .IN3(WX11027), .Q(n2190) );
  XNOR2X1 U5237 ( .IN1(WX11219), .IN2(WX11155), .Q(n3554) );
  XOR3X1 U5238 ( .IN1(n3556), .IN2(n3557), .IN3(WX11025), .Q(n2193) );
  XNOR2X1 U5239 ( .IN1(WX11217), .IN2(WX11153), .Q(n3556) );
  XOR3X1 U5240 ( .IN1(n3558), .IN2(n3559), .IN3(WX11023), .Q(n2196) );
  XNOR2X1 U5241 ( .IN1(WX11215), .IN2(WX11151), .Q(n3558) );
  XOR3X1 U5242 ( .IN1(n3560), .IN2(n3561), .IN3(WX11021), .Q(n2199) );
  XNOR2X1 U5243 ( .IN1(WX11213), .IN2(WX11149), .Q(n3560) );
  XOR3X1 U5244 ( .IN1(n3562), .IN2(n3563), .IN3(WX9758), .Q(n2150) );
  XNOR2X1 U5245 ( .IN1(WX9950), .IN2(WX9886), .Q(n3562) );
  XOR3X1 U5246 ( .IN1(n3564), .IN2(n3565), .IN3(WX9756), .Q(n2155) );
  XNOR2X1 U5247 ( .IN1(WX9948), .IN2(WX9884), .Q(n3564) );
  XOR3X1 U5248 ( .IN1(n3566), .IN2(n3567), .IN3(WX9754), .Q(n2158) );
  XNOR2X1 U5249 ( .IN1(WX9946), .IN2(WX9882), .Q(n3566) );
  XOR3X1 U5250 ( .IN1(n3568), .IN2(n3569), .IN3(test_so81), .Q(n2161) );
  XNOR2X1 U5251 ( .IN1(WX9944), .IN2(WX9880), .Q(n3568) );
  XOR3X1 U5252 ( .IN1(n3570), .IN2(n3571), .IN3(WX9750), .Q(n2164) );
  XNOR2X1 U5253 ( .IN1(WX9942), .IN2(WX9878), .Q(n3570) );
  XOR3X1 U5254 ( .IN1(n3572), .IN2(n3573), .IN3(WX9748), .Q(n2167) );
  XNOR2X1 U5255 ( .IN1(WX9940), .IN2(WX9876), .Q(n3572) );
  XOR3X1 U5256 ( .IN1(n3574), .IN2(n3575), .IN3(WX9746), .Q(n2170) );
  XNOR2X1 U5257 ( .IN1(WX9938), .IN2(WX9874), .Q(n3574) );
  XOR3X1 U5258 ( .IN1(n3576), .IN2(n3577), .IN3(WX9744), .Q(n2173) );
  XNOR2X1 U5259 ( .IN1(WX9936), .IN2(WX9872), .Q(n3576) );
  XOR3X1 U5260 ( .IN1(n3578), .IN2(n3579), .IN3(WX9742), .Q(n2176) );
  XNOR2X1 U5261 ( .IN1(WX9934), .IN2(WX9870), .Q(n3578) );
  XOR3X1 U5262 ( .IN1(n3580), .IN2(n3581), .IN3(WX9740), .Q(n2179) );
  XNOR2X1 U5263 ( .IN1(WX9932), .IN2(WX9868), .Q(n3580) );
  XOR3X1 U5264 ( .IN1(n3582), .IN2(n3583), .IN3(WX9738), .Q(n2182) );
  XNOR2X1 U5265 ( .IN1(WX9930), .IN2(WX9866), .Q(n3582) );
  XOR3X1 U5266 ( .IN1(n3584), .IN2(n3585), .IN3(WX9736), .Q(n2185) );
  XNOR2X1 U5267 ( .IN1(WX9928), .IN2(WX9864), .Q(n3584) );
  XOR3X1 U5268 ( .IN1(n3586), .IN2(n3587), .IN3(WX9734), .Q(n2188) );
  XNOR2X1 U5269 ( .IN1(WX9926), .IN2(WX9862), .Q(n3586) );
  XOR3X1 U5270 ( .IN1(n3588), .IN2(n3589), .IN3(WX9732), .Q(n2191) );
  XNOR2X1 U5271 ( .IN1(WX9924), .IN2(WX9860), .Q(n3588) );
  XOR3X1 U5272 ( .IN1(n3590), .IN2(n3591), .IN3(WX9730), .Q(n2194) );
  XNOR2X1 U5273 ( .IN1(test_so86), .IN2(WX9858), .Q(n3590) );
  XOR3X1 U5274 ( .IN1(n3592), .IN2(n3593), .IN3(WX9728), .Q(n2197) );
  XNOR2X1 U5275 ( .IN1(WX9920), .IN2(WX9856), .Q(n3592) );
  XOR3X1 U5276 ( .IN1(n3594), .IN2(n3595), .IN3(WX8465), .Q(n2281) );
  XNOR2X1 U5277 ( .IN1(WX8657), .IN2(WX8593), .Q(n3594) );
  XOR3X1 U5278 ( .IN1(n3596), .IN2(n3597), .IN3(WX8463), .Q(n2284) );
  XNOR2X1 U5279 ( .IN1(WX8655), .IN2(WX8591), .Q(n3596) );
  XOR3X1 U5280 ( .IN1(n3598), .IN2(n3599), .IN3(WX8461), .Q(n2287) );
  XNOR2X1 U5281 ( .IN1(WX8653), .IN2(WX8589), .Q(n3598) );
  XOR3X1 U5282 ( .IN1(n3600), .IN2(n3601), .IN3(WX8459), .Q(n2290) );
  XNOR2X1 U5283 ( .IN1(WX8651), .IN2(WX8587), .Q(n3600) );
  XOR3X1 U5284 ( .IN1(n3602), .IN2(n3603), .IN3(WX8457), .Q(n2293) );
  XNOR2X1 U5285 ( .IN1(WX8649), .IN2(WX8585), .Q(n3602) );
  XOR3X1 U5286 ( .IN1(n3604), .IN2(n3605), .IN3(WX8455), .Q(n2296) );
  XNOR2X1 U5287 ( .IN1(WX8647), .IN2(WX8583), .Q(n3604) );
  XOR3X1 U5288 ( .IN1(n3606), .IN2(n3607), .IN3(WX8453), .Q(n2299) );
  XNOR2X1 U5289 ( .IN1(WX8645), .IN2(WX8581), .Q(n3606) );
  XOR3X1 U5290 ( .IN1(n3608), .IN2(n3609), .IN3(WX8451), .Q(n2302) );
  XNOR2X1 U5291 ( .IN1(WX8643), .IN2(WX8579), .Q(n3608) );
  XOR3X1 U5292 ( .IN1(n3610), .IN2(n3611), .IN3(WX8449), .Q(n2305) );
  XNOR2X1 U5293 ( .IN1(WX8641), .IN2(WX8577), .Q(n3610) );
  XOR3X1 U5294 ( .IN1(n3612), .IN2(n3613), .IN3(WX8447), .Q(n2308) );
  XNOR2X1 U5295 ( .IN1(test_so75), .IN2(WX8575), .Q(n3612) );
  XOR3X1 U5296 ( .IN1(n3614), .IN2(n3615), .IN3(WX8445), .Q(n2311) );
  XNOR2X1 U5297 ( .IN1(WX8637), .IN2(WX8573), .Q(n3614) );
  XOR3X1 U5298 ( .IN1(n3616), .IN2(n3617), .IN3(WX8443), .Q(n2314) );
  XNOR2X1 U5299 ( .IN1(WX8635), .IN2(test_so73), .Q(n3616) );
  XOR3X1 U5300 ( .IN1(n3618), .IN2(n3619), .IN3(WX8441), .Q(n2317) );
  XNOR2X1 U5301 ( .IN1(WX8633), .IN2(WX8569), .Q(n3618) );
  XOR3X1 U5302 ( .IN1(n3620), .IN2(n3621), .IN3(WX8439), .Q(n2320) );
  XNOR2X1 U5303 ( .IN1(WX8631), .IN2(WX8567), .Q(n3620) );
  XOR3X1 U5304 ( .IN1(n3622), .IN2(n3623), .IN3(WX8437), .Q(n2323) );
  XNOR2X1 U5305 ( .IN1(WX8629), .IN2(WX8565), .Q(n3622) );
  XOR3X1 U5306 ( .IN1(n3624), .IN2(n3625), .IN3(test_so69), .Q(n2326) );
  XNOR2X1 U5307 ( .IN1(WX8627), .IN2(WX8563), .Q(n3624) );
  XOR3X1 U5308 ( .IN1(n3626), .IN2(n3627), .IN3(WX7172), .Q(n2409) );
  XNOR2X1 U5309 ( .IN1(WX7364), .IN2(WX7300), .Q(n3626) );
  XOR3X1 U5310 ( .IN1(n3628), .IN2(n3629), .IN3(WX7170), .Q(n2412) );
  XNOR2X1 U5311 ( .IN1(WX7362), .IN2(WX7298), .Q(n3628) );
  XOR3X1 U5312 ( .IN1(n3630), .IN2(n3631), .IN3(WX7168), .Q(n2415) );
  XNOR2X1 U5313 ( .IN1(WX7360), .IN2(WX7296), .Q(n3630) );
  XOR3X1 U5314 ( .IN1(n3632), .IN2(n3633), .IN3(WX7166), .Q(n2418) );
  XNOR2X1 U5315 ( .IN1(WX7358), .IN2(WX7294), .Q(n3632) );
  XOR3X1 U5316 ( .IN1(n3634), .IN2(n3635), .IN3(WX7164), .Q(n2421) );
  XNOR2X1 U5317 ( .IN1(test_so64), .IN2(WX7292), .Q(n3634) );
  XOR3X1 U5318 ( .IN1(n3636), .IN2(n3637), .IN3(WX7162), .Q(n2424) );
  XNOR2X1 U5319 ( .IN1(WX7354), .IN2(WX7290), .Q(n3636) );
  XOR3X1 U5320 ( .IN1(n3638), .IN2(n3639), .IN3(WX7160), .Q(n2427) );
  XNOR2X1 U5321 ( .IN1(WX7352), .IN2(test_so62), .Q(n3638) );
  XOR3X1 U5322 ( .IN1(n3640), .IN2(n3641), .IN3(WX7158), .Q(n2430) );
  XNOR2X1 U5323 ( .IN1(WX7350), .IN2(WX7286), .Q(n3640) );
  XOR3X1 U5324 ( .IN1(n3642), .IN2(n3643), .IN3(WX7156), .Q(n2433) );
  XNOR2X1 U5325 ( .IN1(WX7348), .IN2(WX7284), .Q(n3642) );
  XOR3X1 U5326 ( .IN1(n3644), .IN2(n3645), .IN3(WX7154), .Q(n2436) );
  XNOR2X1 U5327 ( .IN1(WX7346), .IN2(WX7282), .Q(n3644) );
  XOR3X1 U5328 ( .IN1(n3646), .IN2(n3647), .IN3(test_so58), .Q(n2439) );
  XNOR2X1 U5329 ( .IN1(WX7344), .IN2(WX7280), .Q(n3646) );
  XOR3X1 U5330 ( .IN1(n3648), .IN2(n3649), .IN3(WX7150), .Q(n2442) );
  XNOR2X1 U5331 ( .IN1(WX7342), .IN2(WX7278), .Q(n3648) );
  XOR3X1 U5332 ( .IN1(n3650), .IN2(n3651), .IN3(WX7148), .Q(n2445) );
  XNOR2X1 U5333 ( .IN1(WX7340), .IN2(WX7276), .Q(n3650) );
  XOR3X1 U5334 ( .IN1(n3652), .IN2(n3653), .IN3(WX7146), .Q(n2448) );
  XNOR2X1 U5335 ( .IN1(WX7338), .IN2(WX7274), .Q(n3652) );
  XOR3X1 U5336 ( .IN1(n3654), .IN2(n3655), .IN3(WX7144), .Q(n2451) );
  XNOR2X1 U5337 ( .IN1(WX7336), .IN2(WX7272), .Q(n3654) );
  XOR3X1 U5338 ( .IN1(n3656), .IN2(n3657), .IN3(WX7142), .Q(n2454) );
  XNOR2X1 U5339 ( .IN1(WX7334), .IN2(WX7270), .Q(n3656) );
  XOR3X1 U5340 ( .IN1(n3658), .IN2(n3659), .IN3(WX5879), .Q(n2633) );
  XNOR2X1 U5341 ( .IN1(WX6071), .IN2(WX6007), .Q(n3658) );
  XOR3X1 U5342 ( .IN1(n3660), .IN2(n3661), .IN3(WX5877), .Q(n2636) );
  XNOR2X1 U5343 ( .IN1(WX6069), .IN2(test_so51), .Q(n3660) );
  XOR3X1 U5344 ( .IN1(n3662), .IN2(n3663), .IN3(WX5875), .Q(n2639) );
  XNOR2X1 U5345 ( .IN1(WX6067), .IN2(WX6003), .Q(n3662) );
  XOR3X1 U5346 ( .IN1(n3664), .IN2(n3665), .IN3(WX5873), .Q(n2642) );
  XNOR2X1 U5347 ( .IN1(WX6065), .IN2(WX6001), .Q(n3664) );
  XOR3X1 U5348 ( .IN1(n3666), .IN2(n3667), .IN3(WX5871), .Q(n2645) );
  XNOR2X1 U5349 ( .IN1(WX6063), .IN2(WX5999), .Q(n3666) );
  XOR3X1 U5350 ( .IN1(n3668), .IN2(n3669), .IN3(test_so47), .Q(n2648) );
  XNOR2X1 U5351 ( .IN1(WX6061), .IN2(WX5997), .Q(n3668) );
  XOR3X1 U5352 ( .IN1(n3670), .IN2(n3671), .IN3(WX5867), .Q(n2651) );
  XNOR2X1 U5353 ( .IN1(WX6059), .IN2(WX5995), .Q(n3670) );
  XOR3X1 U5354 ( .IN1(n3672), .IN2(n3673), .IN3(WX5865), .Q(n2654) );
  XNOR2X1 U5355 ( .IN1(WX6057), .IN2(WX5993), .Q(n3672) );
  XOR3X1 U5356 ( .IN1(n3674), .IN2(n3675), .IN3(WX5863), .Q(n2657) );
  XNOR2X1 U5357 ( .IN1(WX6055), .IN2(WX5991), .Q(n3674) );
  XOR3X1 U5358 ( .IN1(n3676), .IN2(n3677), .IN3(WX5861), .Q(n2660) );
  XNOR2X1 U5359 ( .IN1(WX6053), .IN2(WX5989), .Q(n3676) );
  XOR3X1 U5360 ( .IN1(n3678), .IN2(n3679), .IN3(WX5859), .Q(n2663) );
  XNOR2X1 U5361 ( .IN1(WX6051), .IN2(WX5987), .Q(n3678) );
  XOR3X1 U5362 ( .IN1(n3680), .IN2(n3681), .IN3(WX5857), .Q(n2666) );
  XNOR2X1 U5363 ( .IN1(WX6049), .IN2(WX5985), .Q(n3680) );
  XOR3X1 U5364 ( .IN1(n3682), .IN2(n3683), .IN3(WX5855), .Q(n2669) );
  XNOR2X1 U5365 ( .IN1(WX6047), .IN2(WX5983), .Q(n3682) );
  XOR3X1 U5366 ( .IN1(n3684), .IN2(n3685), .IN3(WX5853), .Q(n2672) );
  XNOR2X1 U5367 ( .IN1(WX6045), .IN2(WX5981), .Q(n3684) );
  XOR3X1 U5368 ( .IN1(n3686), .IN2(n3687), .IN3(WX5851), .Q(n2675) );
  XNOR2X1 U5369 ( .IN1(WX6043), .IN2(WX5979), .Q(n3686) );
  XOR3X1 U5370 ( .IN1(n3688), .IN2(n3689), .IN3(WX5849), .Q(n2678) );
  XNOR2X1 U5371 ( .IN1(WX6041), .IN2(WX5977), .Q(n3688) );
  XOR3X1 U5372 ( .IN1(n3690), .IN2(n3691), .IN3(test_so36), .Q(n2761) );
  XNOR2X1 U5373 ( .IN1(WX4778), .IN2(WX4714), .Q(n3690) );
  XOR3X1 U5374 ( .IN1(n3692), .IN2(n3693), .IN3(WX4584), .Q(n2764) );
  XNOR2X1 U5375 ( .IN1(WX4776), .IN2(WX4712), .Q(n3692) );
  XOR3X1 U5376 ( .IN1(n3694), .IN2(n3695), .IN3(WX4582), .Q(n2767) );
  XNOR2X1 U5377 ( .IN1(WX4774), .IN2(WX4710), .Q(n3694) );
  XOR3X1 U5378 ( .IN1(n3696), .IN2(n3697), .IN3(WX4580), .Q(n2770) );
  XNOR2X1 U5379 ( .IN1(WX4772), .IN2(WX4708), .Q(n3696) );
  XOR3X1 U5380 ( .IN1(n3698), .IN2(n3699), .IN3(WX4578), .Q(n2773) );
  XNOR2X1 U5381 ( .IN1(WX4770), .IN2(WX4706), .Q(n3698) );
  XOR3X1 U5382 ( .IN1(n3700), .IN2(n3701), .IN3(WX4576), .Q(n2776) );
  XNOR2X1 U5383 ( .IN1(WX4768), .IN2(WX4704), .Q(n3700) );
  XOR3X1 U5384 ( .IN1(n3702), .IN2(n3703), .IN3(WX4574), .Q(n2779) );
  XNOR2X1 U5385 ( .IN1(WX4766), .IN2(WX4702), .Q(n3702) );
  XOR3X1 U5386 ( .IN1(n3704), .IN2(n3705), .IN3(WX4572), .Q(n2782) );
  XNOR2X1 U5387 ( .IN1(WX4764), .IN2(WX4700), .Q(n3704) );
  XOR3X1 U5388 ( .IN1(n3706), .IN2(n3707), .IN3(WX4570), .Q(n2785) );
  XNOR2X1 U5389 ( .IN1(WX4762), .IN2(WX4698), .Q(n3706) );
  XOR3X1 U5390 ( .IN1(n3708), .IN2(n3709), .IN3(WX4568), .Q(n2788) );
  XNOR2X1 U5391 ( .IN1(WX4760), .IN2(WX4696), .Q(n3708) );
  XOR3X1 U5392 ( .IN1(n3710), .IN2(n3711), .IN3(WX4566), .Q(n2791) );
  XNOR2X1 U5393 ( .IN1(WX4758), .IN2(WX4694), .Q(n3710) );
  XOR3X1 U5394 ( .IN1(n3712), .IN2(n3713), .IN3(WX4564), .Q(n2794) );
  XNOR2X1 U5395 ( .IN1(test_so41), .IN2(WX4692), .Q(n3712) );
  XOR3X1 U5396 ( .IN1(n3714), .IN2(n3715), .IN3(WX4562), .Q(n2797) );
  XNOR2X1 U5397 ( .IN1(WX4754), .IN2(WX4690), .Q(n3714) );
  XOR3X1 U5398 ( .IN1(n3716), .IN2(n3717), .IN3(WX4560), .Q(n2800) );
  XNOR2X1 U5399 ( .IN1(WX4752), .IN2(test_so39), .Q(n3716) );
  XOR3X1 U5400 ( .IN1(n3718), .IN2(n3719), .IN3(WX4558), .Q(n2803) );
  XNOR2X1 U5401 ( .IN1(WX4750), .IN2(WX4686), .Q(n3718) );
  XOR3X1 U5402 ( .IN1(n3720), .IN2(n3721), .IN3(WX4556), .Q(n2806) );
  XNOR2X1 U5403 ( .IN1(WX4748), .IN2(WX4684), .Q(n3720) );
  XOR3X1 U5404 ( .IN1(n3722), .IN2(n3723), .IN3(WX3293), .Q(n2889) );
  XNOR2X1 U5405 ( .IN1(WX3485), .IN2(WX3421), .Q(n3722) );
  XOR3X1 U5406 ( .IN1(n3724), .IN2(n3725), .IN3(WX3291), .Q(n2892) );
  XNOR2X1 U5407 ( .IN1(WX3483), .IN2(WX3419), .Q(n3724) );
  XOR3X1 U5408 ( .IN1(n3726), .IN2(n3727), .IN3(WX3289), .Q(n2895) );
  XNOR2X1 U5409 ( .IN1(WX3481), .IN2(WX3417), .Q(n3726) );
  XOR3X1 U5410 ( .IN1(n3728), .IN2(n3729), .IN3(WX3287), .Q(n2898) );
  XNOR2X1 U5411 ( .IN1(WX3479), .IN2(WX3415), .Q(n3728) );
  XOR3X1 U5412 ( .IN1(n3730), .IN2(n3731), .IN3(WX3285), .Q(n2901) );
  XNOR2X1 U5413 ( .IN1(WX3477), .IN2(WX3413), .Q(n3730) );
  XOR3X1 U5414 ( .IN1(n3732), .IN2(n3733), .IN3(WX3283), .Q(n2904) );
  XNOR2X1 U5415 ( .IN1(WX3475), .IN2(WX3411), .Q(n3732) );
  XOR3X1 U5416 ( .IN1(n3734), .IN2(n3735), .IN3(WX3281), .Q(n2907) );
  XNOR2X1 U5417 ( .IN1(test_so30), .IN2(WX3409), .Q(n3734) );
  XOR3X1 U5418 ( .IN1(n3736), .IN2(n3737), .IN3(WX3279), .Q(n2910) );
  XNOR2X1 U5419 ( .IN1(WX3471), .IN2(WX3407), .Q(n3736) );
  XOR3X1 U5420 ( .IN1(n3738), .IN2(n3739), .IN3(WX3277), .Q(n2913) );
  XNOR2X1 U5421 ( .IN1(WX3469), .IN2(test_so28), .Q(n3738) );
  XOR3X1 U5422 ( .IN1(n3740), .IN2(n3741), .IN3(WX3275), .Q(n2916) );
  XNOR2X1 U5423 ( .IN1(WX3467), .IN2(WX3403), .Q(n3740) );
  XOR3X1 U5424 ( .IN1(n3742), .IN2(n3743), .IN3(WX3273), .Q(n2919) );
  XNOR2X1 U5425 ( .IN1(WX3465), .IN2(WX3401), .Q(n3742) );
  XOR3X1 U5426 ( .IN1(n3744), .IN2(n3745), .IN3(WX3271), .Q(n2922) );
  XNOR2X1 U5427 ( .IN1(WX3463), .IN2(WX3399), .Q(n3744) );
  XOR3X1 U5428 ( .IN1(n3746), .IN2(n3747), .IN3(WX3269), .Q(n2925) );
  XNOR2X1 U5429 ( .IN1(WX3461), .IN2(WX3397), .Q(n3746) );
  XOR3X1 U5430 ( .IN1(n3748), .IN2(n3749), .IN3(WX3267), .Q(n2928) );
  XNOR2X1 U5431 ( .IN1(WX3459), .IN2(WX3395), .Q(n3748) );
  XOR3X1 U5432 ( .IN1(n3750), .IN2(n3751), .IN3(WX3265), .Q(n2931) );
  XNOR2X1 U5433 ( .IN1(WX3457), .IN2(WX3393), .Q(n3750) );
  XOR3X1 U5434 ( .IN1(n3752), .IN2(n3753), .IN3(WX3263), .Q(n2934) );
  XNOR2X1 U5435 ( .IN1(WX3455), .IN2(WX3391), .Q(n3752) );
  XOR3X1 U5436 ( .IN1(n3754), .IN2(n3755), .IN3(WX2000), .Q(n2507) );
  XNOR2X1 U5437 ( .IN1(WX2192), .IN2(WX2128), .Q(n3754) );
  XOR3X1 U5438 ( .IN1(n3756), .IN2(n3757), .IN3(WX1998), .Q(n2510) );
  XNOR2X1 U5439 ( .IN1(WX2190), .IN2(WX2126), .Q(n3756) );
  XOR3X1 U5440 ( .IN1(n3758), .IN2(n3759), .IN3(WX1996), .Q(n2513) );
  XNOR2X1 U5441 ( .IN1(WX2188), .IN2(WX2124), .Q(n3758) );
  XOR3X1 U5442 ( .IN1(n3760), .IN2(n3761), .IN3(WX1994), .Q(n2516) );
  XNOR2X1 U5443 ( .IN1(WX2186), .IN2(WX2122), .Q(n3760) );
  XOR3X1 U5444 ( .IN1(n3762), .IN2(n3763), .IN3(test_so14), .Q(n2519) );
  XNOR2X1 U5445 ( .IN1(WX2184), .IN2(WX2120), .Q(n3762) );
  XOR3X1 U5446 ( .IN1(n3764), .IN2(n3765), .IN3(WX1990), .Q(n2522) );
  XNOR2X1 U5447 ( .IN1(WX2182), .IN2(WX2118), .Q(n3764) );
  XOR3X1 U5448 ( .IN1(n3766), .IN2(n3767), .IN3(WX1988), .Q(n2525) );
  XNOR2X1 U5449 ( .IN1(WX2180), .IN2(WX2116), .Q(n3766) );
  XOR3X1 U5450 ( .IN1(n3768), .IN2(n3769), .IN3(WX1986), .Q(n2528) );
  XNOR2X1 U5451 ( .IN1(WX2178), .IN2(WX2114), .Q(n3768) );
  XOR3X1 U5452 ( .IN1(n3770), .IN2(n3771), .IN3(WX1984), .Q(n2531) );
  XNOR2X1 U5453 ( .IN1(WX2176), .IN2(WX2112), .Q(n3770) );
  XOR3X1 U5454 ( .IN1(n3772), .IN2(n3773), .IN3(WX1982), .Q(n2534) );
  XNOR2X1 U5455 ( .IN1(WX2174), .IN2(WX2110), .Q(n3772) );
  XOR3X1 U5456 ( .IN1(n3774), .IN2(n3775), .IN3(WX1980), .Q(n2537) );
  XNOR2X1 U5457 ( .IN1(test_so19), .IN2(WX2108), .Q(n3774) );
  XOR3X1 U5458 ( .IN1(n3776), .IN2(n3777), .IN3(WX1978), .Q(n2540) );
  XNOR2X1 U5459 ( .IN1(WX2170), .IN2(WX2106), .Q(n3776) );
  XOR3X1 U5460 ( .IN1(n3778), .IN2(n3779), .IN3(WX1976), .Q(n2543) );
  XNOR2X1 U5461 ( .IN1(WX2168), .IN2(WX2104), .Q(n3778) );
  XOR3X1 U5462 ( .IN1(n3780), .IN2(n3781), .IN3(WX1974), .Q(n2546) );
  XNOR2X1 U5463 ( .IN1(WX2166), .IN2(WX2102), .Q(n3780) );
  XOR3X1 U5464 ( .IN1(n3782), .IN2(n3783), .IN3(WX1972), .Q(n2549) );
  XNOR2X1 U5465 ( .IN1(WX2164), .IN2(test_so17), .Q(n3782) );
  XOR3X1 U5466 ( .IN1(n3784), .IN2(n3785), .IN3(WX1970), .Q(n2552) );
  XNOR2X1 U5467 ( .IN1(WX2162), .IN2(WX2098), .Q(n3784) );
  NOR2X0 U5468 ( .IN1(n3786), .IN2(n4586), .QN(WX10888) );
  NOR2X0 U5469 ( .IN1(n3787), .IN2(n4586), .QN(WX10886) );
  NOR2X0 U5470 ( .IN1(n3788), .IN2(n4586), .QN(WX10884) );
  NOR2X0 U5471 ( .IN1(n3789), .IN2(n4586), .QN(WX10882) );
  NOR2X0 U5472 ( .IN1(n3790), .IN2(n4586), .QN(WX10880) );
  NOR2X0 U5473 ( .IN1(n3791), .IN2(n4586), .QN(WX10878) );
  NOR2X0 U5474 ( .IN1(n3792), .IN2(n4586), .QN(WX10876) );
  NOR2X0 U5475 ( .IN1(n3793), .IN2(n4586), .QN(WX10874) );
  NOR2X0 U5476 ( .IN1(n3794), .IN2(n4586), .QN(WX10872) );
  NOR2X0 U5477 ( .IN1(n3795), .IN2(n4586), .QN(WX10870) );
  NOR2X0 U5478 ( .IN1(n3796), .IN2(n4587), .QN(WX10868) );
  NOR2X0 U5479 ( .IN1(n3797), .IN2(n4587), .QN(WX10866) );
  NOR2X0 U5480 ( .IN1(n3798), .IN2(n4587), .QN(WX10864) );
  NOR2X0 U5481 ( .IN1(n3799), .IN2(n4587), .QN(WX10862) );
  NOR2X0 U5482 ( .IN1(n3800), .IN2(n4587), .QN(WX10860) );
  NOR2X0 U5483 ( .IN1(n3801), .IN2(n4587), .QN(WX10858) );
  NOR2X0 U5484 ( .IN1(n3802), .IN2(n4587), .QN(WX10856) );
  NOR2X0 U5485 ( .IN1(n3803), .IN2(n4587), .QN(WX10854) );
  NOR2X0 U5486 ( .IN1(n3804), .IN2(n4587), .QN(WX10852) );
  NOR2X0 U5487 ( .IN1(n3805), .IN2(n4587), .QN(WX10850) );
  NOR2X0 U5488 ( .IN1(n3806), .IN2(n4587), .QN(WX10848) );
  NOR2X0 U5489 ( .IN1(n3807), .IN2(n4587), .QN(WX10846) );
  NOR2X0 U5490 ( .IN1(n3808), .IN2(n4587), .QN(WX10844) );
  NOR2X0 U5491 ( .IN1(n3809), .IN2(n4587), .QN(WX10842) );
  NOR2X0 U5492 ( .IN1(n3810), .IN2(n4587), .QN(WX10840) );
  NOR2X0 U5493 ( .IN1(n3811), .IN2(n4588), .QN(WX10838) );
  NOR2X0 U5494 ( .IN1(n3812), .IN2(n4588), .QN(WX10836) );
  NOR2X0 U5495 ( .IN1(n3813), .IN2(n4588), .QN(WX10834) );
  NOR2X0 U5496 ( .IN1(n3814), .IN2(n4588), .QN(WX10832) );
  NOR2X0 U5497 ( .IN1(n3815), .IN2(n4588), .QN(WX10830) );
  NOR2X0 U5498 ( .IN1(n3816), .IN2(n4588), .QN(WX10828) );
  NOR2X0 U5499 ( .IN1(n3817), .IN2(n4612), .QN(WX9595) );
  NOR2X0 U5500 ( .IN1(n3818), .IN2(n4612), .QN(WX9593) );
  NOR2X0 U5501 ( .IN1(n3819), .IN2(n4612), .QN(WX9591) );
  NOR2X0 U5502 ( .IN1(n3820), .IN2(n4612), .QN(WX9589) );
  NOR2X0 U5503 ( .IN1(n3821), .IN2(n4612), .QN(WX9587) );
  NOR2X0 U5504 ( .IN1(n3822), .IN2(n4612), .QN(WX9585) );
  NOR2X0 U5505 ( .IN1(n3823), .IN2(n4612), .QN(WX9583) );
  NOR2X0 U5506 ( .IN1(n3824), .IN2(n4612), .QN(WX9581) );
  NOR2X0 U5507 ( .IN1(n3825), .IN2(n4612), .QN(WX9579) );
  NOR2X0 U5508 ( .IN1(n3826), .IN2(n4613), .QN(WX9577) );
  NOR2X0 U5509 ( .IN1(n3827), .IN2(n4613), .QN(WX9575) );
  NOR2X0 U5510 ( .IN1(n3828), .IN2(n4613), .QN(WX9573) );
  NOR2X0 U5511 ( .IN1(n3829), .IN2(n4613), .QN(WX9571) );
  NOR2X0 U5512 ( .IN1(n3830), .IN2(n4613), .QN(WX9569) );
  NOR2X0 U5513 ( .IN1(n3831), .IN2(n4613), .QN(WX9567) );
  NOR2X0 U5514 ( .IN1(n3832), .IN2(n4613), .QN(WX9565) );
  NOR2X0 U5515 ( .IN1(n3833), .IN2(n4613), .QN(WX9563) );
  NOR2X0 U5516 ( .IN1(n3834), .IN2(n4613), .QN(WX9561) );
  NOR2X0 U5517 ( .IN1(n3835), .IN2(n4613), .QN(WX9559) );
  NOR2X0 U5518 ( .IN1(n3836), .IN2(n4613), .QN(WX9557) );
  NOR2X0 U5519 ( .IN1(n3837), .IN2(n4613), .QN(WX9555) );
  NOR2X0 U5520 ( .IN1(n3838), .IN2(n4613), .QN(WX9553) );
  NOR2X0 U5521 ( .IN1(n3839), .IN2(n4613), .QN(WX9551) );
  NOR2X0 U5522 ( .IN1(n3840), .IN2(n4613), .QN(WX9549) );
  NOR2X0 U5523 ( .IN1(n3841), .IN2(n4614), .QN(WX9547) );
  NOR2X0 U5524 ( .IN1(n3842), .IN2(n4614), .QN(WX9545) );
  NOR2X0 U5525 ( .IN1(n3843), .IN2(n4614), .QN(WX9543) );
  NOR2X0 U5526 ( .IN1(n3844), .IN2(n4614), .QN(WX9541) );
  NOR2X0 U5527 ( .IN1(n3845), .IN2(n4614), .QN(WX9539) );
  NOR2X0 U5528 ( .IN1(n3846), .IN2(n4614), .QN(WX9537) );
  NOR2X0 U5529 ( .IN1(n3847), .IN2(n4614), .QN(WX9535) );
  NOR2X0 U5530 ( .IN1(n3848), .IN2(n4601), .QN(WX8302) );
  NOR2X0 U5531 ( .IN1(n3849), .IN2(n4601), .QN(WX8300) );
  NOR2X0 U5532 ( .IN1(n3850), .IN2(n4601), .QN(WX8298) );
  NOR2X0 U5533 ( .IN1(n3851), .IN2(n4601), .QN(WX8296) );
  NOR2X0 U5534 ( .IN1(n3852), .IN2(n4601), .QN(WX8294) );
  NOR2X0 U5535 ( .IN1(n3853), .IN2(n4601), .QN(WX8292) );
  NOR2X0 U5536 ( .IN1(n3854), .IN2(n4601), .QN(WX8290) );
  NOR2X0 U5537 ( .IN1(n3855), .IN2(n4601), .QN(WX8288) );
  NOR2X0 U5538 ( .IN1(n3856), .IN2(n4601), .QN(WX8286) );
  NOR2X0 U5539 ( .IN1(n3857), .IN2(n4602), .QN(WX8284) );
  NOR2X0 U5540 ( .IN1(n3858), .IN2(n4602), .QN(WX8282) );
  NOR2X0 U5541 ( .IN1(n3859), .IN2(n4602), .QN(WX8280) );
  NOR2X0 U5542 ( .IN1(n3860), .IN2(n4602), .QN(WX8278) );
  NOR2X0 U5543 ( .IN1(n3861), .IN2(n4602), .QN(WX8276) );
  NOR2X0 U5544 ( .IN1(n3862), .IN2(n4602), .QN(WX8274) );
  NOR2X0 U5545 ( .IN1(n3863), .IN2(n4602), .QN(WX8272) );
  NOR2X0 U5546 ( .IN1(n3864), .IN2(n4602), .QN(WX8270) );
  NOR2X0 U5547 ( .IN1(n3865), .IN2(n4602), .QN(WX8268) );
  NOR2X0 U5548 ( .IN1(n3866), .IN2(n4602), .QN(WX8266) );
  NOR2X0 U5549 ( .IN1(n3867), .IN2(n4602), .QN(WX8264) );
  NOR2X0 U5550 ( .IN1(n3868), .IN2(n4602), .QN(WX8262) );
  NOR2X0 U5551 ( .IN1(n3869), .IN2(n4602), .QN(WX8260) );
  NOR2X0 U5552 ( .IN1(n3870), .IN2(n4603), .QN(WX8258) );
  NOR2X0 U5553 ( .IN1(n3871), .IN2(n4603), .QN(WX8256) );
  NOR2X0 U5554 ( .IN1(n3872), .IN2(n4603), .QN(WX8254) );
  NOR2X0 U5555 ( .IN1(n3873), .IN2(n4603), .QN(WX8252) );
  NOR2X0 U5556 ( .IN1(n3874), .IN2(n4603), .QN(WX8250) );
  NOR2X0 U5557 ( .IN1(n3875), .IN2(n4603), .QN(WX8248) );
  NOR2X0 U5558 ( .IN1(n3876), .IN2(n4603), .QN(WX8246) );
  NOR2X0 U5559 ( .IN1(n3877), .IN2(n4603), .QN(WX8244) );
  NOR2X0 U5560 ( .IN1(n3878), .IN2(n4603), .QN(WX8242) );
  NOR2X0 U5561 ( .IN1(n3879), .IN2(n4633), .QN(WX7009) );
  NOR2X0 U5562 ( .IN1(n3880), .IN2(n4633), .QN(WX7007) );
  NOR2X0 U5563 ( .IN1(n3881), .IN2(n4633), .QN(WX7005) );
  NOR2X0 U5564 ( .IN1(n3882), .IN2(n4633), .QN(WX7003) );
  NOR2X0 U5565 ( .IN1(n3883), .IN2(n4633), .QN(WX7001) );
  NOR2X0 U5566 ( .IN1(n3884), .IN2(n4634), .QN(WX6999) );
  NOR2X0 U5567 ( .IN1(n3885), .IN2(n4634), .QN(WX6997) );
  NOR2X0 U5568 ( .IN1(n3886), .IN2(n4634), .QN(WX6995) );
  NOR2X0 U5569 ( .IN1(n3887), .IN2(n4634), .QN(WX6993) );
  NOR2X0 U5570 ( .IN1(n3888), .IN2(n4634), .QN(WX6991) );
  NOR2X0 U5571 ( .IN1(n3889), .IN2(n4634), .QN(WX6989) );
  NOR2X0 U5572 ( .IN1(n3890), .IN2(n4634), .QN(WX6987) );
  NOR2X0 U5573 ( .IN1(n3891), .IN2(n4634), .QN(WX6985) );
  NOR2X0 U5574 ( .IN1(n3892), .IN2(n4634), .QN(WX6983) );
  NOR2X0 U5575 ( .IN1(n3893), .IN2(n4634), .QN(WX6981) );
  NOR2X0 U5576 ( .IN1(n3894), .IN2(n4634), .QN(WX6979) );
  NOR2X0 U5577 ( .IN1(n3895), .IN2(n4634), .QN(WX6977) );
  NOR2X0 U5578 ( .IN1(n3896), .IN2(n4634), .QN(WX6975) );
  NOR2X0 U5579 ( .IN1(n3897), .IN2(n4634), .QN(WX6973) );
  NOR2X0 U5580 ( .IN1(n3898), .IN2(n4634), .QN(WX6971) );
  NOR2X0 U5581 ( .IN1(n3899), .IN2(n4635), .QN(WX6969) );
  NOR2X0 U5582 ( .IN1(n3900), .IN2(n4635), .QN(WX6967) );
  NOR2X0 U5583 ( .IN1(n3901), .IN2(n4635), .QN(WX6965) );
  NOR2X0 U5584 ( .IN1(n3902), .IN2(n4635), .QN(WX6963) );
  NOR2X0 U5585 ( .IN1(n3903), .IN2(n4635), .QN(WX6961) );
  NOR2X0 U5586 ( .IN1(n3904), .IN2(n4635), .QN(WX6959) );
  NOR2X0 U5587 ( .IN1(n3905), .IN2(n4635), .QN(WX6957) );
  NOR2X0 U5588 ( .IN1(n3906), .IN2(n4635), .QN(WX6955) );
  NOR2X0 U5589 ( .IN1(n3907), .IN2(n4635), .QN(WX6953) );
  NOR2X0 U5590 ( .IN1(n3908), .IN2(n4635), .QN(WX6951) );
  NOR2X0 U5591 ( .IN1(n3909), .IN2(n4635), .QN(WX6949) );
  NOR2X0 U5592 ( .IN1(n3910), .IN2(n4620), .QN(WX5716) );
  NOR2X0 U5593 ( .IN1(n3911), .IN2(n4620), .QN(WX5714) );
  NOR2X0 U5594 ( .IN1(n3912), .IN2(n4620), .QN(WX5712) );
  NOR2X0 U5595 ( .IN1(n3913), .IN2(n4620), .QN(WX5710) );
  NOR2X0 U5596 ( .IN1(n3914), .IN2(n4620), .QN(WX5708) );
  NOR2X0 U5597 ( .IN1(n3915), .IN2(n4620), .QN(WX5706) );
  NOR2X0 U5598 ( .IN1(n3916), .IN2(n4620), .QN(WX5704) );
  NOR2X0 U5599 ( .IN1(n3917), .IN2(n4620), .QN(WX5702) );
  NOR2X0 U5600 ( .IN1(n3918), .IN2(n4620), .QN(WX5700) );
  NOR2X0 U5601 ( .IN1(n3919), .IN2(n4620), .QN(WX5698) );
  NOR2X0 U5602 ( .IN1(n3920), .IN2(n4621), .QN(WX5696) );
  NOR2X0 U5603 ( .IN1(n3921), .IN2(n4621), .QN(WX5694) );
  NOR2X0 U5604 ( .IN1(n3922), .IN2(n4621), .QN(WX5692) );
  NOR2X0 U5605 ( .IN1(n3923), .IN2(n4621), .QN(WX5690) );
  NOR2X0 U5606 ( .IN1(n3924), .IN2(n4621), .QN(WX5688) );
  NOR2X0 U5607 ( .IN1(n3925), .IN2(n4621), .QN(WX5686) );
  NOR2X0 U5608 ( .IN1(n3926), .IN2(n4621), .QN(WX5684) );
  NOR2X0 U5609 ( .IN1(n3927), .IN2(n4621), .QN(WX5682) );
  NOR2X0 U5610 ( .IN1(n3928), .IN2(n4621), .QN(WX5680) );
  NOR2X0 U5611 ( .IN1(n3929), .IN2(n4621), .QN(WX5678) );
  NOR2X0 U5612 ( .IN1(n3930), .IN2(n4621), .QN(WX5676) );
  NOR2X0 U5613 ( .IN1(n3931), .IN2(n4621), .QN(WX5674) );
  NOR2X0 U5614 ( .IN1(n3932), .IN2(n4621), .QN(WX5672) );
  NOR2X0 U5615 ( .IN1(n3933), .IN2(n4621), .QN(WX5670) );
  NOR2X0 U5616 ( .IN1(n3934), .IN2(n4621), .QN(WX5668) );
  NOR2X0 U5617 ( .IN1(n3935), .IN2(n4622), .QN(WX5666) );
  NOR2X0 U5618 ( .IN1(n3936), .IN2(n4622), .QN(WX5664) );
  NOR2X0 U5619 ( .IN1(n3937), .IN2(n4622), .QN(WX5662) );
  NOR2X0 U5620 ( .IN1(n3938), .IN2(n4622), .QN(WX5660) );
  NOR2X0 U5621 ( .IN1(n3939), .IN2(n4622), .QN(WX5658) );
  NOR2X0 U5622 ( .IN1(n3940), .IN2(n4622), .QN(WX5656) );
  NOR2X0 U5623 ( .IN1(n3941), .IN2(n4573), .QN(WX4423) );
  NOR2X0 U5624 ( .IN1(n3942), .IN2(n4572), .QN(WX4421) );
  NOR2X0 U5625 ( .IN1(n3943), .IN2(n4572), .QN(WX4419) );
  NOR2X0 U5626 ( .IN1(n3944), .IN2(n4572), .QN(WX4417) );
  NOR2X0 U5627 ( .IN1(n3945), .IN2(n4572), .QN(WX4415) );
  NOR2X0 U5628 ( .IN1(n3946), .IN2(n4573), .QN(WX4413) );
  NOR2X0 U5629 ( .IN1(n3947), .IN2(n4572), .QN(WX4411) );
  NOR2X0 U5630 ( .IN1(n3948), .IN2(n4572), .QN(WX4409) );
  NOR2X0 U5631 ( .IN1(n3949), .IN2(n4572), .QN(WX4407) );
  NOR2X0 U5632 ( .IN1(n3950), .IN2(n4572), .QN(WX4405) );
  NOR2X0 U5633 ( .IN1(n3951), .IN2(n4571), .QN(WX4403) );
  NOR2X0 U5634 ( .IN1(n3952), .IN2(n4572), .QN(WX4401) );
  NOR2X0 U5635 ( .IN1(n3953), .IN2(n4569), .QN(WX4399) );
  NOR2X0 U5636 ( .IN1(n3954), .IN2(n4568), .QN(WX4397) );
  NOR2X0 U5637 ( .IN1(n3955), .IN2(n4572), .QN(WX4395) );
  NOR2X0 U5638 ( .IN1(n3956), .IN2(n4566), .QN(WX4393) );
  NOR2X0 U5639 ( .IN1(n3957), .IN2(n4571), .QN(WX4391) );
  NOR2X0 U5640 ( .IN1(n3958), .IN2(n4564), .QN(WX4389) );
  NOR2X0 U5641 ( .IN1(n3959), .IN2(n4570), .QN(WX4387) );
  NOR2X0 U5642 ( .IN1(n3960), .IN2(n4560), .QN(WX4385) );
  NOR2X0 U5643 ( .IN1(n3961), .IN2(n4559), .QN(WX4383) );
  NOR2X0 U5644 ( .IN1(n3962), .IN2(n4567), .QN(WX4381) );
  NOR2X0 U5645 ( .IN1(n3963), .IN2(n4571), .QN(WX4379) );
  NOR2X0 U5646 ( .IN1(n3964), .IN2(n4558), .QN(WX4377) );
  NOR2X0 U5647 ( .IN1(n3965), .IN2(n4574), .QN(WX4375) );
  NOR2X0 U5648 ( .IN1(n3966), .IN2(n4565), .QN(WX4373) );
  NOR2X0 U5649 ( .IN1(n3967), .IN2(n4563), .QN(WX4371) );
  NOR2X0 U5650 ( .IN1(n3968), .IN2(n4562), .QN(WX4369) );
  NOR2X0 U5651 ( .IN1(n3969), .IN2(n4561), .QN(WX4367) );
  NOR2X0 U5652 ( .IN1(n3970), .IN2(n4556), .QN(WX4365) );
  NOR2X0 U5653 ( .IN1(n3971), .IN2(n4557), .QN(WX4363) );
  NOR2X0 U5654 ( .IN1(n3972), .IN2(n4592), .QN(WX3130) );
  NOR2X0 U5655 ( .IN1(n3973), .IN2(n4588), .QN(WX3128) );
  NOR2X0 U5656 ( .IN1(n3974), .IN2(n4588), .QN(WX3126) );
  NOR2X0 U5657 ( .IN1(n3975), .IN2(n4588), .QN(WX3124) );
  NOR2X0 U5658 ( .IN1(n3976), .IN2(n4588), .QN(WX3122) );
  NOR2X0 U5659 ( .IN1(n3977), .IN2(n4588), .QN(WX3120) );
  NOR2X0 U5660 ( .IN1(n3978), .IN2(n4588), .QN(WX3118) );
  NOR2X0 U5661 ( .IN1(n3979), .IN2(n4588), .QN(WX3116) );
  NOR2X0 U5662 ( .IN1(n3980), .IN2(n4588), .QN(WX3114) );
  NOR2X0 U5663 ( .IN1(n3981), .IN2(n4588), .QN(WX3112) );
  NOR2X0 U5664 ( .IN1(n3982), .IN2(n4589), .QN(WX3110) );
  NOR2X0 U5665 ( .IN1(n3983), .IN2(n4589), .QN(WX3108) );
  NOR2X0 U5666 ( .IN1(n3984), .IN2(n4589), .QN(WX3106) );
  NOR2X0 U5667 ( .IN1(n3985), .IN2(n4589), .QN(WX3104) );
  NOR2X0 U5668 ( .IN1(n3986), .IN2(n4589), .QN(WX3102) );
  NOR2X0 U5669 ( .IN1(n3987), .IN2(n4589), .QN(WX3100) );
  NOR2X0 U5670 ( .IN1(n3988), .IN2(n4589), .QN(WX3098) );
  NOR2X0 U5671 ( .IN1(n3989), .IN2(n4589), .QN(WX3096) );
  NOR2X0 U5672 ( .IN1(n3990), .IN2(n4589), .QN(WX3094) );
  NOR2X0 U5673 ( .IN1(n3991), .IN2(n4589), .QN(WX3092) );
  NOR2X0 U5674 ( .IN1(n3992), .IN2(n4589), .QN(WX3090) );
  NOR2X0 U5675 ( .IN1(n3993), .IN2(n4589), .QN(WX3088) );
  NOR2X0 U5676 ( .IN1(n3994), .IN2(n4589), .QN(WX3086) );
  NOR2X0 U5677 ( .IN1(n3995), .IN2(n4589), .QN(WX3084) );
  NOR2X0 U5678 ( .IN1(n3996), .IN2(n4589), .QN(WX3082) );
  NOR2X0 U5679 ( .IN1(n3997), .IN2(n4590), .QN(WX3080) );
  NOR2X0 U5680 ( .IN1(n3998), .IN2(n4590), .QN(WX3078) );
  NOR2X0 U5681 ( .IN1(n3999), .IN2(n4590), .QN(WX3076) );
  NOR2X0 U5682 ( .IN1(n4000), .IN2(n4590), .QN(WX3074) );
  NOR2X0 U5683 ( .IN1(n4001), .IN2(n4590), .QN(WX3072) );
  NOR2X0 U5684 ( .IN1(n4002), .IN2(n4590), .QN(WX3070) );
  NOR2X0 U5685 ( .IN1(n4003), .IN2(n4595), .QN(WX1837) );
  NOR2X0 U5686 ( .IN1(n4004), .IN2(n4595), .QN(WX1835) );
  NOR2X0 U5687 ( .IN1(n4005), .IN2(n4595), .QN(WX1833) );
  NOR2X0 U5688 ( .IN1(n4006), .IN2(n4596), .QN(WX1831) );
  NOR2X0 U5689 ( .IN1(n4007), .IN2(n4596), .QN(WX1829) );
  NOR2X0 U5690 ( .IN1(n4008), .IN2(n4596), .QN(WX1827) );
  NOR2X0 U5691 ( .IN1(n4009), .IN2(n4596), .QN(WX1825) );
  NOR2X0 U5692 ( .IN1(n4010), .IN2(n4596), .QN(WX1823) );
  NOR2X0 U5693 ( .IN1(n4011), .IN2(n4596), .QN(WX1821) );
  NOR2X0 U5694 ( .IN1(n4012), .IN2(n4596), .QN(WX1819) );
  NOR2X0 U5695 ( .IN1(n4013), .IN2(n4596), .QN(WX1817) );
  NOR2X0 U5696 ( .IN1(n4014), .IN2(n4596), .QN(WX1815) );
  NOR2X0 U5697 ( .IN1(n4015), .IN2(n4596), .QN(WX1813) );
  NOR2X0 U5698 ( .IN1(n4016), .IN2(n4596), .QN(WX1811) );
  NOR2X0 U5699 ( .IN1(n4017), .IN2(n4596), .QN(WX1809) );
  NOR2X0 U5700 ( .IN1(n4018), .IN2(n4596), .QN(WX1807) );
  NOR2X0 U5701 ( .IN1(n4019), .IN2(n4584), .QN(WX1805) );
  NOR2X0 U5702 ( .IN1(n4020), .IN2(n4579), .QN(WX1803) );
  NOR2X0 U5703 ( .IN1(n4021), .IN2(n4580), .QN(WX1801) );
  NOR2X0 U5704 ( .IN1(n4022), .IN2(n4580), .QN(WX1799) );
  NOR2X0 U5705 ( .IN1(n4023), .IN2(n4580), .QN(WX1797) );
  NOR2X0 U5706 ( .IN1(n4024), .IN2(n4580), .QN(WX1795) );
  NOR2X0 U5707 ( .IN1(n4025), .IN2(n4580), .QN(WX1793) );
  NOR2X0 U5708 ( .IN1(n4026), .IN2(n4580), .QN(WX1791) );
  NOR2X0 U5709 ( .IN1(n4027), .IN2(n4580), .QN(WX1789) );
  NOR2X0 U5710 ( .IN1(n4028), .IN2(n4580), .QN(WX1787) );
  NOR2X0 U5711 ( .IN1(n4029), .IN2(n4580), .QN(WX1785) );
  NOR2X0 U5712 ( .IN1(n4030), .IN2(n4580), .QN(WX1783) );
  NOR2X0 U5713 ( .IN1(n4031), .IN2(n4580), .QN(WX1781) );
  NOR2X0 U5714 ( .IN1(n4032), .IN2(n4580), .QN(WX1779) );
  NOR2X0 U5715 ( .IN1(n4033), .IN2(n4580), .QN(WX1777) );
  ISOLANDX1 U5716 ( .D(WX547), .ISO(n4622), .Q(WX544) );
  ISOLANDX1 U5717 ( .D(WX545), .ISO(n4622), .Q(WX542) );
  ISOLANDX1 U5718 ( .D(WX543), .ISO(n4622), .Q(WX540) );
  ISOLANDX1 U5719 ( .D(WX541), .ISO(n4622), .Q(WX538) );
  ISOLANDX1 U5720 ( .D(WX539), .ISO(n4622), .Q(WX536) );
  ISOLANDX1 U5721 ( .D(WX537), .ISO(n4622), .Q(WX534) );
  ISOLANDX1 U5722 ( .D(WX535), .ISO(n4622), .Q(WX532) );
  ISOLANDX1 U5723 ( .D(WX533), .ISO(n4622), .Q(WX530) );
  ISOLANDX1 U5724 ( .D(WX531), .ISO(n4623), .Q(WX528) );
  ISOLANDX1 U5725 ( .D(WX529), .ISO(n4623), .Q(WX526) );
  ISOLANDX1 U5726 ( .D(WX527), .ISO(n4623), .Q(WX524) );
  ISOLANDX1 U5727 ( .D(WX525), .ISO(n4623), .Q(WX522) );
  ISOLANDX1 U5728 ( .D(WX523), .ISO(n4623), .Q(WX520) );
  ISOLANDX1 U5729 ( .D(WX521), .ISO(n4623), .Q(WX518) );
  ISOLANDX1 U5730 ( .D(test_so1), .ISO(n4623), .Q(WX516) );
  ISOLANDX1 U5731 ( .D(WX517), .ISO(n4623), .Q(WX514) );
  ISOLANDX1 U5732 ( .D(WX515), .ISO(n4623), .Q(WX512) );
  ISOLANDX1 U5733 ( .D(WX513), .ISO(n4623), .Q(WX510) );
  ISOLANDX1 U5734 ( .D(WX511), .ISO(n4623), .Q(WX508) );
  ISOLANDX1 U5735 ( .D(WX509), .ISO(n4623), .Q(WX506) );
  ISOLANDX1 U5736 ( .D(WX507), .ISO(n4623), .Q(WX504) );
  ISOLANDX1 U5737 ( .D(WX505), .ISO(n4623), .Q(WX502) );
  ISOLANDX1 U5738 ( .D(WX503), .ISO(n4623), .Q(WX500) );
  ISOLANDX1 U5739 ( .D(WX501), .ISO(n4624), .Q(WX498) );
  ISOLANDX1 U5740 ( .D(WX499), .ISO(n4624), .Q(WX496) );
  ISOLANDX1 U5741 ( .D(WX497), .ISO(n4624), .Q(WX494) );
  ISOLANDX1 U5742 ( .D(WX495), .ISO(n4624), .Q(WX492) );
  ISOLANDX1 U5743 ( .D(WX493), .ISO(n4624), .Q(WX490) );
  ISOLANDX1 U5744 ( .D(WX491), .ISO(n4624), .Q(WX488) );
  ISOLANDX1 U5745 ( .D(WX489), .ISO(n4624), .Q(WX486) );
  ISOLANDX1 U5746 ( .D(WX487), .ISO(n4624), .Q(WX484) );
  ISOLANDX1 U5747 ( .D(WX5939), .ISO(n4638), .Q(WX6002) );
  ISOLANDX1 U5748 ( .D(test_so49), .ISO(n4638), .Q(WX6000) );
  ISOLANDX1 U5749 ( .D(WX5935), .ISO(n4638), .Q(WX5998) );
  ISOLANDX1 U5750 ( .D(WX5933), .ISO(n4638), .Q(WX5996) );
  ISOLANDX1 U5751 ( .D(WX5931), .ISO(n4638), .Q(WX5994) );
  ISOLANDX1 U5752 ( .D(WX3269), .ISO(n4571), .Q(WX3332) );
  ISOLANDX1 U5753 ( .D(WX3265), .ISO(n4571), .Q(WX3328) );
  ISOLANDX1 U5754 ( .D(WX3263), .ISO(n4571), .Q(WX3326) );
  ISOLANDX1 U5755 ( .D(WX11179), .ISO(n4580), .Q(WX11242) );
  ISOLANDX1 U5756 ( .D(WX11177), .ISO(n4580), .Q(WX11240) );
  ISOLANDX1 U5757 ( .D(WX11175), .ISO(n4581), .Q(WX11238) );
  ISOLANDX1 U5758 ( .D(WX11173), .ISO(n4581), .Q(WX11236) );
  ISOLANDX1 U5759 ( .D(test_so96), .ISO(n4581), .Q(WX11234) );
  ISOLANDX1 U5760 ( .D(WX11169), .ISO(n4581), .Q(WX11232) );
  ISOLANDX1 U5761 ( .D(WX11167), .ISO(n4581), .Q(WX11230) );
  ISOLANDX1 U5762 ( .D(WX11165), .ISO(n4581), .Q(WX11228) );
  ISOLANDX1 U5763 ( .D(WX11163), .ISO(n4581), .Q(WX11226) );
  ISOLANDX1 U5764 ( .D(WX11161), .ISO(n4581), .Q(WX11224) );
  ISOLANDX1 U5765 ( .D(WX11159), .ISO(n4581), .Q(WX11222) );
  ISOLANDX1 U5766 ( .D(WX11157), .ISO(n4581), .Q(WX11220) );
  ISOLANDX1 U5767 ( .D(WX11155), .ISO(n4581), .Q(WX11218) );
  ISOLANDX1 U5768 ( .D(WX11153), .ISO(n4581), .Q(WX11216) );
  ISOLANDX1 U5769 ( .D(WX11151), .ISO(n4581), .Q(WX11214) );
  ISOLANDX1 U5770 ( .D(WX11149), .ISO(n4581), .Q(WX11212) );
  ISOLANDX1 U5771 ( .D(WX11147), .ISO(n4581), .Q(WX11210) );
  ISOLANDX1 U5772 ( .D(WX11145), .ISO(n4582), .Q(WX11208) );
  ISOLANDX1 U5773 ( .D(WX11143), .ISO(n4582), .Q(WX11206) );
  ISOLANDX1 U5774 ( .D(WX11141), .ISO(n4582), .Q(WX11204) );
  ISOLANDX1 U5775 ( .D(WX11139), .ISO(n4582), .Q(WX11202) );
  ISOLANDX1 U5776 ( .D(test_so95), .ISO(n4582), .Q(WX11200) );
  ISOLANDX1 U5777 ( .D(WX11135), .ISO(n4582), .Q(WX11198) );
  ISOLANDX1 U5778 ( .D(WX11133), .ISO(n4582), .Q(WX11196) );
  ISOLANDX1 U5779 ( .D(WX11131), .ISO(n4582), .Q(WX11194) );
  ISOLANDX1 U5780 ( .D(WX11129), .ISO(n4582), .Q(WX11192) );
  ISOLANDX1 U5781 ( .D(WX11127), .ISO(n4582), .Q(WX11190) );
  ISOLANDX1 U5782 ( .D(WX11125), .ISO(n4582), .Q(WX11188) );
  ISOLANDX1 U5783 ( .D(WX11123), .ISO(n4582), .Q(WX11186) );
  ISOLANDX1 U5784 ( .D(WX11121), .ISO(n4582), .Q(WX11184) );
  ISOLANDX1 U5785 ( .D(WX11119), .ISO(n4582), .Q(WX11182) );
  ISOLANDX1 U5786 ( .D(WX11117), .ISO(n4582), .Q(WX11180) );
  ISOLANDX1 U5787 ( .D(WX11115), .ISO(n4583), .Q(WX11178) );
  ISOLANDX1 U5788 ( .D(WX11113), .ISO(n4583), .Q(WX11176) );
  ISOLANDX1 U5789 ( .D(WX11111), .ISO(n4583), .Q(WX11174) );
  ISOLANDX1 U5790 ( .D(WX11109), .ISO(n4583), .Q(WX11172) );
  ISOLANDX1 U5791 ( .D(WX11107), .ISO(n4583), .Q(WX11170) );
  ISOLANDX1 U5792 ( .D(WX11105), .ISO(n4583), .Q(WX11168) );
  ISOLANDX1 U5793 ( .D(test_so94), .ISO(n4583), .Q(WX11166) );
  ISOLANDX1 U5794 ( .D(WX11101), .ISO(n4583), .Q(WX11164) );
  ISOLANDX1 U5795 ( .D(WX11099), .ISO(n4583), .Q(WX11162) );
  ISOLANDX1 U5796 ( .D(WX11097), .ISO(n4583), .Q(WX11160) );
  ISOLANDX1 U5797 ( .D(WX11095), .ISO(n4583), .Q(WX11158) );
  ISOLANDX1 U5798 ( .D(WX11093), .ISO(n4583), .Q(WX11156) );
  ISOLANDX1 U5799 ( .D(WX11091), .ISO(n4583), .Q(WX11154) );
  ISOLANDX1 U5800 ( .D(WX11089), .ISO(n4583), .Q(WX11152) );
  ISOLANDX1 U5801 ( .D(WX11087), .ISO(n4583), .Q(WX11150) );
  ISOLANDX1 U5802 ( .D(WX11085), .ISO(n4584), .Q(WX11148) );
  ISOLANDX1 U5803 ( .D(WX11083), .ISO(n4584), .Q(WX11146) );
  ISOLANDX1 U5804 ( .D(WX11081), .ISO(n4584), .Q(WX11144) );
  ISOLANDX1 U5805 ( .D(WX11079), .ISO(n4584), .Q(WX11142) );
  ISOLANDX1 U5806 ( .D(WX11077), .ISO(n4584), .Q(WX11140) );
  ISOLANDX1 U5807 ( .D(WX11075), .ISO(n4584), .Q(WX11138) );
  ISOLANDX1 U5808 ( .D(WX11073), .ISO(n4584), .Q(WX11136) );
  ISOLANDX1 U5809 ( .D(WX11071), .ISO(n4584), .Q(WX11134) );
  ISOLANDX1 U5810 ( .D(test_so93), .ISO(n4584), .Q(WX11132) );
  ISOLANDX1 U5811 ( .D(WX11067), .ISO(n4584), .Q(WX11130) );
  ISOLANDX1 U5812 ( .D(WX11065), .ISO(n4584), .Q(WX11128) );
  ISOLANDX1 U5813 ( .D(WX11063), .ISO(n4584), .Q(WX11126) );
  ISOLANDX1 U5814 ( .D(WX11061), .ISO(n4584), .Q(WX11124) );
  ISOLANDX1 U5815 ( .D(WX11059), .ISO(n4584), .Q(WX11122) );
  ISOLANDX1 U5816 ( .D(WX11057), .ISO(n4585), .Q(WX11120) );
  ISOLANDX1 U5817 ( .D(WX11055), .ISO(n4585), .Q(WX11118) );
  ISOLANDX1 U5818 ( .D(WX11053), .ISO(n4585), .Q(WX11116) );
  ISOLANDX1 U5819 ( .D(WX11051), .ISO(n4585), .Q(WX11114) );
  ISOLANDX1 U5820 ( .D(WX11049), .ISO(n4585), .Q(WX11112) );
  ISOLANDX1 U5821 ( .D(WX11047), .ISO(n4585), .Q(WX11110) );
  ISOLANDX1 U5822 ( .D(WX11045), .ISO(n4585), .Q(WX11108) );
  ISOLANDX1 U5823 ( .D(WX11043), .ISO(n4585), .Q(WX11106) );
  ISOLANDX1 U5824 ( .D(WX11041), .ISO(n4585), .Q(WX11104) );
  ISOLANDX1 U5825 ( .D(WX11039), .ISO(n4585), .Q(WX11102) );
  ISOLANDX1 U5826 ( .D(WX11037), .ISO(n4585), .Q(WX11100) );
  ISOLANDX1 U5827 ( .D(test_so92), .ISO(n4585), .Q(WX11098) );
  ISOLANDX1 U5828 ( .D(WX11033), .ISO(n4585), .Q(WX11096) );
  ISOLANDX1 U5829 ( .D(WX11031), .ISO(n4585), .Q(WX11094) );
  ISOLANDX1 U5830 ( .D(WX11029), .ISO(n4585), .Q(WX11092) );
  ISOLANDX1 U5831 ( .D(WX11027), .ISO(n4586), .Q(WX11090) );
  ISOLANDX1 U5832 ( .D(WX11025), .ISO(n4586), .Q(WX11088) );
  ISOLANDX1 U5833 ( .D(WX11023), .ISO(n4586), .Q(WX11086) );
  ISOLANDX1 U5834 ( .D(WX11021), .ISO(n4586), .Q(WX11084) );
  ISOLANDX1 U5835 ( .D(WX9886), .ISO(n4596), .Q(WX9949) );
  ISOLANDX1 U5836 ( .D(WX9884), .ISO(n4572), .Q(WX9947) );
  ISOLANDX1 U5837 ( .D(WX9882), .ISO(n4617), .Q(WX9945) );
  ISOLANDX1 U5838 ( .D(WX9880), .ISO(n4612), .Q(WX9943) );
  ISOLANDX1 U5839 ( .D(WX9878), .ISO(n4607), .Q(WX9941) );
  ISOLANDX1 U5840 ( .D(WX9876), .ISO(n4607), .Q(WX9939) );
  ISOLANDX1 U5841 ( .D(WX9874), .ISO(n4607), .Q(WX9937) );
  ISOLANDX1 U5842 ( .D(WX9872), .ISO(n4607), .Q(WX9935) );
  ISOLANDX1 U5843 ( .D(WX9870), .ISO(n4607), .Q(WX9933) );
  ISOLANDX1 U5844 ( .D(WX9868), .ISO(n4607), .Q(WX9931) );
  ISOLANDX1 U5845 ( .D(WX9866), .ISO(n4607), .Q(WX9929) );
  ISOLANDX1 U5846 ( .D(WX9864), .ISO(n4607), .Q(WX9927) );
  ISOLANDX1 U5847 ( .D(WX9862), .ISO(n4607), .Q(WX9925) );
  ISOLANDX1 U5848 ( .D(WX9860), .ISO(n4607), .Q(WX9923) );
  ISOLANDX1 U5849 ( .D(WX9858), .ISO(n4607), .Q(WX9921) );
  ISOLANDX1 U5850 ( .D(WX9856), .ISO(n4608), .Q(WX9919) );
  ISOLANDX1 U5851 ( .D(test_so84), .ISO(n4608), .Q(WX9917) );
  ISOLANDX1 U5852 ( .D(WX9852), .ISO(n4608), .Q(WX9915) );
  ISOLANDX1 U5853 ( .D(WX9850), .ISO(n4608), .Q(WX9913) );
  ISOLANDX1 U5854 ( .D(WX9848), .ISO(n4608), .Q(WX9911) );
  ISOLANDX1 U5855 ( .D(WX9846), .ISO(n4608), .Q(WX9909) );
  ISOLANDX1 U5856 ( .D(WX9844), .ISO(n4608), .Q(WX9907) );
  ISOLANDX1 U5857 ( .D(WX9842), .ISO(n4608), .Q(WX9905) );
  ISOLANDX1 U5858 ( .D(WX9840), .ISO(n4608), .Q(WX9903) );
  ISOLANDX1 U5859 ( .D(WX9838), .ISO(n4608), .Q(WX9901) );
  ISOLANDX1 U5860 ( .D(WX9836), .ISO(n4608), .Q(WX9899) );
  ISOLANDX1 U5861 ( .D(WX9834), .ISO(n4608), .Q(WX9897) );
  ISOLANDX1 U5862 ( .D(WX9832), .ISO(n4608), .Q(WX9895) );
  ISOLANDX1 U5863 ( .D(WX9830), .ISO(n4608), .Q(WX9893) );
  ISOLANDX1 U5864 ( .D(WX9828), .ISO(n4608), .Q(WX9891) );
  ISOLANDX1 U5865 ( .D(WX9826), .ISO(n4609), .Q(WX9889) );
  ISOLANDX1 U5866 ( .D(WX9824), .ISO(n4609), .Q(WX9887) );
  ISOLANDX1 U5867 ( .D(WX9822), .ISO(n4609), .Q(WX9885) );
  ISOLANDX1 U5868 ( .D(test_so83), .ISO(n4609), .Q(WX9883) );
  ISOLANDX1 U5869 ( .D(WX9818), .ISO(n4609), .Q(WX9881) );
  ISOLANDX1 U5870 ( .D(WX9816), .ISO(n4609), .Q(WX9879) );
  ISOLANDX1 U5871 ( .D(WX9814), .ISO(n4609), .Q(WX9877) );
  ISOLANDX1 U5872 ( .D(WX9812), .ISO(n4609), .Q(WX9875) );
  ISOLANDX1 U5873 ( .D(WX9810), .ISO(n4609), .Q(WX9873) );
  ISOLANDX1 U5874 ( .D(WX9808), .ISO(n4609), .Q(WX9871) );
  ISOLANDX1 U5875 ( .D(WX9806), .ISO(n4609), .Q(WX9869) );
  ISOLANDX1 U5876 ( .D(WX9804), .ISO(n4609), .Q(WX9867) );
  ISOLANDX1 U5877 ( .D(WX9802), .ISO(n4609), .Q(WX9865) );
  ISOLANDX1 U5878 ( .D(WX9800), .ISO(n4609), .Q(WX9863) );
  ISOLANDX1 U5879 ( .D(WX9798), .ISO(n4609), .Q(WX9861) );
  ISOLANDX1 U5880 ( .D(WX9796), .ISO(n4610), .Q(WX9859) );
  ISOLANDX1 U5881 ( .D(WX9794), .ISO(n4610), .Q(WX9857) );
  ISOLANDX1 U5882 ( .D(WX9792), .ISO(n4610), .Q(WX9855) );
  ISOLANDX1 U5883 ( .D(WX9790), .ISO(n4610), .Q(WX9853) );
  ISOLANDX1 U5884 ( .D(WX9788), .ISO(n4610), .Q(WX9851) );
  ISOLANDX1 U5885 ( .D(test_so82), .ISO(n4610), .Q(WX9849) );
  ISOLANDX1 U5886 ( .D(WX9784), .ISO(n4610), .Q(WX9847) );
  ISOLANDX1 U5887 ( .D(WX9782), .ISO(n4610), .Q(WX9845) );
  ISOLANDX1 U5888 ( .D(WX9780), .ISO(n4610), .Q(WX9843) );
  ISOLANDX1 U5889 ( .D(WX9778), .ISO(n4610), .Q(WX9841) );
  ISOLANDX1 U5890 ( .D(WX9776), .ISO(n4610), .Q(WX9839) );
  ISOLANDX1 U5891 ( .D(WX9774), .ISO(n4610), .Q(WX9837) );
  ISOLANDX1 U5892 ( .D(WX9772), .ISO(n4610), .Q(WX9835) );
  ISOLANDX1 U5893 ( .D(WX9770), .ISO(n4610), .Q(WX9833) );
  ISOLANDX1 U5894 ( .D(WX9768), .ISO(n4610), .Q(WX9831) );
  ISOLANDX1 U5895 ( .D(WX9766), .ISO(n4611), .Q(WX9829) );
  ISOLANDX1 U5896 ( .D(WX9764), .ISO(n4611), .Q(WX9827) );
  ISOLANDX1 U5897 ( .D(WX9762), .ISO(n4611), .Q(WX9825) );
  ISOLANDX1 U5898 ( .D(WX9760), .ISO(n4611), .Q(WX9823) );
  ISOLANDX1 U5899 ( .D(WX9758), .ISO(n4611), .Q(WX9821) );
  ISOLANDX1 U5900 ( .D(WX9756), .ISO(n4611), .Q(WX9819) );
  ISOLANDX1 U5901 ( .D(WX9754), .ISO(n4611), .Q(WX9817) );
  ISOLANDX1 U5902 ( .D(test_so81), .ISO(n4611), .Q(WX9815) );
  ISOLANDX1 U5903 ( .D(WX9750), .ISO(n4611), .Q(WX9813) );
  ISOLANDX1 U5904 ( .D(WX9748), .ISO(n4611), .Q(WX9811) );
  ISOLANDX1 U5905 ( .D(WX9746), .ISO(n4611), .Q(WX9809) );
  ISOLANDX1 U5906 ( .D(WX9744), .ISO(n4611), .Q(WX9807) );
  ISOLANDX1 U5907 ( .D(WX9742), .ISO(n4611), .Q(WX9805) );
  ISOLANDX1 U5908 ( .D(WX9740), .ISO(n4611), .Q(WX9803) );
  ISOLANDX1 U5909 ( .D(WX9738), .ISO(n4611), .Q(WX9801) );
  ISOLANDX1 U5910 ( .D(WX9736), .ISO(n4612), .Q(WX9799) );
  ISOLANDX1 U5911 ( .D(WX9734), .ISO(n4612), .Q(WX9797) );
  ISOLANDX1 U5912 ( .D(WX9732), .ISO(n4612), .Q(WX9795) );
  ISOLANDX1 U5913 ( .D(WX9730), .ISO(n4612), .Q(WX9793) );
  ISOLANDX1 U5914 ( .D(WX9728), .ISO(n4612), .Q(WX9791) );
  ISOLANDX1 U5915 ( .D(WX8593), .ISO(n4615), .Q(WX8656) );
  ISOLANDX1 U5916 ( .D(WX8591), .ISO(n4615), .Q(WX8654) );
  ISOLANDX1 U5917 ( .D(WX8589), .ISO(n4615), .Q(WX8652) );
  ISOLANDX1 U5918 ( .D(WX8587), .ISO(n4615), .Q(WX8650) );
  ISOLANDX1 U5919 ( .D(WX8585), .ISO(n4615), .Q(WX8648) );
  ISOLANDX1 U5920 ( .D(WX8583), .ISO(n4615), .Q(WX8646) );
  ISOLANDX1 U5921 ( .D(WX8581), .ISO(n4616), .Q(WX8644) );
  ISOLANDX1 U5922 ( .D(WX8579), .ISO(n4616), .Q(WX8642) );
  ISOLANDX1 U5923 ( .D(WX8577), .ISO(n4616), .Q(WX8640) );
  ISOLANDX1 U5924 ( .D(WX8575), .ISO(n4616), .Q(WX8638) );
  ISOLANDX1 U5925 ( .D(WX8573), .ISO(n4616), .Q(WX8636) );
  ISOLANDX1 U5926 ( .D(test_so73), .ISO(n4616), .Q(WX8634) );
  ISOLANDX1 U5927 ( .D(WX8569), .ISO(n4616), .Q(WX8632) );
  ISOLANDX1 U5928 ( .D(WX8567), .ISO(n4616), .Q(WX8630) );
  ISOLANDX1 U5929 ( .D(WX8565), .ISO(n4616), .Q(WX8628) );
  ISOLANDX1 U5930 ( .D(WX8563), .ISO(n4616), .Q(WX8626) );
  ISOLANDX1 U5931 ( .D(WX8561), .ISO(n4616), .Q(WX8624) );
  ISOLANDX1 U5932 ( .D(WX8559), .ISO(n4616), .Q(WX8622) );
  ISOLANDX1 U5933 ( .D(WX8557), .ISO(n4616), .Q(WX8620) );
  ISOLANDX1 U5934 ( .D(WX8555), .ISO(n4617), .Q(WX8618) );
  ISOLANDX1 U5935 ( .D(WX8553), .ISO(n4617), .Q(WX8616) );
  ISOLANDX1 U5936 ( .D(WX8551), .ISO(n4617), .Q(WX8614) );
  ISOLANDX1 U5937 ( .D(WX8549), .ISO(n4617), .Q(WX8612) );
  ISOLANDX1 U5938 ( .D(WX8547), .ISO(n4617), .Q(WX8610) );
  ISOLANDX1 U5939 ( .D(WX8545), .ISO(n4617), .Q(WX8608) );
  ISOLANDX1 U5940 ( .D(WX8543), .ISO(n4617), .Q(WX8606) );
  ISOLANDX1 U5941 ( .D(WX8541), .ISO(n4617), .Q(WX8604) );
  ISOLANDX1 U5942 ( .D(WX8539), .ISO(n4617), .Q(WX8602) );
  ISOLANDX1 U5943 ( .D(test_so72), .ISO(n4602), .Q(WX8600) );
  ISOLANDX1 U5944 ( .D(WX8535), .ISO(n4597), .Q(WX8598) );
  ISOLANDX1 U5945 ( .D(WX8533), .ISO(n4597), .Q(WX8596) );
  ISOLANDX1 U5946 ( .D(WX8531), .ISO(n4597), .Q(WX8594) );
  ISOLANDX1 U5947 ( .D(WX8529), .ISO(n4597), .Q(WX8592) );
  ISOLANDX1 U5948 ( .D(WX8527), .ISO(n4597), .Q(WX8590) );
  ISOLANDX1 U5949 ( .D(WX8525), .ISO(n4597), .Q(WX8588) );
  ISOLANDX1 U5950 ( .D(WX8523), .ISO(n4597), .Q(WX8586) );
  ISOLANDX1 U5951 ( .D(WX8521), .ISO(n4597), .Q(WX8584) );
  ISOLANDX1 U5952 ( .D(WX8519), .ISO(n4597), .Q(WX8582) );
  ISOLANDX1 U5953 ( .D(WX8517), .ISO(n4597), .Q(WX8580) );
  ISOLANDX1 U5954 ( .D(WX8515), .ISO(n4597), .Q(WX8578) );
  ISOLANDX1 U5955 ( .D(WX8513), .ISO(n4597), .Q(WX8576) );
  ISOLANDX1 U5956 ( .D(WX8511), .ISO(n4597), .Q(WX8574) );
  ISOLANDX1 U5957 ( .D(WX8509), .ISO(n4597), .Q(WX8572) );
  ISOLANDX1 U5958 ( .D(WX8507), .ISO(n4598), .Q(WX8570) );
  ISOLANDX1 U5959 ( .D(WX8505), .ISO(n4598), .Q(WX8568) );
  ISOLANDX1 U5960 ( .D(test_so71), .ISO(n4598), .Q(WX8566) );
  ISOLANDX1 U5961 ( .D(WX8501), .ISO(n4598), .Q(WX8564) );
  ISOLANDX1 U5962 ( .D(WX8499), .ISO(n4598), .Q(WX8562) );
  ISOLANDX1 U5963 ( .D(WX8497), .ISO(n4598), .Q(WX8560) );
  ISOLANDX1 U5964 ( .D(WX8495), .ISO(n4598), .Q(WX8558) );
  ISOLANDX1 U5965 ( .D(WX8493), .ISO(n4598), .Q(WX8556) );
  ISOLANDX1 U5966 ( .D(WX8491), .ISO(n4598), .Q(WX8554) );
  ISOLANDX1 U5967 ( .D(WX8489), .ISO(n4598), .Q(WX8552) );
  ISOLANDX1 U5968 ( .D(WX8487), .ISO(n4598), .Q(WX8550) );
  ISOLANDX1 U5969 ( .D(WX8485), .ISO(n4598), .Q(WX8548) );
  ISOLANDX1 U5970 ( .D(WX8483), .ISO(n4598), .Q(WX8546) );
  ISOLANDX1 U5971 ( .D(WX8481), .ISO(n4598), .Q(WX8544) );
  ISOLANDX1 U5972 ( .D(WX8479), .ISO(n4599), .Q(WX8542) );
  ISOLANDX1 U5973 ( .D(WX8477), .ISO(n4599), .Q(WX8540) );
  ISOLANDX1 U5974 ( .D(WX8475), .ISO(n4599), .Q(WX8538) );
  ISOLANDX1 U5975 ( .D(WX8473), .ISO(n4599), .Q(WX8536) );
  ISOLANDX1 U5976 ( .D(WX8471), .ISO(n4599), .Q(WX8534) );
  ISOLANDX1 U5977 ( .D(test_so70), .ISO(n4599), .Q(WX8532) );
  ISOLANDX1 U5978 ( .D(WX8467), .ISO(n4599), .Q(WX8530) );
  ISOLANDX1 U5979 ( .D(WX8465), .ISO(n4599), .Q(WX8528) );
  ISOLANDX1 U5980 ( .D(WX8463), .ISO(n4599), .Q(WX8526) );
  ISOLANDX1 U5981 ( .D(WX8461), .ISO(n4599), .Q(WX8524) );
  ISOLANDX1 U5982 ( .D(WX8459), .ISO(n4599), .Q(WX8522) );
  ISOLANDX1 U5983 ( .D(WX8457), .ISO(n4599), .Q(WX8520) );
  ISOLANDX1 U5984 ( .D(WX8455), .ISO(n4599), .Q(WX8518) );
  ISOLANDX1 U5985 ( .D(WX8453), .ISO(n4600), .Q(WX8516) );
  ISOLANDX1 U5986 ( .D(WX8451), .ISO(n4600), .Q(WX8514) );
  ISOLANDX1 U5987 ( .D(WX8449), .ISO(n4600), .Q(WX8512) );
  ISOLANDX1 U5988 ( .D(WX8447), .ISO(n4600), .Q(WX8510) );
  ISOLANDX1 U5989 ( .D(WX8445), .ISO(n4600), .Q(WX8508) );
  ISOLANDX1 U5990 ( .D(WX8443), .ISO(n4600), .Q(WX8506) );
  ISOLANDX1 U5991 ( .D(WX8441), .ISO(n4600), .Q(WX8504) );
  ISOLANDX1 U5992 ( .D(WX8439), .ISO(n4600), .Q(WX8502) );
  ISOLANDX1 U5993 ( .D(WX8437), .ISO(n4600), .Q(WX8500) );
  ISOLANDX1 U5994 ( .D(test_so69), .ISO(n4600), .Q(WX8498) );
  ISOLANDX1 U5995 ( .D(WX7300), .ISO(n4606), .Q(WX7363) );
  ISOLANDX1 U5996 ( .D(WX7298), .ISO(n4606), .Q(WX7361) );
  ISOLANDX1 U5997 ( .D(WX7296), .ISO(n4606), .Q(WX7359) );
  ISOLANDX1 U5998 ( .D(WX7294), .ISO(n4606), .Q(WX7357) );
  ISOLANDX1 U5999 ( .D(WX7292), .ISO(n4606), .Q(WX7355) );
  ISOLANDX1 U6000 ( .D(WX7290), .ISO(n4607), .Q(WX7353) );
  ISOLANDX1 U6001 ( .D(test_so62), .ISO(n4607), .Q(WX7351) );
  ISOLANDX1 U6002 ( .D(WX7286), .ISO(n4607), .Q(WX7349) );
  ISOLANDX1 U6003 ( .D(WX7284), .ISO(n4607), .Q(WX7347) );
  ISOLANDX1 U6004 ( .D(WX7282), .ISO(n4633), .Q(WX7345) );
  ISOLANDX1 U6005 ( .D(WX7280), .ISO(n4628), .Q(WX7343) );
  ISOLANDX1 U6006 ( .D(WX7278), .ISO(n4628), .Q(WX7341) );
  ISOLANDX1 U6007 ( .D(WX7276), .ISO(n4628), .Q(WX7339) );
  ISOLANDX1 U6008 ( .D(WX7274), .ISO(n4628), .Q(WX7337) );
  ISOLANDX1 U6009 ( .D(WX7272), .ISO(n4628), .Q(WX7335) );
  ISOLANDX1 U6010 ( .D(WX7270), .ISO(n4628), .Q(WX7333) );
  ISOLANDX1 U6011 ( .D(WX7268), .ISO(n4628), .Q(WX7331) );
  ISOLANDX1 U6012 ( .D(WX7266), .ISO(n4628), .Q(WX7329) );
  ISOLANDX1 U6013 ( .D(WX7264), .ISO(n4628), .Q(WX7327) );
  ISOLANDX1 U6014 ( .D(WX7262), .ISO(n4628), .Q(WX7325) );
  ISOLANDX1 U6015 ( .D(WX7260), .ISO(n4628), .Q(WX7323) );
  ISOLANDX1 U6016 ( .D(WX7258), .ISO(n4628), .Q(WX7321) );
  ISOLANDX1 U6017 ( .D(WX7256), .ISO(n4628), .Q(WX7319) );
  ISOLANDX1 U6018 ( .D(test_so61), .ISO(n4629), .Q(WX7317) );
  ISOLANDX1 U6019 ( .D(WX7252), .ISO(n4629), .Q(WX7315) );
  ISOLANDX1 U6020 ( .D(WX7250), .ISO(n4629), .Q(WX7313) );
  ISOLANDX1 U6021 ( .D(WX7248), .ISO(n4629), .Q(WX7311) );
  ISOLANDX1 U6022 ( .D(WX7246), .ISO(n4629), .Q(WX7309) );
  ISOLANDX1 U6023 ( .D(WX7244), .ISO(n4629), .Q(WX7307) );
  ISOLANDX1 U6024 ( .D(WX7242), .ISO(n4629), .Q(WX7305) );
  ISOLANDX1 U6025 ( .D(WX7240), .ISO(n4629), .Q(WX7303) );
  ISOLANDX1 U6026 ( .D(WX7238), .ISO(n4629), .Q(WX7301) );
  ISOLANDX1 U6027 ( .D(WX7236), .ISO(n4629), .Q(WX7299) );
  ISOLANDX1 U6028 ( .D(WX7234), .ISO(n4629), .Q(WX7297) );
  ISOLANDX1 U6029 ( .D(WX7232), .ISO(n4629), .Q(WX7295) );
  ISOLANDX1 U6030 ( .D(WX7230), .ISO(n4629), .Q(WX7293) );
  ISOLANDX1 U6031 ( .D(WX7228), .ISO(n4629), .Q(WX7291) );
  ISOLANDX1 U6032 ( .D(WX7226), .ISO(n4630), .Q(WX7289) );
  ISOLANDX1 U6033 ( .D(WX7224), .ISO(n4630), .Q(WX7287) );
  ISOLANDX1 U6034 ( .D(WX7222), .ISO(n4630), .Q(WX7285) );
  ISOLANDX1 U6035 ( .D(test_so60), .ISO(n4630), .Q(WX7283) );
  ISOLANDX1 U6036 ( .D(WX7218), .ISO(n4630), .Q(WX7281) );
  ISOLANDX1 U6037 ( .D(WX7216), .ISO(n4630), .Q(WX7279) );
  ISOLANDX1 U6038 ( .D(WX7214), .ISO(n4630), .Q(WX7277) );
  ISOLANDX1 U6039 ( .D(WX7212), .ISO(n4630), .Q(WX7275) );
  ISOLANDX1 U6040 ( .D(WX7210), .ISO(n4630), .Q(WX7273) );
  ISOLANDX1 U6041 ( .D(WX7208), .ISO(n4630), .Q(WX7271) );
  ISOLANDX1 U6042 ( .D(WX7206), .ISO(n4630), .Q(WX7269) );
  ISOLANDX1 U6043 ( .D(WX7204), .ISO(n4630), .Q(WX7267) );
  ISOLANDX1 U6044 ( .D(WX7202), .ISO(n4630), .Q(WX7265) );
  ISOLANDX1 U6045 ( .D(WX7200), .ISO(n4630), .Q(WX7263) );
  ISOLANDX1 U6046 ( .D(WX7198), .ISO(n4631), .Q(WX7261) );
  ISOLANDX1 U6047 ( .D(WX7196), .ISO(n4631), .Q(WX7259) );
  ISOLANDX1 U6048 ( .D(WX7194), .ISO(n4631), .Q(WX7257) );
  ISOLANDX1 U6049 ( .D(WX7192), .ISO(n4631), .Q(WX7255) );
  ISOLANDX1 U6050 ( .D(WX7190), .ISO(n4631), .Q(WX7253) );
  ISOLANDX1 U6051 ( .D(WX7188), .ISO(n4631), .Q(WX7251) );
  ISOLANDX1 U6052 ( .D(test_so59), .ISO(n4631), .Q(WX7249) );
  ISOLANDX1 U6053 ( .D(WX7184), .ISO(n4631), .Q(WX7247) );
  ISOLANDX1 U6054 ( .D(WX7182), .ISO(n4631), .Q(WX7245) );
  ISOLANDX1 U6055 ( .D(WX7180), .ISO(n4631), .Q(WX7243) );
  ISOLANDX1 U6056 ( .D(WX7178), .ISO(n4631), .Q(WX7241) );
  ISOLANDX1 U6057 ( .D(WX7176), .ISO(n4631), .Q(WX7239) );
  ISOLANDX1 U6058 ( .D(WX7174), .ISO(n4631), .Q(WX7237) );
  ISOLANDX1 U6059 ( .D(WX7172), .ISO(n4632), .Q(WX7235) );
  ISOLANDX1 U6060 ( .D(WX7170), .ISO(n4632), .Q(WX7233) );
  ISOLANDX1 U6061 ( .D(WX7168), .ISO(n4632), .Q(WX7231) );
  ISOLANDX1 U6062 ( .D(WX7166), .ISO(n4632), .Q(WX7229) );
  ISOLANDX1 U6063 ( .D(WX7164), .ISO(n4632), .Q(WX7227) );
  ISOLANDX1 U6064 ( .D(WX7162), .ISO(n4632), .Q(WX7225) );
  ISOLANDX1 U6065 ( .D(WX7160), .ISO(n4632), .Q(WX7223) );
  ISOLANDX1 U6066 ( .D(WX7158), .ISO(n4632), .Q(WX7221) );
  ISOLANDX1 U6067 ( .D(WX7156), .ISO(n4632), .Q(WX7219) );
  ISOLANDX1 U6068 ( .D(WX7154), .ISO(n4632), .Q(WX7217) );
  ISOLANDX1 U6069 ( .D(test_so58), .ISO(n4632), .Q(WX7215) );
  ISOLANDX1 U6070 ( .D(WX7150), .ISO(n4632), .Q(WX7213) );
  ISOLANDX1 U6071 ( .D(WX7148), .ISO(n4632), .Q(WX7211) );
  ISOLANDX1 U6072 ( .D(WX7146), .ISO(n4632), .Q(WX7209) );
  ISOLANDX1 U6073 ( .D(WX7144), .ISO(n4633), .Q(WX7207) );
  ISOLANDX1 U6074 ( .D(WX7142), .ISO(n4633), .Q(WX7205) );
  ISOLANDX1 U6075 ( .D(WX6007), .ISO(n4635), .Q(WX6070) );
  ISOLANDX1 U6076 ( .D(test_so51), .ISO(n4635), .Q(WX6068) );
  ISOLANDX1 U6077 ( .D(WX6003), .ISO(n4635), .Q(WX6066) );
  ISOLANDX1 U6078 ( .D(WX6001), .ISO(n4635), .Q(WX6064) );
  ISOLANDX1 U6079 ( .D(WX5999), .ISO(n4636), .Q(WX6062) );
  ISOLANDX1 U6080 ( .D(WX5997), .ISO(n4636), .Q(WX6060) );
  ISOLANDX1 U6081 ( .D(WX5995), .ISO(n4636), .Q(WX6058) );
  ISOLANDX1 U6082 ( .D(WX5993), .ISO(n4636), .Q(WX6056) );
  ISOLANDX1 U6083 ( .D(WX5991), .ISO(n4636), .Q(WX6054) );
  ISOLANDX1 U6084 ( .D(WX5989), .ISO(n4636), .Q(WX6052) );
  ISOLANDX1 U6085 ( .D(WX5987), .ISO(n4636), .Q(WX6050) );
  ISOLANDX1 U6086 ( .D(WX5985), .ISO(n4636), .Q(WX6048) );
  ISOLANDX1 U6087 ( .D(WX5983), .ISO(n4636), .Q(WX6046) );
  ISOLANDX1 U6088 ( .D(WX5981), .ISO(n4636), .Q(WX6044) );
  ISOLANDX1 U6089 ( .D(WX5979), .ISO(n4636), .Q(WX6042) );
  ISOLANDX1 U6090 ( .D(WX5977), .ISO(n4636), .Q(WX6040) );
  ISOLANDX1 U6091 ( .D(WX5975), .ISO(n4636), .Q(WX6038) );
  ISOLANDX1 U6092 ( .D(WX5973), .ISO(n4636), .Q(WX6036) );
  ISOLANDX1 U6093 ( .D(test_so50), .ISO(n4636), .Q(WX6034) );
  ISOLANDX1 U6094 ( .D(WX5969), .ISO(n4637), .Q(WX6032) );
  ISOLANDX1 U6095 ( .D(WX5967), .ISO(n4637), .Q(WX6030) );
  ISOLANDX1 U6096 ( .D(WX5965), .ISO(n4637), .Q(WX6028) );
  ISOLANDX1 U6097 ( .D(WX5963), .ISO(n4637), .Q(WX6026) );
  ISOLANDX1 U6098 ( .D(WX5961), .ISO(n4637), .Q(WX6024) );
  ISOLANDX1 U6099 ( .D(WX5959), .ISO(n4637), .Q(WX6022) );
  ISOLANDX1 U6100 ( .D(WX5957), .ISO(n4637), .Q(WX6020) );
  ISOLANDX1 U6101 ( .D(WX5955), .ISO(n4637), .Q(WX6018) );
  ISOLANDX1 U6102 ( .D(WX5953), .ISO(n4637), .Q(WX6016) );
  ISOLANDX1 U6103 ( .D(WX5951), .ISO(n4637), .Q(WX6014) );
  ISOLANDX1 U6104 ( .D(WX5949), .ISO(n4637), .Q(WX6012) );
  ISOLANDX1 U6105 ( .D(WX5947), .ISO(n4637), .Q(WX6010) );
  ISOLANDX1 U6106 ( .D(WX5945), .ISO(n4637), .Q(WX6008) );
  ISOLANDX1 U6107 ( .D(WX5943), .ISO(n4637), .Q(WX6006) );
  ISOLANDX1 U6108 ( .D(WX5941), .ISO(n4637), .Q(WX6004) );
  ISOLANDX1 U6109 ( .D(WX5929), .ISO(n4622), .Q(WX5992) );
  ISOLANDX1 U6110 ( .D(WX5927), .ISO(n4617), .Q(WX5990) );
  ISOLANDX1 U6111 ( .D(WX5925), .ISO(n4617), .Q(WX5988) );
  ISOLANDX1 U6112 ( .D(WX5923), .ISO(n4617), .Q(WX5986) );
  ISOLANDX1 U6113 ( .D(WX5921), .ISO(n4617), .Q(WX5984) );
  ISOLANDX1 U6114 ( .D(WX5919), .ISO(n4617), .Q(WX5982) );
  ISOLANDX1 U6115 ( .D(WX5917), .ISO(n4618), .Q(WX5980) );
  ISOLANDX1 U6116 ( .D(WX5915), .ISO(n4618), .Q(WX5978) );
  ISOLANDX1 U6117 ( .D(WX5913), .ISO(n4618), .Q(WX5976) );
  ISOLANDX1 U6118 ( .D(WX5911), .ISO(n4618), .Q(WX5974) );
  ISOLANDX1 U6119 ( .D(WX5909), .ISO(n4618), .Q(WX5972) );
  ISOLANDX1 U6120 ( .D(WX5907), .ISO(n4618), .Q(WX5970) );
  ISOLANDX1 U6121 ( .D(WX5905), .ISO(n4618), .Q(WX5968) );
  ISOLANDX1 U6122 ( .D(test_so48), .ISO(n4618), .Q(WX5966) );
  ISOLANDX1 U6123 ( .D(WX5901), .ISO(n4618), .Q(WX5964) );
  ISOLANDX1 U6124 ( .D(WX5899), .ISO(n4618), .Q(WX5962) );
  ISOLANDX1 U6125 ( .D(WX5897), .ISO(n4618), .Q(WX5960) );
  ISOLANDX1 U6126 ( .D(WX5895), .ISO(n4618), .Q(WX5958) );
  ISOLANDX1 U6127 ( .D(WX5893), .ISO(n4618), .Q(WX5956) );
  ISOLANDX1 U6128 ( .D(WX5891), .ISO(n4618), .Q(WX5954) );
  ISOLANDX1 U6129 ( .D(WX5889), .ISO(n4618), .Q(WX5952) );
  ISOLANDX1 U6130 ( .D(WX5887), .ISO(n4619), .Q(WX5950) );
  ISOLANDX1 U6131 ( .D(WX5885), .ISO(n4619), .Q(WX5948) );
  ISOLANDX1 U6132 ( .D(WX5883), .ISO(n4619), .Q(WX5946) );
  ISOLANDX1 U6133 ( .D(WX5881), .ISO(n4619), .Q(WX5944) );
  ISOLANDX1 U6134 ( .D(WX5879), .ISO(n4619), .Q(WX5942) );
  ISOLANDX1 U6135 ( .D(WX5877), .ISO(n4619), .Q(WX5940) );
  ISOLANDX1 U6136 ( .D(WX5875), .ISO(n4619), .Q(WX5938) );
  ISOLANDX1 U6137 ( .D(WX5873), .ISO(n4619), .Q(WX5936) );
  ISOLANDX1 U6138 ( .D(WX5871), .ISO(n4619), .Q(WX5934) );
  ISOLANDX1 U6139 ( .D(test_so47), .ISO(n4619), .Q(WX5932) );
  ISOLANDX1 U6140 ( .D(WX5867), .ISO(n4619), .Q(WX5930) );
  ISOLANDX1 U6141 ( .D(WX5865), .ISO(n4619), .Q(WX5928) );
  ISOLANDX1 U6142 ( .D(WX5863), .ISO(n4619), .Q(WX5926) );
  ISOLANDX1 U6143 ( .D(WX5861), .ISO(n4619), .Q(WX5924) );
  ISOLANDX1 U6144 ( .D(WX5859), .ISO(n4619), .Q(WX5922) );
  ISOLANDX1 U6145 ( .D(WX5857), .ISO(n4620), .Q(WX5920) );
  ISOLANDX1 U6146 ( .D(WX5855), .ISO(n4620), .Q(WX5918) );
  ISOLANDX1 U6147 ( .D(WX5853), .ISO(n4620), .Q(WX5916) );
  ISOLANDX1 U6148 ( .D(WX5851), .ISO(n4620), .Q(WX5914) );
  ISOLANDX1 U6149 ( .D(WX5849), .ISO(n4620), .Q(WX5912) );
  ISOLANDX1 U6150 ( .D(WX4714), .ISO(n4624), .Q(WX4777) );
  ISOLANDX1 U6151 ( .D(WX4712), .ISO(n4624), .Q(WX4775) );
  ISOLANDX1 U6152 ( .D(WX4710), .ISO(n4624), .Q(WX4773) );
  ISOLANDX1 U6153 ( .D(WX4708), .ISO(n4624), .Q(WX4771) );
  ISOLANDX1 U6154 ( .D(WX4706), .ISO(n4624), .Q(WX4769) );
  ISOLANDX1 U6155 ( .D(WX4704), .ISO(n4624), .Q(WX4767) );
  ISOLANDX1 U6156 ( .D(WX4702), .ISO(n4624), .Q(WX4765) );
  ISOLANDX1 U6157 ( .D(WX4700), .ISO(n4625), .Q(WX4763) );
  ISOLANDX1 U6158 ( .D(WX4698), .ISO(n4625), .Q(WX4761) );
  ISOLANDX1 U6159 ( .D(WX4696), .ISO(n4625), .Q(WX4759) );
  ISOLANDX1 U6160 ( .D(WX4694), .ISO(n4625), .Q(WX4757) );
  ISOLANDX1 U6161 ( .D(WX4692), .ISO(n4625), .Q(WX4755) );
  ISOLANDX1 U6162 ( .D(WX4690), .ISO(n4625), .Q(WX4753) );
  ISOLANDX1 U6163 ( .D(test_so39), .ISO(n4625), .Q(WX4751) );
  ISOLANDX1 U6164 ( .D(WX4686), .ISO(n4625), .Q(WX4749) );
  ISOLANDX1 U6165 ( .D(WX4684), .ISO(n4625), .Q(WX4747) );
  ISOLANDX1 U6166 ( .D(WX4682), .ISO(n4625), .Q(WX4745) );
  ISOLANDX1 U6167 ( .D(WX4680), .ISO(n4625), .Q(WX4743) );
  ISOLANDX1 U6168 ( .D(WX4678), .ISO(n4625), .Q(WX4741) );
  ISOLANDX1 U6169 ( .D(WX4676), .ISO(n4625), .Q(WX4739) );
  ISOLANDX1 U6170 ( .D(WX4674), .ISO(n4625), .Q(WX4737) );
  ISOLANDX1 U6171 ( .D(WX4672), .ISO(n4625), .Q(WX4735) );
  ISOLANDX1 U6172 ( .D(WX4670), .ISO(n4626), .Q(WX4733) );
  ISOLANDX1 U6173 ( .D(WX4668), .ISO(n4626), .Q(WX4731) );
  ISOLANDX1 U6174 ( .D(WX4666), .ISO(n4626), .Q(WX4729) );
  ISOLANDX1 U6175 ( .D(WX4664), .ISO(n4626), .Q(WX4727) );
  ISOLANDX1 U6176 ( .D(WX4662), .ISO(n4626), .Q(WX4725) );
  ISOLANDX1 U6177 ( .D(WX4660), .ISO(n4626), .Q(WX4723) );
  ISOLANDX1 U6178 ( .D(WX4658), .ISO(n4626), .Q(WX4721) );
  ISOLANDX1 U6179 ( .D(WX4656), .ISO(n4626), .Q(WX4719) );
  ISOLANDX1 U6180 ( .D(test_so38), .ISO(n4626), .Q(WX4717) );
  ISOLANDX1 U6181 ( .D(WX4652), .ISO(n4626), .Q(WX4715) );
  ISOLANDX1 U6182 ( .D(WX4650), .ISO(n4626), .Q(WX4713) );
  ISOLANDX1 U6183 ( .D(WX4648), .ISO(n4626), .Q(WX4711) );
  ISOLANDX1 U6184 ( .D(WX4646), .ISO(n4626), .Q(WX4709) );
  ISOLANDX1 U6185 ( .D(WX4644), .ISO(n4626), .Q(WX4707) );
  ISOLANDX1 U6186 ( .D(WX4642), .ISO(n4626), .Q(WX4705) );
  ISOLANDX1 U6187 ( .D(WX4640), .ISO(n4627), .Q(WX4703) );
  ISOLANDX1 U6188 ( .D(WX4638), .ISO(n4627), .Q(WX4701) );
  ISOLANDX1 U6189 ( .D(WX4636), .ISO(n4627), .Q(WX4699) );
  ISOLANDX1 U6190 ( .D(WX4634), .ISO(n4627), .Q(WX4697) );
  ISOLANDX1 U6191 ( .D(WX4632), .ISO(n4627), .Q(WX4695) );
  ISOLANDX1 U6192 ( .D(WX4630), .ISO(n4627), .Q(WX4693) );
  ISOLANDX1 U6193 ( .D(WX4628), .ISO(n4627), .Q(WX4691) );
  ISOLANDX1 U6194 ( .D(WX4626), .ISO(n4627), .Q(WX4689) );
  ISOLANDX1 U6195 ( .D(WX4624), .ISO(n4627), .Q(WX4687) );
  ISOLANDX1 U6196 ( .D(WX4622), .ISO(n4627), .Q(WX4685) );
  ISOLANDX1 U6197 ( .D(test_so37), .ISO(n4627), .Q(WX4683) );
  ISOLANDX1 U6198 ( .D(WX4618), .ISO(n4627), .Q(WX4681) );
  ISOLANDX1 U6199 ( .D(WX4616), .ISO(n4627), .Q(WX4679) );
  ISOLANDX1 U6200 ( .D(WX4614), .ISO(n4627), .Q(WX4677) );
  ISOLANDX1 U6201 ( .D(WX4612), .ISO(n4627), .Q(WX4675) );
  ISOLANDX1 U6202 ( .D(WX4610), .ISO(n4579), .Q(WX4673) );
  ISOLANDX1 U6203 ( .D(WX4608), .ISO(n4573), .Q(WX4671) );
  ISOLANDX1 U6204 ( .D(WX4606), .ISO(n4573), .Q(WX4669) );
  ISOLANDX1 U6205 ( .D(WX4604), .ISO(n4573), .Q(WX4667) );
  ISOLANDX1 U6206 ( .D(WX4602), .ISO(n4573), .Q(WX4665) );
  ISOLANDX1 U6207 ( .D(WX4600), .ISO(n4573), .Q(WX4663) );
  ISOLANDX1 U6208 ( .D(WX4598), .ISO(n4572), .Q(WX4661) );
  ISOLANDX1 U6209 ( .D(WX4596), .ISO(n4574), .Q(WX4659) );
  ISOLANDX1 U6210 ( .D(WX4594), .ISO(n4574), .Q(WX4657) );
  ISOLANDX1 U6211 ( .D(WX4592), .ISO(n4574), .Q(WX4655) );
  ISOLANDX1 U6212 ( .D(WX4590), .ISO(n4574), .Q(WX4653) );
  ISOLANDX1 U6213 ( .D(WX4588), .ISO(n4574), .Q(WX4651) );
  ISOLANDX1 U6214 ( .D(test_so36), .ISO(n4574), .Q(WX4649) );
  ISOLANDX1 U6215 ( .D(WX4584), .ISO(n4574), .Q(WX4647) );
  ISOLANDX1 U6216 ( .D(WX4582), .ISO(n4574), .Q(WX4645) );
  ISOLANDX1 U6217 ( .D(WX4580), .ISO(n4574), .Q(WX4643) );
  ISOLANDX1 U6218 ( .D(WX4578), .ISO(n4574), .Q(WX4641) );
  ISOLANDX1 U6219 ( .D(WX4576), .ISO(n4574), .Q(WX4639) );
  ISOLANDX1 U6220 ( .D(WX4574), .ISO(n4574), .Q(WX4637) );
  ISOLANDX1 U6221 ( .D(WX4572), .ISO(n4574), .Q(WX4635) );
  ISOLANDX1 U6222 ( .D(WX4570), .ISO(n4575), .Q(WX4633) );
  ISOLANDX1 U6223 ( .D(WX4568), .ISO(n4575), .Q(WX4631) );
  ISOLANDX1 U6224 ( .D(WX4566), .ISO(n4575), .Q(WX4629) );
  ISOLANDX1 U6225 ( .D(WX4564), .ISO(n4575), .Q(WX4627) );
  ISOLANDX1 U6226 ( .D(WX4562), .ISO(n4575), .Q(WX4625) );
  ISOLANDX1 U6227 ( .D(WX4560), .ISO(n4575), .Q(WX4623) );
  ISOLANDX1 U6228 ( .D(WX4558), .ISO(n4575), .Q(WX4621) );
  ISOLANDX1 U6229 ( .D(WX4556), .ISO(n4575), .Q(WX4619) );
  ISOLANDX1 U6230 ( .D(WX3421), .ISO(n4579), .Q(WX3484) );
  ISOLANDX1 U6231 ( .D(WX3419), .ISO(n4579), .Q(WX3482) );
  ISOLANDX1 U6232 ( .D(WX3417), .ISO(n4579), .Q(WX3480) );
  ISOLANDX1 U6233 ( .D(WX3415), .ISO(n4579), .Q(WX3478) );
  ISOLANDX1 U6234 ( .D(WX3413), .ISO(n4579), .Q(WX3476) );
  ISOLANDX1 U6235 ( .D(WX3411), .ISO(n4573), .Q(WX3474) );
  ISOLANDX1 U6236 ( .D(WX3409), .ISO(n4579), .Q(WX3472) );
  ISOLANDX1 U6237 ( .D(WX3407), .ISO(n4579), .Q(WX3470) );
  ISOLANDX1 U6238 ( .D(test_so28), .ISO(n4579), .Q(WX3468) );
  ISOLANDX1 U6239 ( .D(WX3403), .ISO(n4579), .Q(WX3466) );
  ISOLANDX1 U6240 ( .D(WX3401), .ISO(n4579), .Q(WX3464) );
  ISOLANDX1 U6241 ( .D(WX3399), .ISO(n4579), .Q(WX3462) );
  ISOLANDX1 U6242 ( .D(WX3397), .ISO(n4579), .Q(WX3460) );
  ISOLANDX1 U6243 ( .D(WX3395), .ISO(n4579), .Q(WX3458) );
  ISOLANDX1 U6244 ( .D(WX3393), .ISO(n4578), .Q(WX3456) );
  ISOLANDX1 U6245 ( .D(WX3391), .ISO(n4578), .Q(WX3454) );
  ISOLANDX1 U6246 ( .D(WX3389), .ISO(n4578), .Q(WX3452) );
  ISOLANDX1 U6247 ( .D(WX3387), .ISO(n4578), .Q(WX3450) );
  ISOLANDX1 U6248 ( .D(WX3385), .ISO(n4578), .Q(WX3448) );
  ISOLANDX1 U6249 ( .D(WX3383), .ISO(n4578), .Q(WX3446) );
  ISOLANDX1 U6250 ( .D(WX3381), .ISO(n4578), .Q(WX3444) );
  ISOLANDX1 U6251 ( .D(WX3379), .ISO(n4578), .Q(WX3442) );
  ISOLANDX1 U6252 ( .D(WX3377), .ISO(n4578), .Q(WX3440) );
  ISOLANDX1 U6253 ( .D(WX3375), .ISO(n4578), .Q(WX3438) );
  ISOLANDX1 U6254 ( .D(WX3373), .ISO(n4578), .Q(WX3436) );
  ISOLANDX1 U6255 ( .D(WX3371), .ISO(n4578), .Q(WX3434) );
  ISOLANDX1 U6256 ( .D(test_so27), .ISO(n4578), .Q(WX3432) );
  ISOLANDX1 U6257 ( .D(WX3367), .ISO(n4578), .Q(WX3430) );
  ISOLANDX1 U6258 ( .D(WX3365), .ISO(n4578), .Q(WX3428) );
  ISOLANDX1 U6259 ( .D(WX3363), .ISO(n4577), .Q(WX3426) );
  ISOLANDX1 U6260 ( .D(WX3361), .ISO(n4577), .Q(WX3424) );
  ISOLANDX1 U6261 ( .D(WX3359), .ISO(n4577), .Q(WX3422) );
  ISOLANDX1 U6262 ( .D(WX3357), .ISO(n4577), .Q(WX3420) );
  ISOLANDX1 U6263 ( .D(WX3355), .ISO(n4577), .Q(WX3418) );
  ISOLANDX1 U6264 ( .D(WX3353), .ISO(n4577), .Q(WX3416) );
  ISOLANDX1 U6265 ( .D(WX3351), .ISO(n4577), .Q(WX3414) );
  ISOLANDX1 U6266 ( .D(WX3349), .ISO(n4577), .Q(WX3412) );
  ISOLANDX1 U6267 ( .D(WX3347), .ISO(n4577), .Q(WX3410) );
  ISOLANDX1 U6268 ( .D(WX3345), .ISO(n4577), .Q(WX3408) );
  ISOLANDX1 U6269 ( .D(WX3343), .ISO(n4577), .Q(WX3406) );
  ISOLANDX1 U6270 ( .D(WX3341), .ISO(n4577), .Q(WX3404) );
  ISOLANDX1 U6271 ( .D(WX3339), .ISO(n4577), .Q(WX3402) );
  ISOLANDX1 U6272 ( .D(WX3337), .ISO(n4577), .Q(WX3400) );
  ISOLANDX1 U6273 ( .D(WX3335), .ISO(n4577), .Q(WX3398) );
  ISOLANDX1 U6274 ( .D(test_so26), .ISO(n4576), .Q(WX3396) );
  ISOLANDX1 U6275 ( .D(WX3331), .ISO(n4576), .Q(WX3394) );
  ISOLANDX1 U6276 ( .D(WX3329), .ISO(n4576), .Q(WX3392) );
  ISOLANDX1 U6277 ( .D(WX3327), .ISO(n4576), .Q(WX3390) );
  ISOLANDX1 U6278 ( .D(WX3325), .ISO(n4576), .Q(WX3388) );
  ISOLANDX1 U6279 ( .D(WX3323), .ISO(n4576), .Q(WX3386) );
  ISOLANDX1 U6280 ( .D(WX3321), .ISO(n4576), .Q(WX3384) );
  ISOLANDX1 U6281 ( .D(WX3319), .ISO(n4576), .Q(WX3382) );
  ISOLANDX1 U6282 ( .D(WX3317), .ISO(n4576), .Q(WX3380) );
  ISOLANDX1 U6283 ( .D(WX3315), .ISO(n4576), .Q(WX3378) );
  ISOLANDX1 U6284 ( .D(WX3313), .ISO(n4576), .Q(WX3376) );
  ISOLANDX1 U6285 ( .D(WX3311), .ISO(n4576), .Q(WX3374) );
  ISOLANDX1 U6286 ( .D(WX3309), .ISO(n4576), .Q(WX3372) );
  ISOLANDX1 U6287 ( .D(WX3307), .ISO(n4576), .Q(WX3370) );
  ISOLANDX1 U6288 ( .D(WX3305), .ISO(n4576), .Q(WX3368) );
  ISOLANDX1 U6289 ( .D(WX3303), .ISO(n4575), .Q(WX3366) );
  ISOLANDX1 U6290 ( .D(WX3301), .ISO(n4575), .Q(WX3364) );
  ISOLANDX1 U6291 ( .D(WX3299), .ISO(n4575), .Q(WX3362) );
  ISOLANDX1 U6292 ( .D(test_so25), .ISO(n4575), .Q(WX3360) );
  ISOLANDX1 U6293 ( .D(WX3295), .ISO(n4575), .Q(WX3358) );
  ISOLANDX1 U6294 ( .D(WX3293), .ISO(n4575), .Q(WX3356) );
  ISOLANDX1 U6295 ( .D(WX3291), .ISO(n4575), .Q(WX3354) );
  ISOLANDX1 U6296 ( .D(WX3289), .ISO(n4573), .Q(WX3352) );
  ISOLANDX1 U6297 ( .D(WX3287), .ISO(n4573), .Q(WX3350) );
  ISOLANDX1 U6298 ( .D(WX3285), .ISO(n4573), .Q(WX3348) );
  ISOLANDX1 U6299 ( .D(WX3283), .ISO(n4573), .Q(WX3346) );
  ISOLANDX1 U6300 ( .D(WX3281), .ISO(n4573), .Q(WX3344) );
  ISOLANDX1 U6301 ( .D(WX3279), .ISO(n4573), .Q(WX3342) );
  ISOLANDX1 U6302 ( .D(WX3277), .ISO(n4572), .Q(WX3340) );
  ISOLANDX1 U6303 ( .D(WX3275), .ISO(n4573), .Q(WX3338) );
  ISOLANDX1 U6304 ( .D(WX3273), .ISO(n4572), .Q(WX3336) );
  ISOLANDX1 U6305 ( .D(WX3271), .ISO(n4572), .Q(WX3334) );
  ISOLANDX1 U6306 ( .D(WX3267), .ISO(n4574), .Q(WX3330) );
  ISOLANDX1 U6307 ( .D(WX2128), .ISO(n4590), .Q(WX2191) );
  ISOLANDX1 U6308 ( .D(WX2126), .ISO(n4590), .Q(WX2189) );
  ISOLANDX1 U6309 ( .D(WX2124), .ISO(n4590), .Q(WX2187) );
  ISOLANDX1 U6310 ( .D(WX2122), .ISO(n4590), .Q(WX2185) );
  ISOLANDX1 U6311 ( .D(WX2120), .ISO(n4590), .Q(WX2183) );
  ISOLANDX1 U6312 ( .D(WX2118), .ISO(n4590), .Q(WX2181) );
  ISOLANDX1 U6313 ( .D(WX2116), .ISO(n4590), .Q(WX2179) );
  ISOLANDX1 U6314 ( .D(WX2114), .ISO(n4590), .Q(WX2177) );
  ISOLANDX1 U6315 ( .D(WX2112), .ISO(n4590), .Q(WX2175) );
  ISOLANDX1 U6316 ( .D(WX2110), .ISO(n4591), .Q(WX2173) );
  ISOLANDX1 U6317 ( .D(WX2108), .ISO(n4591), .Q(WX2171) );
  ISOLANDX1 U6318 ( .D(WX2106), .ISO(n4591), .Q(WX2169) );
  ISOLANDX1 U6319 ( .D(WX2104), .ISO(n4591), .Q(WX2167) );
  ISOLANDX1 U6320 ( .D(WX2102), .ISO(n4591), .Q(WX2165) );
  ISOLANDX1 U6321 ( .D(test_so17), .ISO(n4591), .Q(WX2163) );
  ISOLANDX1 U6322 ( .D(WX2098), .ISO(n4591), .Q(WX2161) );
  ISOLANDX1 U6323 ( .D(WX2096), .ISO(n4591), .Q(WX2159) );
  ISOLANDX1 U6324 ( .D(WX2094), .ISO(n4591), .Q(WX2157) );
  ISOLANDX1 U6325 ( .D(WX2092), .ISO(n4591), .Q(WX2155) );
  ISOLANDX1 U6326 ( .D(WX2090), .ISO(n4591), .Q(WX2153) );
  ISOLANDX1 U6327 ( .D(WX2088), .ISO(n4591), .Q(WX2151) );
  ISOLANDX1 U6328 ( .D(WX2086), .ISO(n4591), .Q(WX2149) );
  ISOLANDX1 U6329 ( .D(WX2084), .ISO(n4591), .Q(WX2147) );
  ISOLANDX1 U6330 ( .D(WX2082), .ISO(n4591), .Q(WX2145) );
  ISOLANDX1 U6331 ( .D(WX2080), .ISO(n4592), .Q(WX2143) );
  ISOLANDX1 U6332 ( .D(WX2078), .ISO(n4592), .Q(WX2141) );
  ISOLANDX1 U6333 ( .D(WX2076), .ISO(n4592), .Q(WX2139) );
  ISOLANDX1 U6334 ( .D(WX2074), .ISO(n4592), .Q(WX2137) );
  ISOLANDX1 U6335 ( .D(WX2072), .ISO(n4592), .Q(WX2135) );
  ISOLANDX1 U6336 ( .D(WX2070), .ISO(n4592), .Q(WX2133) );
  ISOLANDX1 U6337 ( .D(WX2068), .ISO(n4592), .Q(WX2131) );
  ISOLANDX1 U6338 ( .D(WX2066), .ISO(n4592), .Q(WX2129) );
  ISOLANDX1 U6339 ( .D(test_so16), .ISO(n4592), .Q(WX2127) );
  ISOLANDX1 U6340 ( .D(WX2062), .ISO(n4592), .Q(WX2125) );
  ISOLANDX1 U6341 ( .D(WX2060), .ISO(n4592), .Q(WX2123) );
  ISOLANDX1 U6342 ( .D(WX2058), .ISO(n4592), .Q(WX2121) );
  ISOLANDX1 U6343 ( .D(WX2056), .ISO(n4592), .Q(WX2119) );
  ISOLANDX1 U6344 ( .D(WX2054), .ISO(n4592), .Q(WX2117) );
  ISOLANDX1 U6345 ( .D(WX2052), .ISO(n4593), .Q(WX2115) );
  ISOLANDX1 U6346 ( .D(WX2050), .ISO(n4593), .Q(WX2113) );
  ISOLANDX1 U6347 ( .D(WX2048), .ISO(n4593), .Q(WX2111) );
  ISOLANDX1 U6348 ( .D(WX2046), .ISO(n4593), .Q(WX2109) );
  ISOLANDX1 U6349 ( .D(WX2044), .ISO(n4593), .Q(WX2107) );
  ISOLANDX1 U6350 ( .D(WX2042), .ISO(n4593), .Q(WX2105) );
  ISOLANDX1 U6351 ( .D(WX2040), .ISO(n4593), .Q(WX2103) );
  ISOLANDX1 U6352 ( .D(WX2038), .ISO(n4593), .Q(WX2101) );
  ISOLANDX1 U6353 ( .D(WX2036), .ISO(n4593), .Q(WX2099) );
  ISOLANDX1 U6354 ( .D(WX2034), .ISO(n4593), .Q(WX2097) );
  ISOLANDX1 U6355 ( .D(WX2032), .ISO(n4593), .Q(WX2095) );
  ISOLANDX1 U6356 ( .D(WX2030), .ISO(n4593), .Q(WX2093) );
  ISOLANDX1 U6357 ( .D(test_so15), .ISO(n4593), .Q(WX2091) );
  ISOLANDX1 U6358 ( .D(WX2026), .ISO(n4593), .Q(WX2089) );
  ISOLANDX1 U6359 ( .D(WX2024), .ISO(n4593), .Q(WX2087) );
  ISOLANDX1 U6360 ( .D(WX2022), .ISO(n4594), .Q(WX2085) );
  ISOLANDX1 U6361 ( .D(WX2020), .ISO(n4594), .Q(WX2083) );
  ISOLANDX1 U6362 ( .D(WX2018), .ISO(n4594), .Q(WX2081) );
  ISOLANDX1 U6363 ( .D(WX2016), .ISO(n4594), .Q(WX2079) );
  ISOLANDX1 U6364 ( .D(WX2014), .ISO(n4594), .Q(WX2077) );
  ISOLANDX1 U6365 ( .D(WX2012), .ISO(n4594), .Q(WX2075) );
  ISOLANDX1 U6366 ( .D(WX2010), .ISO(n4594), .Q(WX2073) );
  ISOLANDX1 U6367 ( .D(WX2008), .ISO(n4594), .Q(WX2071) );
  ISOLANDX1 U6368 ( .D(WX2006), .ISO(n4594), .Q(WX2069) );
  ISOLANDX1 U6369 ( .D(WX2004), .ISO(n4594), .Q(WX2067) );
  ISOLANDX1 U6370 ( .D(WX2002), .ISO(n4594), .Q(WX2065) );
  ISOLANDX1 U6371 ( .D(WX2000), .ISO(n4594), .Q(WX2063) );
  ISOLANDX1 U6372 ( .D(WX1998), .ISO(n4594), .Q(WX2061) );
  ISOLANDX1 U6373 ( .D(WX1996), .ISO(n4594), .Q(WX2059) );
  ISOLANDX1 U6374 ( .D(WX1994), .ISO(n4594), .Q(WX2057) );
  ISOLANDX1 U6375 ( .D(test_so14), .ISO(n4595), .Q(WX2055) );
  ISOLANDX1 U6376 ( .D(WX1990), .ISO(n4595), .Q(WX2053) );
  ISOLANDX1 U6377 ( .D(WX1988), .ISO(n4595), .Q(WX2051) );
  ISOLANDX1 U6378 ( .D(WX1986), .ISO(n4595), .Q(WX2049) );
  ISOLANDX1 U6379 ( .D(WX1984), .ISO(n4595), .Q(WX2047) );
  ISOLANDX1 U6380 ( .D(WX1982), .ISO(n4595), .Q(WX2045) );
  ISOLANDX1 U6381 ( .D(WX1980), .ISO(n4595), .Q(WX2043) );
  ISOLANDX1 U6382 ( .D(WX1978), .ISO(n4595), .Q(WX2041) );
  ISOLANDX1 U6383 ( .D(WX1976), .ISO(n4595), .Q(WX2039) );
  ISOLANDX1 U6384 ( .D(WX1974), .ISO(n4595), .Q(WX2037) );
  ISOLANDX1 U6385 ( .D(WX1972), .ISO(n4595), .Q(WX2035) );
  ISOLANDX1 U6386 ( .D(WX1970), .ISO(n4595), .Q(WX2033) );
  ISOLANDX1 U6387 ( .D(WX835), .ISO(n4614), .Q(WX898) );
  ISOLANDX1 U6388 ( .D(WX833), .ISO(n4614), .Q(WX896) );
  ISOLANDX1 U6389 ( .D(test_so7), .ISO(n4614), .Q(WX894) );
  ISOLANDX1 U6390 ( .D(WX829), .ISO(n4614), .Q(WX892) );
  ISOLANDX1 U6391 ( .D(WX827), .ISO(n4614), .Q(WX890) );
  ISOLANDX1 U6392 ( .D(WX825), .ISO(n4614), .Q(WX888) );
  ISOLANDX1 U6393 ( .D(WX823), .ISO(n4614), .Q(WX886) );
  ISOLANDX1 U6394 ( .D(WX821), .ISO(n4614), .Q(WX884) );
  ISOLANDX1 U6395 ( .D(WX819), .ISO(n4615), .Q(WX882) );
  ISOLANDX1 U6396 ( .D(WX817), .ISO(n4615), .Q(WX880) );
  ISOLANDX1 U6397 ( .D(WX815), .ISO(n4615), .Q(WX878) );
  ISOLANDX1 U6398 ( .D(WX813), .ISO(n4615), .Q(WX876) );
  ISOLANDX1 U6399 ( .D(WX811), .ISO(n4615), .Q(WX874) );
  ISOLANDX1 U6400 ( .D(WX809), .ISO(n4615), .Q(WX872) );
  ISOLANDX1 U6401 ( .D(WX807), .ISO(n4615), .Q(WX870) );
  ISOLANDX1 U6402 ( .D(WX805), .ISO(n4615), .Q(WX868) );
  ISOLANDX1 U6403 ( .D(WX803), .ISO(n4615), .Q(WX866) );
  ISOLANDX1 U6404 ( .D(WX801), .ISO(n4616), .Q(WX864) );
  ISOLANDX1 U6405 ( .D(WX799), .ISO(n4616), .Q(WX862) );
  ISOLANDX1 U6406 ( .D(WX797), .ISO(n4596), .Q(WX860) );
  ISOLANDX1 U6407 ( .D(test_so6), .ISO(n4597), .Q(WX858) );
  ISOLANDX1 U6408 ( .D(WX793), .ISO(n4598), .Q(WX856) );
  ISOLANDX1 U6409 ( .D(WX791), .ISO(n4599), .Q(WX854) );
  ISOLANDX1 U6410 ( .D(WX789), .ISO(n4599), .Q(WX852) );
  ISOLANDX1 U6411 ( .D(WX787), .ISO(n4600), .Q(WX850) );
  ISOLANDX1 U6412 ( .D(WX785), .ISO(n4600), .Q(WX848) );
  ISOLANDX1 U6413 ( .D(WX783), .ISO(n4600), .Q(WX846) );
  ISOLANDX1 U6414 ( .D(WX781), .ISO(n4600), .Q(WX844) );
  ISOLANDX1 U6415 ( .D(WX779), .ISO(n4600), .Q(WX842) );
  ISOLANDX1 U6416 ( .D(WX777), .ISO(n4601), .Q(WX840) );
  ISOLANDX1 U6417 ( .D(WX775), .ISO(n4601), .Q(WX838) );
  ISOLANDX1 U6418 ( .D(WX773), .ISO(n4601), .Q(WX836) );
  ISOLANDX1 U6419 ( .D(WX771), .ISO(n4601), .Q(WX834) );
  ISOLANDX1 U6420 ( .D(WX769), .ISO(n4601), .Q(WX832) );
  ISOLANDX1 U6421 ( .D(WX767), .ISO(n4601), .Q(WX830) );
  ISOLANDX1 U6422 ( .D(WX765), .ISO(n4602), .Q(WX828) );
  ISOLANDX1 U6423 ( .D(WX763), .ISO(n4603), .Q(WX826) );
  ISOLANDX1 U6424 ( .D(WX761), .ISO(n4603), .Q(WX824) );
  ISOLANDX1 U6425 ( .D(test_so5), .ISO(n4603), .Q(WX822) );
  ISOLANDX1 U6426 ( .D(WX757), .ISO(n4603), .Q(WX820) );
  ISOLANDX1 U6427 ( .D(WX755), .ISO(n4603), .Q(WX818) );
  ISOLANDX1 U6428 ( .D(WX753), .ISO(n4603), .Q(WX816) );
  ISOLANDX1 U6429 ( .D(WX751), .ISO(n4604), .Q(WX814) );
  ISOLANDX1 U6430 ( .D(WX749), .ISO(n4604), .Q(WX812) );
  ISOLANDX1 U6431 ( .D(WX747), .ISO(n4604), .Q(WX810) );
  ISOLANDX1 U6432 ( .D(WX745), .ISO(n4604), .Q(WX808) );
  ISOLANDX1 U6433 ( .D(WX743), .ISO(n4604), .Q(WX806) );
  ISOLANDX1 U6434 ( .D(WX741), .ISO(n4604), .Q(WX804) );
  ISOLANDX1 U6435 ( .D(WX739), .ISO(n4604), .Q(WX802) );
  ISOLANDX1 U6436 ( .D(WX737), .ISO(n4604), .Q(WX800) );
  ISOLANDX1 U6437 ( .D(WX735), .ISO(n4604), .Q(WX798) );
  ISOLANDX1 U6438 ( .D(WX733), .ISO(n4604), .Q(WX796) );
  ISOLANDX1 U6439 ( .D(WX731), .ISO(n4604), .Q(WX794) );
  ISOLANDX1 U6440 ( .D(WX729), .ISO(n4604), .Q(WX792) );
  ISOLANDX1 U6441 ( .D(WX727), .ISO(n4604), .Q(WX790) );
  ISOLANDX1 U6442 ( .D(WX725), .ISO(n4604), .Q(WX788) );
  ISOLANDX1 U6443 ( .D(test_so4), .ISO(n4604), .Q(WX786) );
  ISOLANDX1 U6444 ( .D(WX721), .ISO(n4605), .Q(WX784) );
  ISOLANDX1 U6445 ( .D(WX719), .ISO(n4605), .Q(WX782) );
  ISOLANDX1 U6446 ( .D(WX717), .ISO(n4605), .Q(WX780) );
  ISOLANDX1 U6447 ( .D(WX715), .ISO(n4605), .Q(WX778) );
  ISOLANDX1 U6448 ( .D(WX713), .ISO(n4605), .Q(WX776) );
  ISOLANDX1 U6449 ( .D(WX711), .ISO(n4605), .Q(WX774) );
  ISOLANDX1 U6450 ( .D(WX709), .ISO(n4605), .Q(WX772) );
  ISOLANDX1 U6451 ( .D(WX707), .ISO(n4605), .Q(WX770) );
  ISOLANDX1 U6452 ( .D(WX705), .ISO(n4605), .Q(WX768) );
  ISOLANDX1 U6453 ( .D(WX703), .ISO(n4605), .Q(WX766) );
  ISOLANDX1 U6454 ( .D(WX701), .ISO(n4605), .Q(WX764) );
  ISOLANDX1 U6455 ( .D(WX699), .ISO(n4605), .Q(WX762) );
  ISOLANDX1 U6456 ( .D(WX697), .ISO(n4605), .Q(WX760) );
  ISOLANDX1 U6457 ( .D(WX695), .ISO(n4605), .Q(WX758) );
  ISOLANDX1 U6458 ( .D(WX693), .ISO(n4605), .Q(WX756) );
  ISOLANDX1 U6459 ( .D(WX691), .ISO(n4606), .Q(WX754) );
  ISOLANDX1 U6460 ( .D(WX689), .ISO(n4606), .Q(WX752) );
  ISOLANDX1 U6461 ( .D(test_so3), .ISO(n4606), .Q(WX750) );
  ISOLANDX1 U6462 ( .D(WX685), .ISO(n4606), .Q(WX748) );
  ISOLANDX1 U6463 ( .D(WX683), .ISO(n4606), .Q(WX746) );
  ISOLANDX1 U6464 ( .D(WX681), .ISO(n4606), .Q(WX744) );
  ISOLANDX1 U6465 ( .D(WX679), .ISO(n4606), .Q(WX742) );
  ISOLANDX1 U6466 ( .D(WX677), .ISO(n4606), .Q(WX740) );
  ISOLANDX1 U6467 ( .D(WX675), .ISO(n4606), .Q(WX738) );
  ISOLANDX1 U6468 ( .D(WX673), .ISO(n4606), .Q(WX736) );
  ISOLANDX1 U6469 ( .D(WX671), .ISO(n4628), .Q(WX734) );
  ISOLANDX1 U6470 ( .D(WX669), .ISO(n4628), .Q(WX732) );
  ISOLANDX1 U6471 ( .D(WX667), .ISO(n4629), .Q(WX730) );
  ISOLANDX1 U6472 ( .D(WX665), .ISO(n4630), .Q(WX728) );
  ISOLANDX1 U6473 ( .D(WX663), .ISO(n4631), .Q(WX726) );
  ISOLANDX1 U6474 ( .D(WX661), .ISO(n4631), .Q(WX724) );
  ISOLANDX1 U6475 ( .D(WX659), .ISO(n4632), .Q(WX722) );
  ISOLANDX1 U6476 ( .D(WX657), .ISO(n4633), .Q(WX720) );
  ISOLANDX1 U6477 ( .D(WX655), .ISO(n4633), .Q(WX718) );
  ISOLANDX1 U6478 ( .D(WX653), .ISO(n4633), .Q(WX716) );
  ISOLANDX1 U6479 ( .D(test_so2), .ISO(n4633), .Q(WX714) );
  ISOLANDX1 U6480 ( .D(WX649), .ISO(n4633), .Q(WX712) );
  ISOLANDX1 U6481 ( .D(WX647), .ISO(n4633), .Q(WX710) );
  ISOLANDX1 U6482 ( .D(WX645), .ISO(n4633), .Q(WX708) );
  NOR2X0 U6483 ( .IN1(WX485), .IN2(n4536), .QN(WX546) );
  NOR2X0 U6484 ( .IN1(WX10829), .IN2(n4548), .QN(WX10890) );
  NOR2X0 U6485 ( .IN1(WX9536), .IN2(n4548), .QN(WX9597) );
  NOR2X0 U6486 ( .IN1(WX8243), .IN2(n4536), .QN(WX8304) );
  NOR2X0 U6487 ( .IN1(WX6950), .IN2(n4545), .QN(WX7011) );
  NOR2X0 U6488 ( .IN1(WX5657), .IN2(n4539), .QN(WX5718) );
  NOR2X0 U6489 ( .IN1(WX4364), .IN2(n4548), .QN(WX4425) );
  NOR2X0 U6490 ( .IN1(WX3071), .IN2(n4546), .QN(WX3132) );
  NOR2X0 U6491 ( .IN1(WX1778), .IN2(n4539), .QN(WX1839) );
  NOR2X0 U6492 ( .IN1(n4567), .IN2(n3178), .QN(WX11640) );
  XNOR3X1 U6493 ( .IN1(WX11211), .IN2(CRC_OUT_1_31), .IN3(DFF_1711_n1), .Q(
        n3178) );
  NOR2X0 U6494 ( .IN1(n4567), .IN2(n3185), .QN(WX11630) );
  XNOR3X1 U6495 ( .IN1(WX11221), .IN2(CRC_OUT_1_31), .IN3(DFF_1706_n1), .Q(
        n3185) );
  NOR2X0 U6496 ( .IN1(n4567), .IN2(n3192), .QN(WX11616) );
  XNOR3X1 U6497 ( .IN1(WX11235), .IN2(CRC_OUT_1_31), .IN3(DFF_1699_n1), .Q(
        n3192) );
  NOR2X0 U6498 ( .IN1(n4563), .IN2(n3313), .QN(WX10347) );
  XNOR3X1 U6499 ( .IN1(WX9918), .IN2(CRC_OUT_2_31), .IN3(DFF_1519_n1), .Q(
        n3313) );
  NOR2X0 U6500 ( .IN1(n4563), .IN2(n3318), .QN(WX10337) );
  XNOR3X1 U6501 ( .IN1(WX9928), .IN2(CRC_OUT_2_31), .IN3(DFF_1514_n1), .Q(
        n3318) );
  NOR2X0 U6502 ( .IN1(n4562), .IN2(n3325), .QN(WX10323) );
  XNOR3X1 U6503 ( .IN1(WX9942), .IN2(CRC_OUT_2_31), .IN3(DFF_1507_n1), .Q(
        n3325) );
  NOR2X0 U6504 ( .IN1(n4567), .IN2(n2264), .QN(WX9054) );
  XNOR3X1 U6505 ( .IN1(WX8625), .IN2(CRC_OUT_3_31), .IN3(DFF_1327_n1), .Q(
        n2264) );
  NOR2X0 U6506 ( .IN1(n4567), .IN2(n2269), .QN(WX9044) );
  XNOR3X1 U6507 ( .IN1(WX8635), .IN2(CRC_OUT_3_31), .IN3(DFF_1322_n1), .Q(
        n2269) );
  NOR2X0 U6508 ( .IN1(n4567), .IN2(n2276), .QN(WX9030) );
  XNOR3X1 U6509 ( .IN1(WX8649), .IN2(CRC_OUT_3_31), .IN3(DFF_1315_n1), .Q(
        n2276) );
  NOR2X0 U6510 ( .IN1(n4557), .IN2(n2392), .QN(WX7761) );
  XNOR3X1 U6511 ( .IN1(WX7332), .IN2(CRC_OUT_4_31), .IN3(DFF_1135_n1), .Q(
        n2392) );
  NOR2X0 U6512 ( .IN1(n4558), .IN2(n2397), .QN(WX7751) );
  XNOR3X1 U6513 ( .IN1(WX7342), .IN2(CRC_OUT_4_31), .IN3(DFF_1130_n1), .Q(
        n2397) );
  NOR2X0 U6514 ( .IN1(n4558), .IN2(n2404), .QN(WX7737) );
  XNOR3X1 U6515 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .IN3(DFF_1123_n1), .Q(
        n2404) );
  NOR2X0 U6516 ( .IN1(n4562), .IN2(n2610), .QN(WX6468) );
  XNOR3X1 U6517 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .IN3(DFF_943_n1), .Q(
        n2610) );
  NOR2X0 U6518 ( .IN1(n4562), .IN2(n2618), .QN(WX6458) );
  XNOR3X1 U6519 ( .IN1(WX6049), .IN2(CRC_OUT_5_31), .IN3(DFF_938_n1), .Q(n2618) );
  NOR2X0 U6520 ( .IN1(n4562), .IN2(n2625), .QN(WX6444) );
  XNOR3X1 U6521 ( .IN1(WX6063), .IN2(CRC_OUT_5_31), .IN3(DFF_931_n1), .Q(n2625) );
  NOR2X0 U6522 ( .IN1(n4571), .IN2(n2744), .QN(WX5175) );
  XNOR3X1 U6523 ( .IN1(WX4746), .IN2(CRC_OUT_6_31), .IN3(DFF_751_n1), .Q(n2744) );
  NOR2X0 U6524 ( .IN1(n4567), .IN2(n2749), .QN(WX5165) );
  XNOR3X1 U6525 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .IN3(DFF_746_n1), .Q(
        n2749) );
  NOR2X0 U6526 ( .IN1(n4567), .IN2(n2756), .QN(WX5151) );
  XNOR3X1 U6527 ( .IN1(WX4770), .IN2(CRC_OUT_6_31), .IN3(DFF_739_n1), .Q(n2756) );
  NOR2X0 U6528 ( .IN1(n4564), .IN2(n2872), .QN(WX3882) );
  XNOR3X1 U6529 ( .IN1(WX3453), .IN2(CRC_OUT_7_31), .IN3(DFF_559_n1), .Q(n2872) );
  NOR2X0 U6530 ( .IN1(n4565), .IN2(n2877), .QN(WX3872) );
  XNOR3X1 U6531 ( .IN1(WX3463), .IN2(CRC_OUT_7_31), .IN3(DFF_554_n1), .Q(n2877) );
  NOR2X0 U6532 ( .IN1(n4568), .IN2(n2884), .QN(WX3858) );
  XNOR3X1 U6533 ( .IN1(WX3477), .IN2(CRC_OUT_7_31), .IN3(DFF_547_n1), .Q(n2884) );
  NOR2X0 U6534 ( .IN1(n4560), .IN2(n3000), .QN(WX2589) );
  XNOR3X1 U6535 ( .IN1(WX2160), .IN2(CRC_OUT_8_31), .IN3(DFF_367_n1), .Q(n3000) );
  NOR2X0 U6536 ( .IN1(n4560), .IN2(n3005), .QN(WX2579) );
  XNOR3X1 U6537 ( .IN1(WX2170), .IN2(CRC_OUT_8_31), .IN3(DFF_362_n1), .Q(n3005) );
  NOR2X0 U6538 ( .IN1(n4560), .IN2(n3012), .QN(WX2565) );
  XNOR3X1 U6539 ( .IN1(WX2184), .IN2(CRC_OUT_8_31), .IN3(DFF_355_n1), .Q(n3012) );
  NOR2X0 U6540 ( .IN1(n4566), .IN2(n3128), .QN(WX1296) );
  XNOR3X1 U6541 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .IN3(DFF_175_n1), .Q(
        n3128) );
  NOR2X0 U6542 ( .IN1(n4567), .IN2(n3133), .QN(WX1286) );
  XNOR3X1 U6543 ( .IN1(WX877), .IN2(CRC_OUT_9_31), .IN3(DFF_170_n1), .Q(n3133)
         );
  NOR2X0 U6544 ( .IN1(n4567), .IN2(n3140), .QN(WX1272) );
  XNOR3X1 U6545 ( .IN1(WX891), .IN2(CRC_OUT_9_31), .IN3(DFF_163_n1), .Q(n3140)
         );
  NOR2X0 U6546 ( .IN1(n3196), .IN2(n4530), .QN(WX11608) );
  XNOR2X1 U6547 ( .IN1(WX11243), .IN2(DFF_1727_n1), .Q(n3196) );
  NOR2X0 U6548 ( .IN1(n3329), .IN2(n4548), .QN(WX10315) );
  XNOR2X1 U6549 ( .IN1(WX9950), .IN2(DFF_1535_n1), .Q(n3329) );
  NOR2X0 U6550 ( .IN1(n2280), .IN2(n4552), .QN(WX9022) );
  XNOR2X1 U6551 ( .IN1(WX8657), .IN2(DFF_1343_n1), .Q(n2280) );
  NOR2X0 U6552 ( .IN1(n2408), .IN2(n4542), .QN(WX7729) );
  XNOR2X1 U6553 ( .IN1(WX7364), .IN2(DFF_1151_n1), .Q(n2408) );
  NOR2X0 U6554 ( .IN1(n2632), .IN2(n4545), .QN(WX6436) );
  XNOR2X1 U6555 ( .IN1(WX6071), .IN2(DFF_959_n1), .Q(n2632) );
  NOR2X0 U6556 ( .IN1(n2760), .IN2(n4553), .QN(WX5143) );
  XNOR2X1 U6557 ( .IN1(WX4778), .IN2(DFF_767_n1), .Q(n2760) );
  NOR2X0 U6558 ( .IN1(n2888), .IN2(n4538), .QN(WX3850) );
  XNOR2X1 U6559 ( .IN1(WX3485), .IN2(DFF_575_n1), .Q(n2888) );
  NOR2X0 U6560 ( .IN1(n3016), .IN2(n4542), .QN(WX2557) );
  XNOR2X1 U6561 ( .IN1(WX2192), .IN2(DFF_383_n1), .Q(n3016) );
  NOR2X0 U6562 ( .IN1(n3144), .IN2(n4533), .QN(WX1264) );
  XNOR2X1 U6563 ( .IN1(WX899), .IN2(DFF_191_n1), .Q(n3144) );
  NOR2X0 U6564 ( .IN1(n3163), .IN2(n4533), .QN(WX11670) );
  XNOR2X1 U6565 ( .IN1(DFF_1726_n1), .IN2(WX11181), .Q(n3163) );
  NOR2X0 U6566 ( .IN1(n3164), .IN2(n4533), .QN(WX11668) );
  XNOR2X1 U6567 ( .IN1(DFF_1725_n1), .IN2(WX11183), .Q(n3164) );
  NOR2X0 U6568 ( .IN1(n3165), .IN2(n4533), .QN(WX11666) );
  XNOR2X1 U6569 ( .IN1(DFF_1724_n1), .IN2(WX11185), .Q(n3165) );
  NOR2X0 U6570 ( .IN1(n3166), .IN2(n4533), .QN(WX11664) );
  XNOR2X1 U6571 ( .IN1(DFF_1723_n1), .IN2(WX11187), .Q(n3166) );
  NOR2X0 U6572 ( .IN1(n3167), .IN2(n4532), .QN(WX11662) );
  XNOR2X1 U6573 ( .IN1(DFF_1722_n1), .IN2(WX11189), .Q(n3167) );
  NOR2X0 U6574 ( .IN1(n3168), .IN2(n4532), .QN(WX11660) );
  XNOR2X1 U6575 ( .IN1(DFF_1721_n1), .IN2(WX11191), .Q(n3168) );
  NOR2X0 U6576 ( .IN1(n3169), .IN2(n4532), .QN(WX11658) );
  XNOR2X1 U6577 ( .IN1(DFF_1720_n1), .IN2(WX11193), .Q(n3169) );
  NOR2X0 U6578 ( .IN1(n3170), .IN2(n4532), .QN(WX11656) );
  XNOR2X1 U6579 ( .IN1(DFF_1719_n1), .IN2(WX11195), .Q(n3170) );
  NOR2X0 U6580 ( .IN1(n3171), .IN2(n4532), .QN(WX11654) );
  XNOR2X1 U6581 ( .IN1(DFF_1718_n1), .IN2(WX11197), .Q(n3171) );
  NOR2X0 U6582 ( .IN1(n3172), .IN2(n4532), .QN(WX11652) );
  XNOR2X1 U6583 ( .IN1(DFF_1717_n1), .IN2(WX11199), .Q(n3172) );
  NOR2X0 U6584 ( .IN1(n3173), .IN2(n4532), .QN(WX11650) );
  XNOR2X1 U6585 ( .IN1(DFF_1716_n1), .IN2(WX11201), .Q(n3173) );
  NOR2X0 U6586 ( .IN1(n3174), .IN2(n4532), .QN(WX11648) );
  XNOR2X1 U6587 ( .IN1(DFF_1715_n1), .IN2(WX11203), .Q(n3174) );
  NOR2X0 U6588 ( .IN1(n3175), .IN2(n4532), .QN(WX11646) );
  XNOR2X1 U6589 ( .IN1(DFF_1714_n1), .IN2(test_so97), .Q(n3175) );
  NOR2X0 U6590 ( .IN1(n3176), .IN2(n4532), .QN(WX11644) );
  XNOR2X1 U6591 ( .IN1(DFF_1713_n1), .IN2(WX11207), .Q(n3176) );
  NOR2X0 U6592 ( .IN1(n3177), .IN2(n4531), .QN(WX11642) );
  XNOR2X1 U6593 ( .IN1(DFF_1712_n1), .IN2(WX11209), .Q(n3177) );
  NOR2X0 U6594 ( .IN1(n3181), .IN2(n4531), .QN(WX11638) );
  XNOR2X1 U6595 ( .IN1(DFF_1710_n1), .IN2(WX11213), .Q(n3181) );
  NOR2X0 U6596 ( .IN1(n3182), .IN2(n4531), .QN(WX11636) );
  XNOR2X1 U6597 ( .IN1(DFF_1709_n1), .IN2(WX11215), .Q(n3182) );
  NOR2X0 U6598 ( .IN1(n3183), .IN2(n4531), .QN(WX11634) );
  XNOR2X1 U6599 ( .IN1(DFF_1708_n1), .IN2(WX11217), .Q(n3183) );
  NOR2X0 U6600 ( .IN1(n3184), .IN2(n4531), .QN(WX11632) );
  XNOR2X1 U6601 ( .IN1(DFF_1707_n1), .IN2(WX11219), .Q(n3184) );
  NOR2X0 U6602 ( .IN1(n3186), .IN2(n4531), .QN(WX11628) );
  XNOR2X1 U6603 ( .IN1(DFF_1705_n1), .IN2(WX11223), .Q(n3186) );
  NOR2X0 U6604 ( .IN1(n3187), .IN2(n4531), .QN(WX11626) );
  XNOR2X1 U6605 ( .IN1(DFF_1704_n1), .IN2(WX11225), .Q(n3187) );
  NOR2X0 U6606 ( .IN1(n3188), .IN2(n4531), .QN(WX11624) );
  XNOR2X1 U6607 ( .IN1(DFF_1703_n1), .IN2(WX11227), .Q(n3188) );
  NOR2X0 U6608 ( .IN1(n3189), .IN2(n4531), .QN(WX11622) );
  XNOR2X1 U6609 ( .IN1(DFF_1702_n1), .IN2(WX11229), .Q(n3189) );
  NOR2X0 U6610 ( .IN1(n3190), .IN2(n4531), .QN(WX11620) );
  XNOR2X1 U6611 ( .IN1(DFF_1701_n1), .IN2(WX11231), .Q(n3190) );
  NOR2X0 U6612 ( .IN1(n3191), .IN2(n4530), .QN(WX11618) );
  XNOR2X1 U6613 ( .IN1(DFF_1700_n1), .IN2(WX11233), .Q(n3191) );
  NOR2X0 U6614 ( .IN1(n3193), .IN2(n4530), .QN(WX11614) );
  XNOR2X1 U6615 ( .IN1(DFF_1698_n1), .IN2(WX11237), .Q(n3193) );
  NOR2X0 U6616 ( .IN1(n3194), .IN2(n4530), .QN(WX11612) );
  XNOR2X1 U6617 ( .IN1(DFF_1697_n1), .IN2(test_so98), .Q(n3194) );
  NOR2X0 U6618 ( .IN1(n3195), .IN2(n4530), .QN(WX11610) );
  XNOR2X1 U6619 ( .IN1(DFF_1696_n1), .IN2(WX11241), .Q(n3195) );
  NOR2X0 U6620 ( .IN1(n3298), .IN2(n4548), .QN(WX10377) );
  XNOR2X1 U6621 ( .IN1(DFF_1534_n1), .IN2(test_so85), .Q(n3298) );
  NOR2X0 U6622 ( .IN1(n3299), .IN2(n4548), .QN(WX10375) );
  XNOR2X1 U6623 ( .IN1(DFF_1533_n1), .IN2(WX9890), .Q(n3299) );
  NOR2X0 U6624 ( .IN1(n3300), .IN2(n4548), .QN(WX10373) );
  XNOR2X1 U6625 ( .IN1(DFF_1532_n1), .IN2(WX9892), .Q(n3300) );
  NOR2X0 U6626 ( .IN1(n3301), .IN2(n4548), .QN(WX10371) );
  XNOR2X1 U6627 ( .IN1(DFF_1531_n1), .IN2(WX9894), .Q(n3301) );
  NOR2X0 U6628 ( .IN1(n3302), .IN2(n4548), .QN(WX10369) );
  XNOR2X1 U6629 ( .IN1(DFF_1530_n1), .IN2(WX9896), .Q(n3302) );
  NOR2X0 U6630 ( .IN1(n3303), .IN2(n4548), .QN(WX10367) );
  XNOR2X1 U6631 ( .IN1(DFF_1529_n1), .IN2(WX9898), .Q(n3303) );
  NOR2X0 U6632 ( .IN1(n3304), .IN2(n4549), .QN(WX10365) );
  XNOR2X1 U6633 ( .IN1(DFF_1528_n1), .IN2(WX9900), .Q(n3304) );
  NOR2X0 U6634 ( .IN1(n3305), .IN2(n4549), .QN(WX10363) );
  XNOR2X1 U6635 ( .IN1(DFF_1527_n1), .IN2(WX9902), .Q(n3305) );
  NOR2X0 U6636 ( .IN1(n3306), .IN2(n4549), .QN(WX10361) );
  XNOR2X1 U6637 ( .IN1(DFF_1526_n1), .IN2(WX9904), .Q(n3306) );
  NOR2X0 U6638 ( .IN1(n3307), .IN2(n4549), .QN(WX10359) );
  XNOR2X1 U6639 ( .IN1(DFF_1525_n1), .IN2(WX9906), .Q(n3307) );
  NOR2X0 U6640 ( .IN1(n3308), .IN2(n4549), .QN(WX10357) );
  XNOR2X1 U6641 ( .IN1(DFF_1524_n1), .IN2(WX9908), .Q(n3308) );
  NOR2X0 U6642 ( .IN1(n3309), .IN2(n4549), .QN(WX10355) );
  XNOR2X1 U6643 ( .IN1(DFF_1523_n1), .IN2(WX9910), .Q(n3309) );
  NOR2X0 U6644 ( .IN1(n3310), .IN2(n4549), .QN(WX10353) );
  XNOR2X1 U6645 ( .IN1(DFF_1522_n1), .IN2(WX9912), .Q(n3310) );
  NOR2X0 U6646 ( .IN1(n3311), .IN2(n4552), .QN(WX10351) );
  XNOR2X1 U6647 ( .IN1(DFF_1521_n1), .IN2(WX9914), .Q(n3311) );
  NOR2X0 U6648 ( .IN1(n3312), .IN2(n4552), .QN(WX10349) );
  XNOR2X1 U6649 ( .IN1(DFF_1520_n1), .IN2(WX9916), .Q(n3312) );
  NOR2X0 U6650 ( .IN1(n3314), .IN2(n4553), .QN(WX10345) );
  XNOR2X1 U6651 ( .IN1(DFF_1518_n1), .IN2(WX9920), .Q(n3314) );
  NOR2X0 U6652 ( .IN1(n3315), .IN2(n4553), .QN(WX10343) );
  XNOR2X1 U6653 ( .IN1(DFF_1517_n1), .IN2(test_so86), .Q(n3315) );
  NOR2X0 U6654 ( .IN1(n3316), .IN2(n4553), .QN(WX10341) );
  XNOR2X1 U6655 ( .IN1(DFF_1516_n1), .IN2(WX9924), .Q(n3316) );
  NOR2X0 U6656 ( .IN1(n3317), .IN2(n4553), .QN(WX10339) );
  XNOR2X1 U6657 ( .IN1(DFF_1515_n1), .IN2(WX9926), .Q(n3317) );
  NOR2X0 U6658 ( .IN1(n3319), .IN2(n4553), .QN(WX10335) );
  XNOR2X1 U6659 ( .IN1(DFF_1513_n1), .IN2(WX9930), .Q(n3319) );
  NOR2X0 U6660 ( .IN1(n3320), .IN2(n4554), .QN(WX10333) );
  XNOR2X1 U6661 ( .IN1(DFF_1512_n1), .IN2(WX9932), .Q(n3320) );
  NOR2X0 U6662 ( .IN1(n3321), .IN2(n4555), .QN(WX10331) );
  XNOR2X1 U6663 ( .IN1(DFF_1511_n1), .IN2(WX9934), .Q(n3321) );
  NOR2X0 U6664 ( .IN1(n3322), .IN2(n4555), .QN(WX10329) );
  XNOR2X1 U6665 ( .IN1(DFF_1510_n1), .IN2(WX9936), .Q(n3322) );
  NOR2X0 U6666 ( .IN1(n3323), .IN2(n4554), .QN(WX10327) );
  XNOR2X1 U6667 ( .IN1(DFF_1509_n1), .IN2(WX9938), .Q(n3323) );
  NOR2X0 U6668 ( .IN1(n3324), .IN2(n4555), .QN(WX10325) );
  XNOR2X1 U6669 ( .IN1(DFF_1508_n1), .IN2(WX9940), .Q(n3324) );
  NOR2X0 U6670 ( .IN1(n3326), .IN2(n4552), .QN(WX10321) );
  XNOR2X1 U6671 ( .IN1(DFF_1506_n1), .IN2(WX9944), .Q(n3326) );
  NOR2X0 U6672 ( .IN1(n3327), .IN2(n4555), .QN(WX10319) );
  XNOR2X1 U6673 ( .IN1(DFF_1505_n1), .IN2(WX9946), .Q(n3327) );
  NOR2X0 U6674 ( .IN1(n3328), .IN2(n4555), .QN(WX10317) );
  XNOR2X1 U6675 ( .IN1(DFF_1504_n1), .IN2(WX9948), .Q(n3328) );
  NOR2X0 U6676 ( .IN1(n2249), .IN2(n4549), .QN(WX9084) );
  XNOR2X1 U6677 ( .IN1(DFF_1342_n1), .IN2(WX8595), .Q(n2249) );
  NOR2X0 U6678 ( .IN1(n2250), .IN2(n4549), .QN(WX9082) );
  XNOR2X1 U6679 ( .IN1(DFF_1341_n1), .IN2(WX8597), .Q(n2250) );
  NOR2X0 U6680 ( .IN1(n2251), .IN2(n4549), .QN(WX9080) );
  XNOR2X1 U6681 ( .IN1(DFF_1340_n1), .IN2(WX8599), .Q(n2251) );
  NOR2X0 U6682 ( .IN1(n2252), .IN2(n4550), .QN(WX9078) );
  XNOR2X1 U6683 ( .IN1(DFF_1339_n1), .IN2(WX8601), .Q(n2252) );
  NOR2X0 U6684 ( .IN1(n2253), .IN2(n4550), .QN(WX9076) );
  XNOR2X1 U6685 ( .IN1(DFF_1338_n1), .IN2(WX8603), .Q(n2253) );
  NOR2X0 U6686 ( .IN1(n2254), .IN2(n4550), .QN(WX9074) );
  XNOR2X1 U6687 ( .IN1(DFF_1337_n1), .IN2(test_so74), .Q(n2254) );
  NOR2X0 U6688 ( .IN1(n2255), .IN2(n4550), .QN(WX9072) );
  XNOR2X1 U6689 ( .IN1(DFF_1336_n1), .IN2(WX8607), .Q(n2255) );
  NOR2X0 U6690 ( .IN1(n2256), .IN2(n4550), .QN(WX9070) );
  XNOR2X1 U6691 ( .IN1(DFF_1335_n1), .IN2(WX8609), .Q(n2256) );
  NOR2X0 U6692 ( .IN1(n2257), .IN2(n4550), .QN(WX9068) );
  XNOR2X1 U6693 ( .IN1(DFF_1334_n1), .IN2(WX8611), .Q(n2257) );
  NOR2X0 U6694 ( .IN1(n2258), .IN2(n4550), .QN(WX9066) );
  XNOR2X1 U6695 ( .IN1(DFF_1333_n1), .IN2(WX8613), .Q(n2258) );
  NOR2X0 U6696 ( .IN1(n2259), .IN2(n4550), .QN(WX9064) );
  XNOR2X1 U6697 ( .IN1(DFF_1332_n1), .IN2(WX8615), .Q(n2259) );
  NOR2X0 U6698 ( .IN1(n2260), .IN2(n4550), .QN(WX9062) );
  XNOR2X1 U6699 ( .IN1(DFF_1331_n1), .IN2(WX8617), .Q(n2260) );
  NOR2X0 U6700 ( .IN1(n2261), .IN2(n4550), .QN(WX9060) );
  XNOR2X1 U6701 ( .IN1(DFF_1330_n1), .IN2(WX8619), .Q(n2261) );
  NOR2X0 U6702 ( .IN1(n2262), .IN2(n4551), .QN(WX9058) );
  XNOR2X1 U6703 ( .IN1(DFF_1329_n1), .IN2(WX8621), .Q(n2262) );
  NOR2X0 U6704 ( .IN1(n2263), .IN2(n4551), .QN(WX9056) );
  XNOR2X1 U6705 ( .IN1(DFF_1328_n1), .IN2(WX8623), .Q(n2263) );
  NOR2X0 U6706 ( .IN1(n2265), .IN2(n4551), .QN(WX9052) );
  XNOR2X1 U6707 ( .IN1(DFF_1326_n1), .IN2(WX8627), .Q(n2265) );
  NOR2X0 U6708 ( .IN1(n2266), .IN2(n4551), .QN(WX9050) );
  XNOR2X1 U6709 ( .IN1(DFF_1325_n1), .IN2(WX8629), .Q(n2266) );
  NOR2X0 U6710 ( .IN1(n2267), .IN2(n4551), .QN(WX9048) );
  XNOR2X1 U6711 ( .IN1(DFF_1324_n1), .IN2(WX8631), .Q(n2267) );
  NOR2X0 U6712 ( .IN1(n2268), .IN2(n4551), .QN(WX9046) );
  XNOR2X1 U6713 ( .IN1(DFF_1323_n1), .IN2(WX8633), .Q(n2268) );
  NOR2X0 U6714 ( .IN1(n2270), .IN2(n4551), .QN(WX9042) );
  XNOR2X1 U6715 ( .IN1(DFF_1321_n1), .IN2(WX8637), .Q(n2270) );
  NOR2X0 U6716 ( .IN1(n2271), .IN2(n4551), .QN(WX9040) );
  XNOR2X1 U6717 ( .IN1(DFF_1320_n1), .IN2(test_so75), .Q(n2271) );
  NOR2X0 U6718 ( .IN1(n2272), .IN2(n4551), .QN(WX9038) );
  XNOR2X1 U6719 ( .IN1(DFF_1319_n1), .IN2(WX8641), .Q(n2272) );
  NOR2X0 U6720 ( .IN1(n2273), .IN2(n4551), .QN(WX9036) );
  XNOR2X1 U6721 ( .IN1(DFF_1318_n1), .IN2(WX8643), .Q(n2273) );
  NOR2X0 U6722 ( .IN1(n2274), .IN2(n4552), .QN(WX9034) );
  XNOR2X1 U6723 ( .IN1(DFF_1317_n1), .IN2(WX8645), .Q(n2274) );
  NOR2X0 U6724 ( .IN1(n2275), .IN2(n4552), .QN(WX9032) );
  XNOR2X1 U6725 ( .IN1(DFF_1316_n1), .IN2(WX8647), .Q(n2275) );
  NOR2X0 U6726 ( .IN1(n2277), .IN2(n4552), .QN(WX9028) );
  XNOR2X1 U6727 ( .IN1(DFF_1314_n1), .IN2(WX8651), .Q(n2277) );
  NOR2X0 U6728 ( .IN1(n2278), .IN2(n4552), .QN(WX9026) );
  XNOR2X1 U6729 ( .IN1(DFF_1313_n1), .IN2(WX8653), .Q(n2278) );
  NOR2X0 U6730 ( .IN1(n2279), .IN2(n4552), .QN(WX9024) );
  XNOR2X1 U6731 ( .IN1(DFF_1312_n1), .IN2(WX8655), .Q(n2279) );
  NOR2X0 U6732 ( .IN1(n2377), .IN2(n4539), .QN(WX7791) );
  XNOR2X1 U6733 ( .IN1(DFF_1150_n1), .IN2(WX7302), .Q(n2377) );
  NOR2X0 U6734 ( .IN1(n2378), .IN2(n4539), .QN(WX7789) );
  XNOR2X1 U6735 ( .IN1(DFF_1149_n1), .IN2(WX7304), .Q(n2378) );
  NOR2X0 U6736 ( .IN1(n2379), .IN2(n4539), .QN(WX7787) );
  XNOR2X1 U6737 ( .IN1(DFF_1148_n1), .IN2(WX7306), .Q(n2379) );
  NOR2X0 U6738 ( .IN1(n2380), .IN2(n4539), .QN(WX7785) );
  XNOR2X1 U6739 ( .IN1(DFF_1147_n1), .IN2(WX7308), .Q(n2380) );
  NOR2X0 U6740 ( .IN1(n2381), .IN2(n4539), .QN(WX7783) );
  XNOR2X1 U6741 ( .IN1(DFF_1146_n1), .IN2(WX7310), .Q(n2381) );
  NOR2X0 U6742 ( .IN1(n2382), .IN2(n4539), .QN(WX7781) );
  XNOR2X1 U6743 ( .IN1(DFF_1145_n1), .IN2(WX7312), .Q(n2382) );
  NOR2X0 U6744 ( .IN1(n2383), .IN2(n4539), .QN(WX7779) );
  XNOR2X1 U6745 ( .IN1(DFF_1144_n1), .IN2(WX7314), .Q(n2383) );
  NOR2X0 U6746 ( .IN1(n2384), .IN2(n4539), .QN(WX7777) );
  XNOR2X1 U6747 ( .IN1(DFF_1143_n1), .IN2(WX7316), .Q(n2384) );
  NOR2X0 U6748 ( .IN1(n2385), .IN2(n4540), .QN(WX7775) );
  XNOR2X1 U6749 ( .IN1(DFF_1142_n1), .IN2(WX7318), .Q(n2385) );
  NOR2X0 U6750 ( .IN1(n2386), .IN2(n4540), .QN(WX7773) );
  XNOR2X1 U6751 ( .IN1(DFF_1141_n1), .IN2(WX7320), .Q(n2386) );
  NOR2X0 U6752 ( .IN1(n2387), .IN2(n4540), .QN(WX7771) );
  XNOR2X1 U6753 ( .IN1(DFF_1140_n1), .IN2(test_so63), .Q(n2387) );
  NOR2X0 U6754 ( .IN1(n2388), .IN2(n4540), .QN(WX7769) );
  XNOR2X1 U6755 ( .IN1(DFF_1139_n1), .IN2(WX7324), .Q(n2388) );
  NOR2X0 U6756 ( .IN1(n2389), .IN2(n4540), .QN(WX7767) );
  XNOR2X1 U6757 ( .IN1(DFF_1138_n1), .IN2(WX7326), .Q(n2389) );
  NOR2X0 U6758 ( .IN1(n2390), .IN2(n4540), .QN(WX7765) );
  XNOR2X1 U6759 ( .IN1(DFF_1137_n1), .IN2(WX7328), .Q(n2390) );
  NOR2X0 U6760 ( .IN1(n2391), .IN2(n4540), .QN(WX7763) );
  XNOR2X1 U6761 ( .IN1(DFF_1136_n1), .IN2(WX7330), .Q(n2391) );
  NOR2X0 U6762 ( .IN1(n2393), .IN2(n4540), .QN(WX7759) );
  XNOR2X1 U6763 ( .IN1(DFF_1134_n1), .IN2(WX7334), .Q(n2393) );
  NOR2X0 U6764 ( .IN1(n2394), .IN2(n4540), .QN(WX7757) );
  XNOR2X1 U6765 ( .IN1(DFF_1133_n1), .IN2(WX7336), .Q(n2394) );
  NOR2X0 U6766 ( .IN1(n2395), .IN2(n4540), .QN(WX7755) );
  XNOR2X1 U6767 ( .IN1(DFF_1132_n1), .IN2(WX7338), .Q(n2395) );
  NOR2X0 U6768 ( .IN1(n2396), .IN2(n4541), .QN(WX7753) );
  XNOR2X1 U6769 ( .IN1(DFF_1131_n1), .IN2(WX7340), .Q(n2396) );
  NOR2X0 U6770 ( .IN1(n2398), .IN2(n4541), .QN(WX7749) );
  XNOR2X1 U6771 ( .IN1(DFF_1129_n1), .IN2(WX7344), .Q(n2398) );
  NOR2X0 U6772 ( .IN1(n2399), .IN2(n4541), .QN(WX7747) );
  XNOR2X1 U6773 ( .IN1(DFF_1128_n1), .IN2(WX7346), .Q(n2399) );
  NOR2X0 U6774 ( .IN1(n2400), .IN2(n4541), .QN(WX7745) );
  XNOR2X1 U6775 ( .IN1(DFF_1127_n1), .IN2(WX7348), .Q(n2400) );
  NOR2X0 U6776 ( .IN1(n2401), .IN2(n4541), .QN(WX7743) );
  XNOR2X1 U6777 ( .IN1(DFF_1126_n1), .IN2(WX7350), .Q(n2401) );
  NOR2X0 U6778 ( .IN1(n2402), .IN2(n4541), .QN(WX7741) );
  XNOR2X1 U6779 ( .IN1(DFF_1125_n1), .IN2(WX7352), .Q(n2402) );
  NOR2X0 U6780 ( .IN1(n2403), .IN2(n4541), .QN(WX7739) );
  XNOR2X1 U6781 ( .IN1(DFF_1124_n1), .IN2(WX7354), .Q(n2403) );
  NOR2X0 U6782 ( .IN1(n2405), .IN2(n4541), .QN(WX7735) );
  XNOR2X1 U6783 ( .IN1(DFF_1122_n1), .IN2(WX7358), .Q(n2405) );
  NOR2X0 U6784 ( .IN1(n2406), .IN2(n4541), .QN(WX7733) );
  XNOR2X1 U6785 ( .IN1(DFF_1121_n1), .IN2(WX7360), .Q(n2406) );
  NOR2X0 U6786 ( .IN1(n2407), .IN2(n4541), .QN(WX7731) );
  XNOR2X1 U6787 ( .IN1(DFF_1120_n1), .IN2(WX7362), .Q(n2407) );
  NOR2X0 U6788 ( .IN1(n2592), .IN2(n4546), .QN(WX6498) );
  XNOR2X1 U6789 ( .IN1(DFF_958_n1), .IN2(WX6009), .Q(n2592) );
  NOR2X0 U6790 ( .IN1(n2593), .IN2(n4546), .QN(WX6496) );
  XNOR2X1 U6791 ( .IN1(DFF_957_n1), .IN2(WX6011), .Q(n2593) );
  NOR2X0 U6792 ( .IN1(n2594), .IN2(n4546), .QN(WX6494) );
  XNOR2X1 U6793 ( .IN1(DFF_956_n1), .IN2(WX6013), .Q(n2594) );
  NOR2X0 U6794 ( .IN1(n2595), .IN2(n4546), .QN(WX6492) );
  XNOR2X1 U6795 ( .IN1(DFF_955_n1), .IN2(WX6015), .Q(n2595) );
  NOR2X0 U6796 ( .IN1(n2596), .IN2(n4546), .QN(WX6490) );
  XNOR2X1 U6797 ( .IN1(DFF_954_n1), .IN2(WX6017), .Q(n2596) );
  NOR2X0 U6798 ( .IN1(n2597), .IN2(n4546), .QN(WX6488) );
  XNOR2X1 U6799 ( .IN1(DFF_953_n1), .IN2(WX6019), .Q(n2597) );
  NOR2X0 U6800 ( .IN1(n2598), .IN2(n4546), .QN(WX6486) );
  XNOR2X1 U6801 ( .IN1(DFF_952_n1), .IN2(WX6021), .Q(n2598) );
  NOR2X0 U6802 ( .IN1(n2599), .IN2(n4546), .QN(WX6484) );
  XNOR2X1 U6803 ( .IN1(DFF_951_n1), .IN2(WX6023), .Q(n2599) );
  NOR2X0 U6804 ( .IN1(n2600), .IN2(n4547), .QN(WX6482) );
  XNOR2X1 U6805 ( .IN1(DFF_950_n1), .IN2(WX6025), .Q(n2600) );
  NOR2X0 U6806 ( .IN1(n2601), .IN2(n4547), .QN(WX6480) );
  XNOR2X1 U6807 ( .IN1(DFF_949_n1), .IN2(WX6027), .Q(n2601) );
  NOR2X0 U6808 ( .IN1(n2605), .IN2(n4547), .QN(WX6478) );
  XNOR2X1 U6809 ( .IN1(DFF_948_n1), .IN2(WX6029), .Q(n2605) );
  NOR2X0 U6810 ( .IN1(n2606), .IN2(n4547), .QN(WX6476) );
  XNOR2X1 U6811 ( .IN1(DFF_947_n1), .IN2(WX6031), .Q(n2606) );
  NOR2X0 U6812 ( .IN1(n2607), .IN2(n4547), .QN(WX6474) );
  XNOR2X1 U6813 ( .IN1(DFF_946_n1), .IN2(WX6033), .Q(n2607) );
  NOR2X0 U6814 ( .IN1(n2608), .IN2(n4547), .QN(WX6472) );
  XNOR2X1 U6815 ( .IN1(DFF_945_n1), .IN2(WX6035), .Q(n2608) );
  NOR2X0 U6816 ( .IN1(n2609), .IN2(n4547), .QN(WX6470) );
  XNOR2X1 U6817 ( .IN1(DFF_944_n1), .IN2(WX6037), .Q(n2609) );
  NOR2X0 U6818 ( .IN1(n2611), .IN2(n4547), .QN(WX6466) );
  XNOR2X1 U6819 ( .IN1(DFF_942_n1), .IN2(WX6041), .Q(n2611) );
  NOR2X0 U6820 ( .IN1(n2612), .IN2(n4547), .QN(WX6464) );
  XNOR2X1 U6821 ( .IN1(DFF_941_n1), .IN2(WX6043), .Q(n2612) );
  NOR2X0 U6822 ( .IN1(n2613), .IN2(n4547), .QN(WX6462) );
  XNOR2X1 U6823 ( .IN1(DFF_940_n1), .IN2(WX6045), .Q(n2613) );
  NOR2X0 U6824 ( .IN1(n2614), .IN2(n4529), .QN(WX6460) );
  XNOR2X1 U6825 ( .IN1(DFF_939_n1), .IN2(WX6047), .Q(n2614) );
  NOR2X0 U6826 ( .IN1(n2619), .IN2(n4546), .QN(WX6456) );
  XNOR2X1 U6827 ( .IN1(DFF_937_n1), .IN2(WX6051), .Q(n2619) );
  NOR2X0 U6828 ( .IN1(n2620), .IN2(n4545), .QN(WX6454) );
  XNOR2X1 U6829 ( .IN1(DFF_936_n1), .IN2(WX6053), .Q(n2620) );
  NOR2X0 U6830 ( .IN1(n2621), .IN2(n4545), .QN(WX6452) );
  XNOR2X1 U6831 ( .IN1(DFF_935_n1), .IN2(WX6055), .Q(n2621) );
  NOR2X0 U6832 ( .IN1(n2622), .IN2(n4545), .QN(WX6450) );
  XNOR2X1 U6833 ( .IN1(DFF_934_n1), .IN2(WX6057), .Q(n2622) );
  NOR2X0 U6834 ( .IN1(n2623), .IN2(n4545), .QN(WX6448) );
  XNOR2X1 U6835 ( .IN1(DFF_933_n1), .IN2(WX6059), .Q(n2623) );
  NOR2X0 U6836 ( .IN1(n2624), .IN2(n4545), .QN(WX6446) );
  XNOR2X1 U6837 ( .IN1(DFF_932_n1), .IN2(WX6061), .Q(n2624) );
  NOR2X0 U6838 ( .IN1(n2626), .IN2(n4545), .QN(WX6442) );
  XNOR2X1 U6839 ( .IN1(DFF_930_n1), .IN2(WX6065), .Q(n2626) );
  NOR2X0 U6840 ( .IN1(n2627), .IN2(n4545), .QN(WX6440) );
  XNOR2X1 U6841 ( .IN1(DFF_929_n1), .IN2(WX6067), .Q(n2627) );
  NOR2X0 U6842 ( .IN1(n2631), .IN2(n4545), .QN(WX6438) );
  XNOR2X1 U6843 ( .IN1(DFF_928_n1), .IN2(WX6069), .Q(n2631) );
  NOR2X0 U6844 ( .IN1(n2729), .IN2(n4529), .QN(WX5205) );
  XNOR2X1 U6845 ( .IN1(DFF_766_n1), .IN2(WX4716), .Q(n2729) );
  NOR2X0 U6846 ( .IN1(n2730), .IN2(n4529), .QN(WX5203) );
  XNOR2X1 U6847 ( .IN1(DFF_765_n1), .IN2(WX4718), .Q(n2730) );
  NOR2X0 U6848 ( .IN1(n2731), .IN2(n4529), .QN(WX5201) );
  XNOR2X1 U6849 ( .IN1(DFF_764_n1), .IN2(WX4720), .Q(n2731) );
  NOR2X0 U6850 ( .IN1(n2732), .IN2(n4529), .QN(WX5199) );
  XNOR2X1 U6851 ( .IN1(DFF_763_n1), .IN2(test_so40), .Q(n2732) );
  NOR2X0 U6852 ( .IN1(n2733), .IN2(n4529), .QN(WX5197) );
  XNOR2X1 U6853 ( .IN1(DFF_762_n1), .IN2(WX4724), .Q(n2733) );
  NOR2X0 U6854 ( .IN1(n2734), .IN2(n4529), .QN(WX5195) );
  XNOR2X1 U6855 ( .IN1(DFF_761_n1), .IN2(WX4726), .Q(n2734) );
  NOR2X0 U6856 ( .IN1(n2735), .IN2(n4529), .QN(WX5193) );
  XNOR2X1 U6857 ( .IN1(DFF_760_n1), .IN2(WX4728), .Q(n2735) );
  NOR2X0 U6858 ( .IN1(n2736), .IN2(n4529), .QN(WX5191) );
  XNOR2X1 U6859 ( .IN1(DFF_759_n1), .IN2(WX4730), .Q(n2736) );
  NOR2X0 U6860 ( .IN1(n2737), .IN2(n4529), .QN(WX5189) );
  XNOR2X1 U6861 ( .IN1(DFF_758_n1), .IN2(WX4732), .Q(n2737) );
  NOR2X0 U6862 ( .IN1(n2738), .IN2(n4538), .QN(WX5187) );
  XNOR2X1 U6863 ( .IN1(DFF_757_n1), .IN2(WX4734), .Q(n2738) );
  NOR2X0 U6864 ( .IN1(n2739), .IN2(n4554), .QN(WX5185) );
  XNOR2X1 U6865 ( .IN1(DFF_756_n1), .IN2(WX4736), .Q(n2739) );
  NOR2X0 U6866 ( .IN1(n2740), .IN2(n4555), .QN(WX5183) );
  XNOR2X1 U6867 ( .IN1(DFF_755_n1), .IN2(WX4738), .Q(n2740) );
  NOR2X0 U6868 ( .IN1(n2741), .IN2(n4555), .QN(WX5181) );
  XNOR2X1 U6869 ( .IN1(DFF_754_n1), .IN2(WX4740), .Q(n2741) );
  NOR2X0 U6870 ( .IN1(n2742), .IN2(n4555), .QN(WX5179) );
  XNOR2X1 U6871 ( .IN1(DFF_753_n1), .IN2(WX4742), .Q(n2742) );
  NOR2X0 U6872 ( .IN1(n2743), .IN2(n4555), .QN(WX5177) );
  XNOR2X1 U6873 ( .IN1(DFF_752_n1), .IN2(WX4744), .Q(n2743) );
  NOR2X0 U6874 ( .IN1(n2745), .IN2(n4555), .QN(WX5173) );
  XNOR2X1 U6875 ( .IN1(DFF_750_n1), .IN2(WX4748), .Q(n2745) );
  NOR2X0 U6876 ( .IN1(n2746), .IN2(n4554), .QN(WX5171) );
  XNOR2X1 U6877 ( .IN1(DFF_749_n1), .IN2(WX4750), .Q(n2746) );
  NOR2X0 U6878 ( .IN1(n2747), .IN2(n4554), .QN(WX5169) );
  XNOR2X1 U6879 ( .IN1(DFF_748_n1), .IN2(WX4752), .Q(n2747) );
  NOR2X0 U6880 ( .IN1(n2748), .IN2(n4554), .QN(WX5167) );
  XNOR2X1 U6881 ( .IN1(DFF_747_n1), .IN2(WX4754), .Q(n2748) );
  NOR2X0 U6882 ( .IN1(n2750), .IN2(n4554), .QN(WX5163) );
  XNOR2X1 U6883 ( .IN1(DFF_745_n1), .IN2(WX4758), .Q(n2750) );
  NOR2X0 U6884 ( .IN1(n2751), .IN2(n4552), .QN(WX5161) );
  XNOR2X1 U6885 ( .IN1(DFF_744_n1), .IN2(WX4760), .Q(n2751) );
  NOR2X0 U6886 ( .IN1(n2752), .IN2(n4554), .QN(WX5159) );
  XNOR2X1 U6887 ( .IN1(DFF_743_n1), .IN2(WX4762), .Q(n2752) );
  NOR2X0 U6888 ( .IN1(n2753), .IN2(n4554), .QN(WX5157) );
  XNOR2X1 U6889 ( .IN1(DFF_742_n1), .IN2(WX4764), .Q(n2753) );
  NOR2X0 U6890 ( .IN1(n2754), .IN2(n4553), .QN(WX5155) );
  XNOR2X1 U6891 ( .IN1(DFF_741_n1), .IN2(WX4766), .Q(n2754) );
  NOR2X0 U6892 ( .IN1(n2755), .IN2(n4554), .QN(WX5153) );
  XNOR2X1 U6893 ( .IN1(DFF_740_n1), .IN2(WX4768), .Q(n2755) );
  NOR2X0 U6894 ( .IN1(n2757), .IN2(n4553), .QN(WX5149) );
  XNOR2X1 U6895 ( .IN1(DFF_738_n1), .IN2(WX4772), .Q(n2757) );
  NOR2X0 U6896 ( .IN1(n2758), .IN2(n4553), .QN(WX5147) );
  XNOR2X1 U6897 ( .IN1(DFF_737_n1), .IN2(WX4774), .Q(n2758) );
  NOR2X0 U6898 ( .IN1(n2759), .IN2(n4553), .QN(WX5145) );
  XNOR2X1 U6899 ( .IN1(DFF_736_n1), .IN2(WX4776), .Q(n2759) );
  NOR2X0 U6900 ( .IN1(n2857), .IN2(n4530), .QN(WX3912) );
  XNOR2X1 U6901 ( .IN1(DFF_574_n1), .IN2(WX3423), .Q(n2857) );
  NOR2X0 U6902 ( .IN1(n2858), .IN2(n4530), .QN(WX3910) );
  XNOR2X1 U6903 ( .IN1(DFF_573_n1), .IN2(WX3425), .Q(n2858) );
  NOR2X0 U6904 ( .IN1(n2859), .IN2(n4530), .QN(WX3908) );
  XNOR2X1 U6905 ( .IN1(DFF_572_n1), .IN2(WX3427), .Q(n2859) );
  NOR2X0 U6906 ( .IN1(n2860), .IN2(n4530), .QN(WX3906) );
  XNOR2X1 U6907 ( .IN1(DFF_571_n1), .IN2(WX3429), .Q(n2860) );
  NOR2X0 U6908 ( .IN1(n2861), .IN2(n4530), .QN(WX3904) );
  XNOR2X1 U6909 ( .IN1(DFF_570_n1), .IN2(WX3431), .Q(n2861) );
  NOR2X0 U6910 ( .IN1(n2862), .IN2(n4536), .QN(WX3902) );
  XNOR2X1 U6911 ( .IN1(DFF_569_n1), .IN2(WX3433), .Q(n2862) );
  NOR2X0 U6912 ( .IN1(n2863), .IN2(n4536), .QN(WX3900) );
  XNOR2X1 U6913 ( .IN1(DFF_568_n1), .IN2(WX3435), .Q(n2863) );
  NOR2X0 U6914 ( .IN1(n2864), .IN2(n4536), .QN(WX3898) );
  XNOR2X1 U6915 ( .IN1(DFF_567_n1), .IN2(WX3437), .Q(n2864) );
  NOR2X0 U6916 ( .IN1(n2865), .IN2(n4536), .QN(WX3896) );
  XNOR2X1 U6917 ( .IN1(DFF_566_n1), .IN2(test_so29), .Q(n2865) );
  NOR2X0 U6918 ( .IN1(n2866), .IN2(n4536), .QN(WX3894) );
  XNOR2X1 U6919 ( .IN1(DFF_565_n1), .IN2(WX3441), .Q(n2866) );
  NOR2X0 U6920 ( .IN1(n2867), .IN2(n4537), .QN(WX3892) );
  XNOR2X1 U6921 ( .IN1(DFF_564_n1), .IN2(WX3443), .Q(n2867) );
  NOR2X0 U6922 ( .IN1(n2868), .IN2(n4537), .QN(WX3890) );
  XNOR2X1 U6923 ( .IN1(DFF_563_n1), .IN2(WX3445), .Q(n2868) );
  NOR2X0 U6924 ( .IN1(n2869), .IN2(n4537), .QN(WX3888) );
  XNOR2X1 U6925 ( .IN1(DFF_562_n1), .IN2(WX3447), .Q(n2869) );
  NOR2X0 U6926 ( .IN1(n2870), .IN2(n4537), .QN(WX3886) );
  XNOR2X1 U6927 ( .IN1(DFF_561_n1), .IN2(WX3449), .Q(n2870) );
  NOR2X0 U6928 ( .IN1(n2871), .IN2(n4537), .QN(WX3884) );
  XNOR2X1 U6929 ( .IN1(DFF_560_n1), .IN2(WX3451), .Q(n2871) );
  NOR2X0 U6930 ( .IN1(n2873), .IN2(n4537), .QN(WX3880) );
  XNOR2X1 U6931 ( .IN1(DFF_558_n1), .IN2(WX3455), .Q(n2873) );
  NOR2X0 U6932 ( .IN1(n2874), .IN2(n4537), .QN(WX3878) );
  XNOR2X1 U6933 ( .IN1(DFF_557_n1), .IN2(WX3457), .Q(n2874) );
  NOR2X0 U6934 ( .IN1(n2875), .IN2(n4537), .QN(WX3876) );
  XNOR2X1 U6935 ( .IN1(DFF_556_n1), .IN2(WX3459), .Q(n2875) );
  NOR2X0 U6936 ( .IN1(n2876), .IN2(n4537), .QN(WX3874) );
  XNOR2X1 U6937 ( .IN1(DFF_555_n1), .IN2(WX3461), .Q(n2876) );
  NOR2X0 U6938 ( .IN1(n2878), .IN2(n4537), .QN(WX3870) );
  XNOR2X1 U6939 ( .IN1(DFF_553_n1), .IN2(WX3465), .Q(n2878) );
  NOR2X0 U6940 ( .IN1(n2879), .IN2(n4538), .QN(WX3868) );
  XNOR2X1 U6941 ( .IN1(DFF_552_n1), .IN2(WX3467), .Q(n2879) );
  NOR2X0 U6942 ( .IN1(n2880), .IN2(n4538), .QN(WX3866) );
  XNOR2X1 U6943 ( .IN1(DFF_551_n1), .IN2(WX3469), .Q(n2880) );
  NOR2X0 U6944 ( .IN1(n2881), .IN2(n4538), .QN(WX3864) );
  XNOR2X1 U6945 ( .IN1(DFF_550_n1), .IN2(WX3471), .Q(n2881) );
  NOR2X0 U6946 ( .IN1(n2882), .IN2(n4538), .QN(WX3862) );
  XNOR2X1 U6947 ( .IN1(DFF_549_n1), .IN2(test_so30), .Q(n2882) );
  NOR2X0 U6948 ( .IN1(n2883), .IN2(n4538), .QN(WX3860) );
  XNOR2X1 U6949 ( .IN1(DFF_548_n1), .IN2(WX3475), .Q(n2883) );
  NOR2X0 U6950 ( .IN1(n2885), .IN2(n4538), .QN(WX3856) );
  XNOR2X1 U6951 ( .IN1(DFF_546_n1), .IN2(WX3479), .Q(n2885) );
  NOR2X0 U6952 ( .IN1(n2886), .IN2(n4538), .QN(WX3854) );
  XNOR2X1 U6953 ( .IN1(DFF_545_n1), .IN2(WX3481), .Q(n2886) );
  NOR2X0 U6954 ( .IN1(n2887), .IN2(n4538), .QN(WX3852) );
  XNOR2X1 U6955 ( .IN1(DFF_544_n1), .IN2(WX3483), .Q(n2887) );
  NOR2X0 U6956 ( .IN1(n2985), .IN2(n4544), .QN(WX2619) );
  XNOR2X1 U6957 ( .IN1(DFF_382_n1), .IN2(WX2130), .Q(n2985) );
  NOR2X0 U6958 ( .IN1(n2986), .IN2(n4544), .QN(WX2617) );
  XNOR2X1 U6959 ( .IN1(DFF_381_n1), .IN2(WX2132), .Q(n2986) );
  NOR2X0 U6960 ( .IN1(n2987), .IN2(n4544), .QN(WX2615) );
  XNOR2X1 U6961 ( .IN1(DFF_380_n1), .IN2(WX2134), .Q(n2987) );
  NOR2X0 U6962 ( .IN1(n2988), .IN2(n4544), .QN(WX2613) );
  XNOR2X1 U6963 ( .IN1(DFF_379_n1), .IN2(test_so18), .Q(n2988) );
  NOR2X0 U6964 ( .IN1(n2989), .IN2(n4544), .QN(WX2611) );
  XNOR2X1 U6965 ( .IN1(DFF_378_n1), .IN2(WX2138), .Q(n2989) );
  NOR2X0 U6966 ( .IN1(n2990), .IN2(n4544), .QN(WX2609) );
  XNOR2X1 U6967 ( .IN1(DFF_377_n1), .IN2(WX2140), .Q(n2990) );
  NOR2X0 U6968 ( .IN1(n2991), .IN2(n4544), .QN(WX2607) );
  XNOR2X1 U6969 ( .IN1(DFF_376_n1), .IN2(WX2142), .Q(n2991) );
  NOR2X0 U6970 ( .IN1(n2992), .IN2(n4544), .QN(WX2605) );
  XNOR2X1 U6971 ( .IN1(DFF_375_n1), .IN2(WX2144), .Q(n2992) );
  NOR2X0 U6972 ( .IN1(n2993), .IN2(n4544), .QN(WX2603) );
  XNOR2X1 U6973 ( .IN1(DFF_374_n1), .IN2(WX2146), .Q(n2993) );
  NOR2X0 U6974 ( .IN1(n2994), .IN2(n4544), .QN(WX2601) );
  XNOR2X1 U6975 ( .IN1(DFF_373_n1), .IN2(WX2148), .Q(n2994) );
  NOR2X0 U6976 ( .IN1(n2995), .IN2(n4543), .QN(WX2599) );
  XNOR2X1 U6977 ( .IN1(DFF_372_n1), .IN2(WX2150), .Q(n2995) );
  NOR2X0 U6978 ( .IN1(n2996), .IN2(n4543), .QN(WX2597) );
  XNOR2X1 U6979 ( .IN1(DFF_371_n1), .IN2(WX2152), .Q(n2996) );
  NOR2X0 U6980 ( .IN1(n2997), .IN2(n4543), .QN(WX2595) );
  XNOR2X1 U6981 ( .IN1(DFF_370_n1), .IN2(WX2154), .Q(n2997) );
  NOR2X0 U6982 ( .IN1(n2998), .IN2(n4543), .QN(WX2593) );
  XNOR2X1 U6983 ( .IN1(DFF_369_n1), .IN2(WX2156), .Q(n2998) );
  NOR2X0 U6984 ( .IN1(n2999), .IN2(n4543), .QN(WX2591) );
  XNOR2X1 U6985 ( .IN1(DFF_368_n1), .IN2(WX2158), .Q(n2999) );
  NOR2X0 U6986 ( .IN1(n3001), .IN2(n4543), .QN(WX2587) );
  XNOR2X1 U6987 ( .IN1(DFF_366_n1), .IN2(WX2162), .Q(n3001) );
  NOR2X0 U6988 ( .IN1(n3002), .IN2(n4543), .QN(WX2585) );
  XNOR2X1 U6989 ( .IN1(DFF_365_n1), .IN2(WX2164), .Q(n3002) );
  NOR2X0 U6990 ( .IN1(n3003), .IN2(n4543), .QN(WX2583) );
  XNOR2X1 U6991 ( .IN1(DFF_364_n1), .IN2(WX2166), .Q(n3003) );
  NOR2X0 U6992 ( .IN1(n3004), .IN2(n4543), .QN(WX2581) );
  XNOR2X1 U6993 ( .IN1(DFF_363_n1), .IN2(WX2168), .Q(n3004) );
  NOR2X0 U6994 ( .IN1(n3006), .IN2(n4543), .QN(WX2577) );
  XNOR2X1 U6995 ( .IN1(DFF_361_n1), .IN2(test_so19), .Q(n3006) );
  NOR2X0 U6996 ( .IN1(n3007), .IN2(n4542), .QN(WX2575) );
  XNOR2X1 U6997 ( .IN1(DFF_360_n1), .IN2(WX2174), .Q(n3007) );
  NOR2X0 U6998 ( .IN1(n3008), .IN2(n4542), .QN(WX2573) );
  XNOR2X1 U6999 ( .IN1(DFF_359_n1), .IN2(WX2176), .Q(n3008) );
  NOR2X0 U7000 ( .IN1(n3009), .IN2(n4542), .QN(WX2571) );
  XNOR2X1 U7001 ( .IN1(DFF_358_n1), .IN2(WX2178), .Q(n3009) );
  NOR2X0 U7002 ( .IN1(n3010), .IN2(n4542), .QN(WX2569) );
  XNOR2X1 U7003 ( .IN1(DFF_357_n1), .IN2(WX2180), .Q(n3010) );
  NOR2X0 U7004 ( .IN1(n3011), .IN2(n4542), .QN(WX2567) );
  XNOR2X1 U7005 ( .IN1(DFF_356_n1), .IN2(WX2182), .Q(n3011) );
  NOR2X0 U7006 ( .IN1(n3013), .IN2(n4542), .QN(WX2563) );
  XNOR2X1 U7007 ( .IN1(DFF_354_n1), .IN2(WX2186), .Q(n3013) );
  NOR2X0 U7008 ( .IN1(n3014), .IN2(n4542), .QN(WX2561) );
  XNOR2X1 U7009 ( .IN1(DFF_353_n1), .IN2(WX2188), .Q(n3014) );
  NOR2X0 U7010 ( .IN1(n3015), .IN2(n4542), .QN(WX2559) );
  XNOR2X1 U7011 ( .IN1(DFF_352_n1), .IN2(WX2190), .Q(n3015) );
  NOR2X0 U7012 ( .IN1(n3113), .IN2(n4536), .QN(WX1326) );
  XNOR2X1 U7013 ( .IN1(DFF_190_n1), .IN2(WX837), .Q(n3113) );
  NOR2X0 U7014 ( .IN1(n3114), .IN2(n4536), .QN(WX1324) );
  XNOR2X1 U7015 ( .IN1(DFF_189_n1), .IN2(WX839), .Q(n3114) );
  NOR2X0 U7016 ( .IN1(n3115), .IN2(n4536), .QN(WX1322) );
  XNOR2X1 U7017 ( .IN1(DFF_188_n1), .IN2(WX841), .Q(n3115) );
  NOR2X0 U7018 ( .IN1(n3116), .IN2(n4535), .QN(WX1320) );
  XNOR2X1 U7019 ( .IN1(DFF_187_n1), .IN2(WX843), .Q(n3116) );
  NOR2X0 U7020 ( .IN1(n3117), .IN2(n4535), .QN(WX1318) );
  XNOR2X1 U7021 ( .IN1(DFF_186_n1), .IN2(WX845), .Q(n3117) );
  NOR2X0 U7022 ( .IN1(n3118), .IN2(n4535), .QN(WX1316) );
  XNOR2X1 U7023 ( .IN1(DFF_185_n1), .IN2(WX847), .Q(n3118) );
  NOR2X0 U7024 ( .IN1(n3119), .IN2(n4535), .QN(WX1314) );
  XNOR2X1 U7025 ( .IN1(DFF_184_n1), .IN2(WX849), .Q(n3119) );
  NOR2X0 U7026 ( .IN1(n3120), .IN2(n4535), .QN(WX1312) );
  XNOR2X1 U7027 ( .IN1(DFF_183_n1), .IN2(WX851), .Q(n3120) );
  NOR2X0 U7028 ( .IN1(n3121), .IN2(n4535), .QN(WX1310) );
  XNOR2X1 U7029 ( .IN1(DFF_182_n1), .IN2(WX853), .Q(n3121) );
  NOR2X0 U7030 ( .IN1(n3122), .IN2(n4535), .QN(WX1308) );
  XNOR2X1 U7031 ( .IN1(DFF_181_n1), .IN2(WX855), .Q(n3122) );
  NOR2X0 U7032 ( .IN1(n3123), .IN2(n4535), .QN(WX1306) );
  XNOR2X1 U7033 ( .IN1(DFF_180_n1), .IN2(WX857), .Q(n3123) );
  NOR2X0 U7034 ( .IN1(n3124), .IN2(n4535), .QN(WX1304) );
  XNOR2X1 U7035 ( .IN1(DFF_179_n1), .IN2(WX859), .Q(n3124) );
  NOR2X0 U7036 ( .IN1(n3125), .IN2(n4535), .QN(WX1302) );
  XNOR2X1 U7037 ( .IN1(DFF_178_n1), .IN2(WX861), .Q(n3125) );
  NOR2X0 U7038 ( .IN1(n3126), .IN2(n4534), .QN(WX1300) );
  XNOR2X1 U7039 ( .IN1(DFF_177_n1), .IN2(WX863), .Q(n3126) );
  NOR2X0 U7040 ( .IN1(n3127), .IN2(n4534), .QN(WX1298) );
  XNOR2X1 U7041 ( .IN1(DFF_176_n1), .IN2(WX865), .Q(n3127) );
  NOR2X0 U7042 ( .IN1(n3129), .IN2(n4534), .QN(WX1294) );
  XNOR2X1 U7043 ( .IN1(DFF_174_n1), .IN2(WX869), .Q(n3129) );
  NOR2X0 U7044 ( .IN1(n3130), .IN2(n4534), .QN(WX1292) );
  XNOR2X1 U7045 ( .IN1(DFF_173_n1), .IN2(WX871), .Q(n3130) );
  NOR2X0 U7046 ( .IN1(n3131), .IN2(n4534), .QN(WX1290) );
  XNOR2X1 U7047 ( .IN1(DFF_172_n1), .IN2(WX873), .Q(n3131) );
  NOR2X0 U7048 ( .IN1(n3132), .IN2(n4534), .QN(WX1288) );
  XNOR2X1 U7049 ( .IN1(DFF_171_n1), .IN2(WX875), .Q(n3132) );
  NOR2X0 U7050 ( .IN1(n3134), .IN2(n4534), .QN(WX1284) );
  XNOR2X1 U7051 ( .IN1(DFF_169_n1), .IN2(WX879), .Q(n3134) );
  NOR2X0 U7052 ( .IN1(n3135), .IN2(n4534), .QN(WX1282) );
  XNOR2X1 U7053 ( .IN1(DFF_168_n1), .IN2(WX881), .Q(n3135) );
  NOR2X0 U7054 ( .IN1(n3136), .IN2(n4534), .QN(WX1280) );
  XNOR2X1 U7055 ( .IN1(DFF_167_n1), .IN2(WX883), .Q(n3136) );
  NOR2X0 U7056 ( .IN1(n3137), .IN2(n4534), .QN(WX1278) );
  XNOR2X1 U7057 ( .IN1(DFF_166_n1), .IN2(WX885), .Q(n3137) );
  NOR2X0 U7058 ( .IN1(n3138), .IN2(n4533), .QN(WX1276) );
  XNOR2X1 U7059 ( .IN1(DFF_165_n1), .IN2(WX887), .Q(n3138) );
  NOR2X0 U7060 ( .IN1(n3139), .IN2(n4533), .QN(WX1274) );
  XNOR2X1 U7061 ( .IN1(DFF_164_n1), .IN2(WX889), .Q(n3139) );
  NOR2X0 U7062 ( .IN1(n3141), .IN2(n4533), .QN(WX1270) );
  XNOR2X1 U7063 ( .IN1(DFF_162_n1), .IN2(WX893), .Q(n3141) );
  NOR2X0 U7064 ( .IN1(n3142), .IN2(n4533), .QN(WX1268) );
  XNOR2X1 U7065 ( .IN1(DFF_161_n1), .IN2(WX895), .Q(n3142) );
  NOR2X0 U7066 ( .IN1(n3143), .IN2(n4533), .QN(WX1266) );
  XNOR2X1 U7067 ( .IN1(DFF_160_n1), .IN2(WX897), .Q(n3143) );


  // Trigger -----------------------
  AND2X1 Trojan1 ( .IN1(WX742), .IN2(WX7249), .Q(Tj_OUT1) );
  AND2X1 Trojan2 ( .IN1(WX5922), .IN2(WX5960), .Q(Tj_OUT2) );
  AND2X1 Trojan3 ( .IN1(WX4697), .IN2(WX9032), .Q(Tj_OUT3) );
  AND2X1 Trojan4 ( .IN1(WX8298), .IN2(WX10846), .Q(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT1), .IN3(Tj_OUT3), .IN4(Tj_OUT4), .QN(Tj_OUT1234) );
  AND2X1 Trojan5 ( .IN1(WX3340), .IN2(WX6476), .Q(Tj_OUT5) );
  AND2X1 Trojan6 ( .IN1(WX9819), .IN2(WX1813), .Q(Tj_OUT6) );
  AND2X1 Trojan7 ( .IN1(WX5710), .IN2(WX3458), .Q(Tj_OUT7) );
  AND2X1 Trojan8 ( .IN1(WX9060), .IN2(WX7749), .Q(Tj_OUT8) );
  NOR4X0 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(Tj_OUT8), .QN(Tj_OUT5678) );

  INVX0 TrojanINV_test_se ( .IN(test_se), .QN(test_se_NOT) );  
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  DFFX2 TrojanScanEnable ( .CLK(Tj_Trigger), .D(1'b1), .Q(Trojan_SE) );

  // Payload -----------------------
  MUX21X1 Trojan_Payload1 ( .IN1(test_se), .IN2(1'b1), .S(Trojan_SE), .Q(test_se_Trojan) );
  MUX21X1 Trojan_Payload2 ( .IN1(WX11155), .IN2(WX3442), .S(Trojan_SE), .Q(WX11155_Tj_Payload) );

endmodule
