module top(n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [2:0] n6;
    wire [63:0] n7;
    wire [7:0] n8;
    wire [19:0] n9;
    wire n10, n11, n12, n13, n14, n15, n16, n17;
    wire n18, n19, n20, n21, n22, n23, n24, n25;
    wire n26, n27, n28, n29, n30, n31, n32, n33;
    wire n34, n35, n36, n37, n38, n39, n40, n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    wire n442, n443, n444, n445, n446, n447, n448, n449;
    wire n450, n451, n452, n453, n454, n455, n456, n457;
    wire n458, n459, n460, n461, n462, n463, n464, n465;
    wire n466, n467, n468, n469, n470, n471, n472, n473;
    wire n474, n475, n476, n477, n478, n479, n480, n481;
    wire n482, n483, n484, n485, n486, n487, n488, n489;
    wire n490, n491, n492, n493, n494, n495, n496, n497;
    wire n498, n499, n500, n501, n502, n503, n504, n505;
    wire n506, n507, n508, n509, n510, n511, n512, n513;
    wire n514, n515, n516, n517, n518, n519, n520, n521;
    wire n522, n523, n524, n525, n526, n527, n528, n529;
    wire n530, n531, n532, n533, n534, n535, n536, n537;
    wire n538, n539, n540, n541, n542, n543, n544, n545;
    wire n546, n547, n548, n549, n550, n551, n552, n553;
    wire n554, n555, n556, n557, n558, n559, n560, n561;
    wire n562, n563, n564, n565, n566, n567, n568, n569;
    wire n570, n571, n572, n573, n574, n575, n576, n577;
    wire n578, n579, n580, n581, n582, n583, n584, n585;
    wire n586, n587, n588, n589, n590, n591, n592, n593;
    wire n594, n595, n596, n597, n598, n599, n600, n601;
    wire n602, n603, n604, n605, n606, n607, n608, n609;
    wire n610, n611, n612, n613, n614, n615, n616, n617;
    wire n618, n619, n620, n621, n622, n623, n624, n625;
    wire n626, n627, n628, n629, n630, n631, n632, n633;
    wire n634, n635, n636, n637, n638, n639, n640, n641;
    wire n642, n643, n644, n645, n646, n647, n648, n649;
    wire n650, n651, n652, n653, n654, n655, n656, n657;
    wire n658, n659, n660, n661, n662, n663, n664, n665;
    wire n666, n667, n668, n669, n670, n671, n672, n673;
    wire n674, n675, n676, n677, n678, n679, n680, n681;
    wire n682, n683, n684, n685, n686, n687, n688, n689;
    wire n690, n691, n692, n693, n694, n695, n696, n697;
    wire n698, n699, n700, n701, n702, n703, n704, n705;
    wire n706, n707, n708, n709, n710, n711, n712, n713;
    wire n714, n715, n716, n717, n718, n719, n720, n721;
    wire n722, n723, n724, n725, n726, n727, n728, n729;
    wire n730, n731, n732, n733, n734, n735, n736, n737;
    wire n738, n739, n740, n741, n742, n743, n744, n745;
    wire n746, n747, n748, n749, n750, n751, n752, n753;
    wire n754, n755, n756, n757, n758, n759, n760, n761;
    wire n762, n763, n764, n765, n766, n767, n768, n769;
    wire n770, n771, n772, n773, n774, n775, n776, n777;
    wire n778, n779, n780, n781, n782, n783, n784, n785;
    wire n786, n787, n788, n789, n790, n791, n792, n793;
    wire n794, n795, n796, n797, n798, n799, n800, n801;
    wire n802, n803, n804, n805, n806, n807, n808, n809;
    wire n810, n811, n812, n813, n814, n815, n816, n817;
    wire n818, n819, n820, n821, n822, n823, n824, n825;
    wire n826, n827, n828, n829, n830, n831, n832, n833;
    wire n834, n835, n836, n837, n838, n839, n840, n841;
    wire n842, n843, n844, n845, n846, n847, n848, n849;
    wire n850, n851, n852, n853, n854, n855, n856, n857;
    wire n858, n859, n860, n861, n862, n863, n864, n865;
    wire n866, n867, n868, n869, n870, n871, n872, n873;
    wire n874, n875, n876, n877, n878, n879, n880, n881;
    wire n882, n883, n884, n885, n886, n887, n888, n889;
    wire n890, n891, n892, n893, n894, n895, n896, n897;
    wire n898, n899, n900, n901, n902, n903, n904, n905;
    wire n906, n907, n908, n909, n910, n911, n912, n913;
    wire n914, n915, n916, n917, n918, n919, n920, n921;
    wire n922, n923, n924, n925, n926, n927, n928, n929;
    wire n930, n931, n932, n933, n934, n935, n936, n937;
    wire n938, n939, n940, n941, n942, n943, n944, n945;
    wire n946, n947, n948, n949, n950, n951, n952, n953;
    wire n954, n955, n956, n957, n958, n959, n960, n961;
    wire n962, n963, n964, n965, n966, n967, n968, n969;
    wire n970, n971, n972, n973, n974, n975, n976, n977;
    wire n978, n979, n980, n981, n982, n983, n984, n985;
    wire n986, n987, n988, n989, n990, n991, n992, n993;
    wire n994, n995, n996, n997, n998, n999, n1000, n1001;
    wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
    wire n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
    wire n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
    wire n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
    wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
    wire n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049;
    wire n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
    wire n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065;
    wire n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
    wire n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081;
    wire n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089;
    wire n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097;
    wire n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105;
    wire n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113;
    wire n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121;
    wire n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129;
    wire n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137;
    wire n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145;
    wire n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153;
    wire n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161;
    wire n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169;
    wire n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177;
    wire n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185;
    wire n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193;
    wire n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201;
    wire n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209;
    wire n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217;
    wire n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225;
    wire n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;
    wire n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241;
    wire n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249;
    wire n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;
    wire n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265;
    wire n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;
    wire n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;
    wire n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289;
    wire n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297;
    wire n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;
    wire n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313;
    wire n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321;
    wire n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329;
    wire n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;
    wire n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;
    wire n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;
    wire n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;
    wire n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369;
    wire n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;
    wire n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;
    wire n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393;
    wire n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401;
    wire n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;
    wire n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417;
    wire n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425;
    wire n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433;
    wire n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441;
    wire n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449;
    wire n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457;
    wire n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465;
    wire n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473;
    wire n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481;
    wire n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
    wire n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497;
    wire n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505;
    wire n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513;
    wire n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
    wire n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529;
    wire n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537;
    wire n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545;
    wire n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553;
    wire n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561;
    wire n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569;
    wire n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577;
    wire n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585;
    wire n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593;
    wire n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601;
    wire n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609;
    wire n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617;
    wire n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625;
    wire n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633;
    wire n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
    wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
    wire n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657;
    wire n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665;
    wire n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673;
    wire n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681;
    wire n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689;
    wire n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
    wire n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705;
    wire n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713;
    wire n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721;
    wire n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729;
    wire n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737;
    wire n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745;
    wire n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753;
    wire n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
    wire n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769;
    wire n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777;
    wire n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785;
    wire n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793;
    wire n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801;
    wire n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809;
    wire n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817;
    wire n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825;
    wire n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833;
    wire n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
    wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
    wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857;
    wire n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865;
    wire n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
    wire n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
    wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
    wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897;
    wire n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905;
    wire n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913;
    wire n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
    wire n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929;
    wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
    wire n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945;
    wire n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953;
    wire n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961;
    wire n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969;
    wire n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977;
    wire n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985;
    wire n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993;
    wire n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001;
    wire n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
    wire n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017;
    wire n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025;
    wire n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033;
    wire n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
    wire n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049;
    wire n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057;
    wire n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065;
    wire n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073;
    wire n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081;
    wire n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089;
    wire n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097;
    wire n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105;
    wire n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113;
    wire n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
    wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
    wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137;
    wire n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145;
    wire n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153;
    wire n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
    wire n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169;
    wire n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177;
    wire n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185;
    wire n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193;
    wire n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201;
    wire n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209;
    wire n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217;
    wire n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225;
    wire n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233;
    wire n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241;
    wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
    wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257;
    wire n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265;
    wire n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273;
    wire n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281;
    wire n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289;
    wire n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297;
    wire n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305;
    wire n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313;
    wire n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321;
    wire n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329;
    wire n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337;
    wire n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345;
    wire n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353;
    wire n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361;
    wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
    wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377;
    wire n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385;
    wire n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
    wire n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
    wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
    wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417;
    wire n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425;
    wire n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433;
    wire n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
    wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
    wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457;
    wire n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465;
    wire n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473;
    wire n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
    wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
    wire n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497;
    wire n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505;
    wire n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513;
    wire n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521;
    wire n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529;
    wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537;
    wire n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545;
    wire n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
    wire n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
    wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569;
    wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
    wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
    wire n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593;
    wire n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
    wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609;
    wire n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617;
    wire n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625;
    wire n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633;
    wire n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641;
    wire n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649;
    wire n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657;
    wire n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665;
    wire n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673;
    wire n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681;
    wire n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689;
    wire n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697;
    wire n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705;
    wire n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713;
    wire n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721;
    wire n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729;
    wire n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737;
    wire n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745;
    wire n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753;
    wire n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761;
    wire n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769;
    wire n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777;
    wire n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785;
    wire n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793;
    wire n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
    wire n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809;
    wire n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817;
    wire n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825;
    wire n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833;
    wire n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841;
    wire n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849;
    wire n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857;
    wire n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865;
    wire n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873;
    wire n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881;
    wire n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889;
    wire n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897;
    wire n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905;
    wire n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913;
    wire n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921;
    wire n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929;
    wire n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937;
    wire n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945;
    wire n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953;
    wire n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961;
    wire n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969;
    wire n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977;
    wire n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985;
    wire n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993;
    wire n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001;
    wire n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009;
    wire n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017;
    wire n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025;
    wire n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033;
    wire n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041;
    wire n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049;
    wire n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057;
    wire n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065;
    wire n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073;
    wire n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081;
    wire n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089;
    wire n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097;
    wire n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105;
    wire n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113;
    wire n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121;
    wire n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129;
    wire n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137;
    wire n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145;
    wire n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153;
    wire n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161;
    wire n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169;
    wire n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177;
    wire n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185;
    wire n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193;
    wire n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201;
    wire n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209;
    wire n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217;
    wire n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225;
    wire n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233;
    wire n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241;
    wire n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249;
    wire n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257;
    wire n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265;
    wire n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273;
    wire n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281;
    wire n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289;
    wire n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297;
    wire n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305;
    wire n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313;
    wire n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321;
    wire n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329;
    wire n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337;
    wire n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345;
    wire n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353;
    wire n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361;
    wire n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369;
    wire n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377;
    wire n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385;
    wire n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393;
    wire n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401;
    wire n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409;
    wire n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417;
    wire n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425;
    wire n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433;
    wire n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441;
    wire n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449;
    wire n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457;
    wire n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465;
    wire n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473;
    wire n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481;
    wire n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489;
    wire n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497;
    wire n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505;
    wire n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513;
    wire n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521;
    wire n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529;
    wire n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537;
    wire n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545;
    wire n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553;
    wire n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561;
    wire n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569;
    wire n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577;
    wire n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585;
    wire n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593;
    wire n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601;
    wire n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609;
    wire n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617;
    wire n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625;
    wire n3626, n3627, n3628, n3629, n3630;
    not g0(n2959 ,n6[1]);
    or g1(n3089 ,n2926 ,n2852);
    or g2(n3150 ,n2938 ,n2821);
    or g3(n3148 ,n2931 ,n2838);
    or g4(n3145 ,n2942 ,n2890);
    or g5(n3126 ,n2949 ,n2870);
    or g6(n3100 ,n2948 ,n2872);
    or g7(n3157 ,n2954 ,n2876);
    or g8(n3156 ,n2954 ,n2874);
    or g9(n3155 ,n2954 ,n2873);
    or g10(n3099 ,n2947 ,n2867);
    or g11(n3154 ,n2954 ,n2871);
    or g12(n3153 ,n2954 ,n2869);
    or g13(n3125 ,n2946 ,n2865);
    or g14(n3152 ,n2954 ,n2878);
    or g15(n3098 ,n2945 ,n2866);
    or g16(n3138 ,n2943 ,n2861);
    or g17(n3124 ,n2941 ,n2862);
    or g18(n3097 ,n2944 ,n2864);
    or g19(n3096 ,n2940 ,n2863);
    or g20(n3123 ,n2937 ,n2895);
    or g21(n3095 ,n2939 ,n2860);
    or g22(n3144 ,n2927 ,n2845);
    or g23(n3137 ,n2934 ,n2759);
    or g24(n3094 ,n2936 ,n2884);
    or g25(n3093 ,n2935 ,n2901);
    or g26(n3122 ,n2933 ,n2950);
    or g27(n3092 ,n2932 ,n2916);
    or g28(n3091 ,n2930 ,n2857);
    or g29(n3136 ,n2925 ,n2847);
    or g30(n3121 ,n2929 ,n2854);
    or g31(n3090 ,n2928 ,n2855);
    or g32(n3120 ,n2923 ,n2848);
    or g33(n3151 ,n2924 ,n2827);
    or g34(n3088 ,n2922 ,n2849);
    or g35(n3147 ,n2906 ,n2794);
    or g36(n3143 ,n2914 ,n2818);
    or g37(n3135 ,n2919 ,n2833);
    or g38(n3119 ,n2920 ,n2841);
    or g39(n3215 ,n2951 ,n2846);
    or g40(n3214 ,n2951 ,n2844);
    or g41(n3213 ,n2951 ,n2842);
    or g42(n3212 ,n2951 ,n2770);
    or g43(n3118 ,n2918 ,n2836);
    or g44(n3211 ,n2951 ,n2837);
    or g45(n3210 ,n2951 ,n2835);
    or g46(n3209 ,n2951 ,n2834);
    or g47(n3117 ,n2917 ,n2830);
    or g48(n3208 ,n2951 ,n2832);
    or g49(n3207 ,n2952 ,n2831);
    or g50(n3134 ,n2913 ,n2822);
    or g51(n3116 ,n2912 ,n2825);
    or g52(n3206 ,n2952 ,n2829);
    or g53(n3205 ,n2952 ,n2797);
    or g54(n3115 ,n2910 ,n2851);
    or g55(n3204 ,n2952 ,n2824);
    or g56(n3203 ,n2952 ,n2823);
    or g57(n3202 ,n2952 ,n2816);
    or g58(n3133 ,n2909 ,n2811);
    or g59(n3201 ,n2952 ,n2820);
    or g60(n3200 ,n2952 ,n2840);
    or g61(n3199 ,n2953 ,n2859);
    or g62(n3114 ,n2907 ,n2815);
    or g63(n3198 ,n2953 ,n2814);
    or g64(n3197 ,n2953 ,n2812);
    or g65(n3177 ,n2955 ,n2778);
    or g66(n3142 ,n2903 ,n2800);
    or g67(n3132 ,n2904 ,n2802);
    or g68(n3113 ,n2905 ,n2808);
    or g69(n3196 ,n2953 ,n2856);
    or g70(n3195 ,n2953 ,n2810);
    or g71(n3112 ,n2902 ,n2804);
    or g72(n3194 ,n2953 ,n2880);
    or g73(n3193 ,n2953 ,n2807);
    or g74(n3192 ,n2953 ,n2806);
    or g75(n3131 ,n2898 ,n2790);
    or g76(n3111 ,n2900 ,n2796);
    or g77(n3191 ,n2958 ,n2803);
    or g78(n3190 ,n2958 ,n2766);
    or g79(n3189 ,n2958 ,n2798);
    or g80(n3188 ,n2958 ,n2763);
    or g81(n3187 ,n2958 ,n2795);
    or g82(n3141 ,n2893 ,n2777);
    or g83(n3110 ,n2897 ,n2792);
    or g84(n3186 ,n2958 ,n2793);
    or g85(n3185 ,n2958 ,n2791);
    or g86(n3109 ,n2896 ,n2786);
    or g87(n3184 ,n2958 ,n2789);
    or g88(n3183 ,n2955 ,n2787);
    or g89(n3130 ,n2894 ,n2779);
    or g90(n3108 ,n2892 ,n2781);
    or g91(n3182 ,n2955 ,n2784);
    or g92(n3181 ,n2955 ,n2775);
    or g93(n3180 ,n2955 ,n2782);
    or g94(n3107 ,n2891 ,n2776);
    or g95(n3179 ,n2955 ,n2780);
    or g96(n3178 ,n2955 ,n2783);
    or g97(n3149 ,n2885 ,n2875);
    or g98(n3146 ,n2888 ,n2850);
    or g99(n3140 ,n2886 ,n2799);
    or g100(n3129 ,n2889 ,n2813);
    or g101(n3176 ,n2955 ,n2788);
    or g102(n3175 ,n2956 ,n2774);
    or g103(n3106 ,n2899 ,n2773);
    or g104(n3174 ,n2956 ,n2805);
    or g105(n3173 ,n2956 ,n2785);
    or g106(n3128 ,n2911 ,n2767);
    or g107(n3105 ,n2887 ,n2817);
    or g108(n3172 ,n2956 ,n2809);
    or g109(n3171 ,n2956 ,n2772);
    or g110(n3170 ,n2956 ,n2826);
    or g111(n3104 ,n2915 ,n2769);
    or g112(n3169 ,n2956 ,n2771);
    or g113(n3168 ,n2956 ,n2819);
    or g114(n3167 ,n2957 ,n2768);
    or g115(n3139 ,n2921 ,n2868);
    or g116(n3127 ,n2881 ,n2760);
    or g117(n3103 ,n2883 ,n2764);
    or g118(n3166 ,n2957 ,n2828);
    or g119(n3165 ,n2957 ,n2765);
    or g120(n3164 ,n2957 ,n2839);
    or g121(n3163 ,n2957 ,n2801);
    or g122(n3102 ,n2882 ,n2761);
    or g123(n3162 ,n2957 ,n2843);
    or g124(n3161 ,n2957 ,n2762);
    or g125(n3160 ,n2957 ,n2853);
    or g126(n3101 ,n2879 ,n2877);
    or g127(n3159 ,n2954 ,n2858);
    or g128(n3158 ,n2954 ,n2908);
    nor g129(n2950 ,n2621 ,n2648);
    nor g130(n2949 ,n2656 ,n2686);
    nor g131(n2948 ,n2657 ,n2691);
    nor g132(n2947 ,n2656 ,n2638);
    nor g133(n2946 ,n2651 ,n2566);
    nor g134(n2945 ,n2655 ,n2740);
    nor g135(n2944 ,n2659 ,n2633);
    nor g136(n2943 ,n2653 ,n2629);
    nor g137(n2942 ,n2651 ,n2628);
    nor g138(n2941 ,n2651 ,n2565);
    nor g139(n2940 ,n2659 ,n2554);
    nor g140(n2939 ,n2653 ,n2586);
    nor g141(n2938 ,n2651 ,n2666);
    nor g142(n2937 ,n2656 ,n2585);
    nor g143(n2936 ,n2655 ,n2564);
    nor g144(n2935 ,n2656 ,n2719);
    nor g145(n2934 ,n2657 ,n2622);
    nor g146(n2933 ,n2659 ,n2563);
    nor g147(n2932 ,n2655 ,n2553);
    nor g148(n2931 ,n2655 ,n2549);
    nor g149(n2930 ,n2656 ,n2582);
    nor g150(n2929 ,n2656 ,n2705);
    nor g151(n2928 ,n2658 ,n2618);
    nor g152(n2927 ,n2652 ,n2609);
    nor g153(n2926 ,n2657 ,n2700);
    nor g154(n2925 ,n2658 ,n2560);
    nor g155(n2924 ,n2653 ,n2744);
    nor g156(n2923 ,n2658 ,n2613);
    nor g157(n2922 ,n2659 ,n2697);
    nor g158(n2921 ,n2657 ,n2636);
    nor g159(n2920 ,n2658 ,n2684);
    nor g160(n2919 ,n2658 ,n2672);
    nor g161(n2918 ,n2659 ,n2674);
    nor g162(n2917 ,n2658 ,n2676);
    nor g163(n2916 ,n2583 ,n2545);
    nor g164(n2915 ,n2652 ,n2734);
    nor g165(n2914 ,n2658 ,n2742);
    nor g166(n2913 ,n2656 ,n2631);
    nor g167(n2912 ,n2655 ,n2750);
    nor g168(n2911 ,n2657 ,n2607);
    nor g169(n2910 ,n2652 ,n2639);
    nor g170(n2909 ,n2653 ,n2614);
    nor g171(n2908 ,n2723 ,n2650);
    nor g172(n2907 ,n2653 ,n2711);
    nor g173(n2906 ,n2652 ,n2646);
    nor g174(n2905 ,n2652 ,n2703);
    nor g175(n2904 ,n2653 ,n2682);
    nor g176(n2903 ,n2655 ,n2668);
    nor g177(n2902 ,n2651 ,n2732);
    nor g178(n2901 ,n2624 ,n2545);
    nor g179(n2900 ,n2651 ,n2568);
    nor g180(n2899 ,n2652 ,n2755);
    nor g181(n2898 ,n2652 ,n2663);
    nor g182(n2897 ,n2652 ,n2599);
    nor g183(n2896 ,n2659 ,n2597);
    nor g184(n2895 ,n2625 ,n2544);
    nor g185(n2894 ,n2657 ,n2600);
    nor g186(n2893 ,n2653 ,n2603);
    nor g187(n2892 ,n2656 ,n2572);
    nor g188(n2891 ,n2655 ,n2660);
    nor g189(n2890 ,n2584 ,n2648);
    nor g190(n2889 ,n2657 ,n2749);
    nor g191(n2888 ,n2651 ,n2725);
    nor g192(n2887 ,n2653 ,n2715);
    nor g193(n2886 ,n2655 ,n2722);
    nor g194(n2885 ,n2651 ,n2706);
    nor g195(n2884 ,n2626 ,n2650);
    nor g196(n2883 ,n2657 ,n2726);
    nor g197(n2882 ,n2659 ,n2642);
    nor g198(n2881 ,n2658 ,n2620);
    nor g199(n2880 ,n2721 ,n2545);
    nor g200(n2879 ,n2659 ,n2704);
    nor g201(n2878 ,n2696 ,n2650);
    nor g202(n2877 ,n2592 ,n2650);
    nor g203(n2876 ,n2733 ,n2650);
    nor g204(n2875 ,n2634 ,n2650);
    nor g205(n2874 ,n2690 ,n2648);
    nor g206(n2873 ,n2694 ,n2544);
    nor g207(n2872 ,n2641 ,n2545);
    nor g208(n2871 ,n2590 ,n2650);
    nor g209(n2870 ,n2546 ,n2648);
    nor g210(n2869 ,n2555 ,n2544);
    nor g211(n2868 ,n2589 ,n2648);
    nor g212(n2867 ,n2637 ,n2648);
    nor g213(n2866 ,n2588 ,n2544);
    nor g214(n2865 ,n2737 ,n2648);
    nor g215(n2864 ,n2632 ,n2544);
    nor g216(n2863 ,n2587 ,n2544);
    nor g217(n2862 ,n2727 ,n2545);
    nor g218(n2861 ,n2627 ,n2648);
    nor g219(n2860 ,n2724 ,n2545);
    nor g220(n2859 ,n2619 ,n2650);
    nor g221(n2958 ,n2687 ,n2654);
    nor g222(n2957 ,n2736 ,n2654);
    nor g223(n2956 ,n2754 ,n2654);
    nor g224(n2955 ,n2664 ,n2654);
    nor g225(n2954 ,n2581 ,n2654);
    nor g226(n2953 ,n2683 ,n2654);
    nor g227(n2952 ,n2675 ,n2654);
    nor g228(n2951 ,n2610 ,n2654);
    nor g229(n2858 ,n2548 ,n2648);
    nor g230(n2857 ,n2709 ,n2544);
    nor g231(n2856 ,n2708 ,n2544);
    nor g232(n2855 ,n2617 ,n2650);
    nor g233(n2854 ,n2616 ,n2544);
    nor g234(n2853 ,n2552 ,n2648);
    nor g235(n2852 ,n2561 ,n2545);
    nor g236(n2851 ,n2630 ,n2544);
    nor g237(n2850 ,n2701 ,n2545);
    nor g238(n2849 ,n2578 ,n2545);
    nor g239(n2848 ,n2577 ,n2648);
    nor g240(n2847 ,n2608 ,n2545);
    nor g241(n2846 ,n2576 ,n2545);
    nor g242(n2845 ,n2680 ,n2545);
    nor g243(n2844 ,n2567 ,n2648);
    nor g244(n2843 ,n2716 ,n2648);
    nor g245(n2842 ,n2591 ,n2545);
    nor g246(n2841 ,n2667 ,n2545);
    nor g247(n2840 ,n2640 ,n2545);
    nor g248(n2839 ,n2557 ,n2648);
    nor g249(n2838 ,n2606 ,n2545);
    nor g250(n2837 ,n2551 ,n2544);
    nor g251(n2836 ,n2673 ,n2650);
    nor g252(n2835 ,n2601 ,n2544);
    nor g253(n2834 ,n2671 ,n2648);
    nor g254(n2833 ,n2662 ,n2648);
    nor g255(n2832 ,n2717 ,n2545);
    nor g256(n2831 ,n2679 ,n2544);
    nor g257(n2830 ,n2677 ,n2648);
    nor g258(n2829 ,n2643 ,n2544);
    nor g259(n2828 ,n2718 ,n2648);
    nor g260(n2827 ,n2670 ,n2545);
    nor g261(n2826 ,n2738 ,n2544);
    nor g262(n2825 ,n2635 ,n2650);
    nor g263(n2824 ,n2623 ,n2650);
    nor g264(n2823 ,n2743 ,n2545);
    nor g265(n2822 ,n2731 ,n2650);
    nor g266(n2821 ,n2707 ,n2545);
    nor g267(n2820 ,n2547 ,n2545);
    nor g268(n2819 ,n2741 ,n2544);
    nor g269(n2818 ,n2757 ,n2650);
    nor g270(n2817 ,n2712 ,n2650);
    nor g271(n2816 ,n2739 ,n2545);
    nor g272(n2815 ,n2579 ,n2650);
    nor g273(n2814 ,n2713 ,n2650);
    nor g274(n2813 ,n2748 ,n2648);
    nor g275(n2812 ,n2710 ,n2544);
    nor g276(n2811 ,n2615 ,n2650);
    nor g277(n2810 ,n2702 ,n2650);
    nor g278(n2809 ,n2751 ,n2544);
    nor g279(n2808 ,n2753 ,n2544);
    nor g280(n2807 ,n2695 ,n2648);
    nor g281(n2806 ,n2693 ,n2650);
    nor g282(n2805 ,n2756 ,n2544);
    nor g283(n2804 ,n2689 ,n2650);
    nor g284(n2803 ,n2752 ,n2545);
    nor g285(n2802 ,n2593 ,n2545);
    nor g286(n2801 ,n2685 ,n2648);
    nor g287(n2800 ,n2556 ,n2545);
    nor g288(n2799 ,n2720 ,n2545);
    nor g289(n2798 ,n2644 ,n2545);
    nor g290(n2797 ,n2747 ,n2544);
    nor g291(n2796 ,n2595 ,n2650);
    nor g292(n2795 ,n2569 ,n2544);
    nor g293(n2794 ,n2571 ,n2544);
    nor g294(n2793 ,n2605 ,n2650);
    nor g295(n2792 ,n2661 ,n2648);
    nor g296(n2791 ,n2596 ,n2650);
    nor g297(n2790 ,n2558 ,n2648);
    nor g298(n2789 ,n2570 ,n2544);
    nor g299(n2788 ,n2574 ,n2650);
    nor g300(n2787 ,n2550 ,n2545);
    nor g301(n2786 ,n2669 ,n2650);
    nor g302(n2785 ,n2611 ,n2544);
    nor g303(n2784 ,n2598 ,n2648);
    nor g304(n2783 ,n2665 ,n2648);
    nor g305(n2782 ,n2602 ,n2650);
    nor g306(n2781 ,n2681 ,n2650);
    nor g307(n2780 ,n2573 ,n2544);
    nor g308(n2779 ,n2575 ,n2648);
    nor g309(n2778 ,n2604 ,n2544);
    nor g310(n2777 ,n2758 ,n2545);
    nor g311(n2776 ,n2746 ,n2648);
    nor g312(n2775 ,n2692 ,n2650);
    nor g313(n2774 ,n2559 ,n2544);
    nor g314(n2773 ,n2612 ,n2650);
    nor g315(n2772 ,n2688 ,n2650);
    nor g316(n2771 ,n2745 ,n2648);
    nor g317(n2770 ,n2645 ,n2544);
    nor g318(n2769 ,n2730 ,n2544);
    nor g319(n2768 ,n2735 ,n2545);
    nor g320(n2767 ,n2729 ,n2648);
    nor g321(n2766 ,n2678 ,n2545);
    nor g322(n2765 ,n2728 ,n2648);
    nor g323(n2764 ,n2714 ,n2544);
    nor g324(n2763 ,n2594 ,n2648);
    nor g325(n2762 ,n2699 ,n2650);
    nor g326(n2761 ,n2580 ,n2544);
    nor g327(n2760 ,n2698 ,n2648);
    nor g328(n2759 ,n2562 ,n2545);
    not g329(n2758 ,n2[53]);
    not g330(n2757 ,n2[55]);
    not g331(n2756 ,n2[86]);
    not g332(n2755 ,n3[18]);
    not g333(n2754 ,n7[23]);
    not g334(n2753 ,n2[25]);
    not g335(n2752 ,n2[103]);
    not g336(n2751 ,n2[84]);
    not g337(n2750 ,n3[28]);
    not g338(n2749 ,n3[41]);
    not g339(n2748 ,n2[41]);
    not g340(n2747 ,n2[117]);
    not g341(n2746 ,n2[19]);
    not g342(n2745 ,n2[81]);
    not g343(n2744 ,n3[63]);
    not g344(n2743 ,n2[115]);
    not g345(n2742 ,n3[55]);
    not g346(n2741 ,n2[80]);
    not g347(n2740 ,n3[10]);
    not g348(n2739 ,n2[114]);
    not g349(n2738 ,n2[82]);
    not g350(n2737 ,n2[37]);
    not g351(n2736 ,n7[15]);
    not g352(n2735 ,n2[79]);
    not g353(n2734 ,n3[16]);
    not g354(n2733 ,n2[69]);
    not g355(n2732 ,n3[24]);
    not g356(n2731 ,n2[46]);
    not g357(n2730 ,n2[16]);
    not g358(n2729 ,n2[40]);
    not g359(n2728 ,n2[77]);
    not g360(n2727 ,n2[36]);
    not g361(n2726 ,n3[15]);
    not g362(n2725 ,n3[58]);
    not g363(n2724 ,n2[7]);
    not g364(n2723 ,n2[70]);
    not g365(n2722 ,n3[52]);
    not g366(n2721 ,n2[106]);
    not g367(n2720 ,n2[52]);
    not g368(n2719 ,n3[5]);
    not g369(n2718 ,n2[78]);
    not g370(n2717 ,n2[120]);
    not g371(n2716 ,n2[74]);
    not g372(n2715 ,n3[17]);
    not g373(n2714 ,n2[15]);
    not g374(n2713 ,n2[110]);
    not g375(n2712 ,n2[17]);
    not g376(n2711 ,n3[26]);
    not g377(n2710 ,n2[109]);
    not g378(n2709 ,n2[3]);
    not g379(n2708 ,n2[108]);
    not g380(n2707 ,n2[62]);
    not g381(n2706 ,n3[61]);
    not g382(n2705 ,n3[33]);
    not g383(n2704 ,n3[13]);
    not g384(n2703 ,n3[25]);
    not g385(n2702 ,n2[107]);
    not g386(n2701 ,n2[58]);
    not g387(n2700 ,n3[1]);
    not g388(n2699 ,n2[73]);
    not g389(n2698 ,n2[39]);
    not g390(n2697 ,n3[0]);
    not g391(n2696 ,n2[64]);
    not g392(n2695 ,n2[105]);
    not g393(n2694 ,n2[67]);
    not g394(n2693 ,n2[104]);
    not g395(n2692 ,n2[93]);
    not g396(n2691 ,n3[12]);
    not g397(n2690 ,n2[68]);
    not g398(n2689 ,n2[24]);
    not g399(n2688 ,n2[83]);
    not g400(n2687 ,n7[39]);
    not g401(n2686 ,n3[38]);
    not g402(n2685 ,n2[75]);
    not g403(n2684 ,n3[31]);
    not g404(n2683 ,n7[47]);
    not g405(n2682 ,n3[44]);
    not g406(n2681 ,n2[20]);
    not g407(n2680 ,n2[56]);
    not g408(n2679 ,n2[119]);
    not g409(n2678 ,n2[102]);
    not g410(n2677 ,n2[29]);
    not g411(n2676 ,n3[29]);
    not g412(n2675 ,n7[55]);
    not g413(n2674 ,n3[30]);
    not g414(n2673 ,n2[30]);
    not g415(n2672 ,n3[47]);
    not g416(n2671 ,n2[121]);
    not g417(n2670 ,n2[63]);
    not g418(n2669 ,n2[21]);
    not g419(n2668 ,n3[54]);
    not g420(n2667 ,n2[31]);
    not g421(n2666 ,n3[62]);
    not g422(n2665 ,n2[90]);
    not g423(n2664 ,n7[31]);
    not g424(n2663 ,n3[43]);
    not g425(n2662 ,n2[47]);
    not g426(n2661 ,n2[22]);
    not g427(n2660 ,n3[19]);
    not g428(n2659 ,n6[2]);
    not g429(n2658 ,n6[2]);
    not g430(n2657 ,n6[2]);
    not g431(n2656 ,n6[2]);
    not g432(n2655 ,n6[2]);
    not g433(n2654 ,n6[2]);
    not g434(n2653 ,n6[2]);
    not g435(n2652 ,n6[2]);
    not g436(n2651 ,n6[2]);
    not g437(n2650 ,n2649);
    not g438(n2545 ,n2649);
    not g439(n2649 ,n2959);
    not g440(n2648 ,n2647);
    not g441(n2544 ,n2647);
    not g442(n2647 ,n2959);
    not g443(n2646 ,n3[59]);
    not g444(n2645 ,n2[124]);
    not g445(n2644 ,n2[101]);
    not g446(n2643 ,n2[118]);
    not g447(n2642 ,n3[14]);
    not g448(n2641 ,n2[12]);
    not g449(n2640 ,n2[112]);
    not g450(n2639 ,n3[27]);
    not g451(n2638 ,n3[11]);
    not g452(n2637 ,n2[11]);
    not g453(n2636 ,n3[51]);
    not g454(n2635 ,n2[28]);
    not g455(n2634 ,n2[61]);
    not g456(n2633 ,n3[9]);
    not g457(n2632 ,n2[9]);
    not g458(n2631 ,n3[46]);
    not g459(n2630 ,n2[27]);
    not g460(n2629 ,n3[50]);
    not g461(n2628 ,n3[57]);
    not g462(n2627 ,n2[50]);
    not g463(n2626 ,n2[6]);
    not g464(n2625 ,n2[35]);
    not g465(n2624 ,n2[5]);
    not g466(n2623 ,n2[116]);
    not g467(n2622 ,n3[49]);
    not g468(n2621 ,n2[34]);
    not g469(n2620 ,n3[39]);
    not g470(n2619 ,n2[111]);
    not g471(n2618 ,n3[2]);
    not g472(n2617 ,n2[2]);
    not g473(n2616 ,n2[33]);
    not g474(n2615 ,n2[45]);
    not g475(n2614 ,n3[45]);
    not g476(n2613 ,n3[32]);
    not g477(n2612 ,n2[18]);
    not g478(n2611 ,n2[85]);
    not g479(n2610 ,n7[63]);
    not g480(n2609 ,n3[56]);
    not g481(n2608 ,n2[48]);
    not g482(n2607 ,n3[40]);
    not g483(n2606 ,n2[60]);
    not g484(n2605 ,n2[98]);
    not g485(n2604 ,n2[89]);
    not g486(n2603 ,n3[53]);
    not g487(n2602 ,n2[92]);
    not g488(n2601 ,n2[122]);
    not g489(n2600 ,n3[42]);
    not g490(n2599 ,n3[22]);
    not g491(n2598 ,n2[94]);
    not g492(n2597 ,n3[21]);
    not g493(n2596 ,n2[97]);
    not g494(n2595 ,n2[23]);
    not g495(n2594 ,n2[100]);
    not g496(n2593 ,n2[44]);
    not g497(n2592 ,n2[13]);
    not g498(n2591 ,n2[125]);
    not g499(n2590 ,n2[66]);
    not g500(n2589 ,n2[51]);
    not g501(n2588 ,n2[10]);
    not g502(n2587 ,n2[8]);
    not g503(n2586 ,n3[7]);
    not g504(n2585 ,n3[35]);
    not g505(n2584 ,n2[57]);
    not g506(n2583 ,n2[4]);
    not g507(n2582 ,n3[3]);
    not g508(n2581 ,n7[7]);
    not g509(n2580 ,n2[14]);
    not g510(n2579 ,n2[26]);
    not g511(n2578 ,n2[0]);
    not g512(n2577 ,n2[32]);
    not g513(n2576 ,n2[127]);
    not g514(n2575 ,n2[42]);
    not g515(n2574 ,n2[88]);
    not g516(n2573 ,n2[91]);
    not g517(n2572 ,n3[20]);
    not g518(n2571 ,n2[59]);
    not g519(n2570 ,n2[96]);
    not g520(n2569 ,n2[99]);
    not g521(n2568 ,n3[23]);
    not g522(n2567 ,n2[126]);
    not g523(n2566 ,n3[37]);
    not g524(n2565 ,n3[36]);
    not g525(n2564 ,n3[6]);
    not g526(n2563 ,n3[34]);
    not g527(n2562 ,n2[49]);
    not g528(n2561 ,n2[1]);
    not g529(n2560 ,n3[48]);
    not g530(n2559 ,n2[87]);
    not g531(n2558 ,n2[43]);
    not g532(n2557 ,n2[76]);
    not g533(n2556 ,n2[54]);
    not g534(n2555 ,n2[65]);
    not g535(n2554 ,n3[8]);
    not g536(n2553 ,n3[4]);
    not g537(n2552 ,n2[72]);
    not g538(n2551 ,n2[123]);
    not g539(n2550 ,n2[95]);
    not g540(n2549 ,n3[60]);
    not g541(n2548 ,n2[71]);
    not g542(n2547 ,n2[113]);
    not g543(n2546 ,n2[38]);
    dff g544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2471), .Q(n5[0]));
    dff g545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2447), .Q(n5[1]));
    dff g546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2527), .Q(n5[2]));
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2541), .Q(n5[3]));
    dff g548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2531), .Q(n5[4]));
    dff g549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2523), .Q(n5[5]));
    dff g550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2518), .Q(n5[6]));
    dff g551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2516), .Q(n5[7]));
    dff g552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2513), .Q(n5[8]));
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2506), .Q(n5[9]));
    dff g554(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2502), .Q(n5[10]));
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2498), .Q(n5[11]));
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2494), .Q(n5[12]));
    dff g557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2489), .Q(n5[13]));
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2490), .Q(n5[14]));
    dff g559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2488), .Q(n5[15]));
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2487), .Q(n5[16]));
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2485), .Q(n5[17]));
    dff g562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2486), .Q(n5[18]));
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2484), .Q(n5[19]));
    dff g564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2483), .Q(n5[20]));
    dff g565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2482), .Q(n5[21]));
    dff g566(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2481), .Q(n5[22]));
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2480), .Q(n5[23]));
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2477), .Q(n5[24]));
    dff g569(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2479), .Q(n5[25]));
    dff g570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2478), .Q(n5[26]));
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2476), .Q(n5[27]));
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2475), .Q(n5[28]));
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2474), .Q(n5[29]));
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2473), .Q(n5[30]));
    dff g575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2472), .Q(n5[31]));
    dff g576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2470), .Q(n5[32]));
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2468), .Q(n5[33]));
    dff g578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2469), .Q(n5[34]));
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2466), .Q(n5[35]));
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2467), .Q(n5[36]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2465), .Q(n5[37]));
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2464), .Q(n5[38]));
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2463), .Q(n5[39]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2462), .Q(n5[40]));
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2509), .Q(n5[41]));
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2460), .Q(n5[42]));
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2459), .Q(n5[43]));
    dff g588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2458), .Q(n5[44]));
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2457), .Q(n5[45]));
    dff g590(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2454), .Q(n5[46]));
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2452), .Q(n5[47]));
    dff g592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2450), .Q(n5[48]));
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2445), .Q(n5[49]));
    dff g594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2441), .Q(n5[50]));
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2439), .Q(n5[51]));
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2437), .Q(n5[52]));
    dff g597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2434), .Q(n5[53]));
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2431), .Q(n5[54]));
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2429), .Q(n5[55]));
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2427), .Q(n5[56]));
    dff g601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2420), .Q(n5[57]));
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2421), .Q(n5[58]));
    dff g603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2418), .Q(n5[59]));
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2416), .Q(n5[60]));
    dff g605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2539), .Q(n5[61]));
    dff g606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2538), .Q(n5[62]));
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2536), .Q(n5[63]));
    dff g608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n771), .Q(n8[0]));
    dff g609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n775), .Q(n8[1]));
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n774), .Q(n8[2]));
    dff g611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n779), .Q(n8[3]));
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n778), .Q(n8[4]));
    dff g613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n783), .Q(n8[5]));
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n773), .Q(n8[6]));
    dff g615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n776), .Q(n8[7]));
    dff g616(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2365), .Q(n3[0]));
    dff g617(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2412), .Q(n3[1]));
    dff g618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2411), .Q(n3[2]));
    dff g619(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2410), .Q(n3[3]));
    dff g620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2409), .Q(n3[4]));
    dff g621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2408), .Q(n3[5]));
    dff g622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2407), .Q(n3[6]));
    dff g623(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2406), .Q(n3[7]));
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2405), .Q(n3[8]));
    dff g625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2404), .Q(n3[9]));
    dff g626(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2403), .Q(n3[10]));
    dff g627(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2402), .Q(n3[11]));
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2401), .Q(n3[12]));
    dff g629(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2400), .Q(n3[13]));
    dff g630(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2399), .Q(n3[14]));
    dff g631(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2398), .Q(n3[15]));
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2397), .Q(n3[16]));
    dff g633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2396), .Q(n3[17]));
    dff g634(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2395), .Q(n3[18]));
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n3[19]));
    dff g636(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2393), .Q(n3[20]));
    dff g637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n3[21]));
    dff g638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n3[22]));
    dff g639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2390), .Q(n3[23]));
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2389), .Q(n3[24]));
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2388), .Q(n3[25]));
    dff g642(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2387), .Q(n3[26]));
    dff g643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2386), .Q(n3[27]));
    dff g644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2385), .Q(n3[28]));
    dff g645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2384), .Q(n3[29]));
    dff g646(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2383), .Q(n3[30]));
    dff g647(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2382), .Q(n3[31]));
    dff g648(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2381), .Q(n3[32]));
    dff g649(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2380), .Q(n3[33]));
    dff g650(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n3[34]));
    dff g651(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n3[35]));
    dff g652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n3[36]));
    dff g653(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2376), .Q(n3[37]));
    dff g654(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2375), .Q(n3[38]));
    dff g655(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2374), .Q(n3[39]));
    dff g656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2373), .Q(n3[40]));
    dff g657(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2372), .Q(n3[41]));
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2371), .Q(n3[42]));
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2370), .Q(n3[43]));
    dff g660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2369), .Q(n3[44]));
    dff g661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2368), .Q(n3[45]));
    dff g662(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2367), .Q(n3[46]));
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2366), .Q(n3[47]));
    dff g664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2413), .Q(n3[48]));
    dff g665(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2364), .Q(n3[49]));
    dff g666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2363), .Q(n3[50]));
    dff g667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2362), .Q(n3[51]));
    dff g668(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2361), .Q(n3[52]));
    dff g669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2360), .Q(n3[53]));
    dff g670(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2359), .Q(n3[54]));
    dff g671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2358), .Q(n3[55]));
    dff g672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2357), .Q(n3[56]));
    dff g673(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2356), .Q(n3[57]));
    dff g674(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2355), .Q(n3[58]));
    dff g675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2354), .Q(n3[59]));
    dff g676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2353), .Q(n3[60]));
    dff g677(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n3[61]));
    dff g678(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2351), .Q(n3[62]));
    dff g679(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2350), .Q(n3[63]));
    dff g680(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n949), .Q(n6[0]));
    dff g681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n950), .Q(n2542));
    dff g682(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n951), .Q(n2543));
    dff g683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2456), .Q(n4[0]));
    dff g684(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2455), .Q(n4[1]));
    dff g685(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2453), .Q(n4[2]));
    dff g686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2451), .Q(n4[3]));
    dff g687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2449), .Q(n4[4]));
    dff g688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2448), .Q(n4[5]));
    dff g689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2446), .Q(n4[6]));
    dff g690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2444), .Q(n4[7]));
    dff g691(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2443), .Q(n4[8]));
    dff g692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2442), .Q(n4[9]));
    dff g693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2440), .Q(n4[10]));
    dff g694(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2438), .Q(n4[11]));
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2436), .Q(n4[12]));
    dff g696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2435), .Q(n4[13]));
    dff g697(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2433), .Q(n4[14]));
    dff g698(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2432), .Q(n4[15]));
    dff g699(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2430), .Q(n4[16]));
    dff g700(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2428), .Q(n4[17]));
    dff g701(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2426), .Q(n4[18]));
    dff g702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2425), .Q(n4[19]));
    dff g703(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2424), .Q(n4[20]));
    dff g704(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2423), .Q(n4[21]));
    dff g705(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2422), .Q(n4[22]));
    dff g706(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2419), .Q(n4[23]));
    dff g707(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n4[24]));
    dff g708(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2415), .Q(n4[25]));
    dff g709(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2414), .Q(n4[26]));
    dff g710(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2525), .Q(n4[27]));
    dff g711(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2540), .Q(n4[28]));
    dff g712(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2537), .Q(n4[29]));
    dff g713(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2535), .Q(n4[30]));
    dff g714(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2534), .Q(n4[31]));
    dff g715(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2533), .Q(n4[32]));
    dff g716(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2532), .Q(n4[33]));
    dff g717(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2530), .Q(n4[34]));
    dff g718(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2529), .Q(n4[35]));
    dff g719(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2528), .Q(n4[36]));
    dff g720(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2526), .Q(n4[37]));
    dff g721(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2524), .Q(n4[38]));
    dff g722(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2522), .Q(n4[39]));
    dff g723(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2521), .Q(n4[40]));
    dff g724(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2520), .Q(n4[41]));
    dff g725(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2519), .Q(n4[42]));
    dff g726(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2517), .Q(n4[43]));
    dff g727(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2515), .Q(n4[44]));
    dff g728(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2514), .Q(n4[45]));
    dff g729(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2512), .Q(n4[46]));
    dff g730(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2511), .Q(n4[47]));
    dff g731(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2510), .Q(n4[48]));
    dff g732(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2461), .Q(n4[49]));
    dff g733(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2508), .Q(n4[50]));
    dff g734(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2507), .Q(n4[51]));
    dff g735(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2505), .Q(n4[52]));
    dff g736(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2504), .Q(n4[53]));
    dff g737(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2503), .Q(n4[54]));
    dff g738(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2501), .Q(n4[55]));
    dff g739(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2500), .Q(n4[56]));
    dff g740(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2499), .Q(n4[57]));
    dff g741(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2497), .Q(n4[58]));
    dff g742(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2496), .Q(n4[59]));
    dff g743(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2495), .Q(n4[60]));
    dff g744(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2493), .Q(n4[61]));
    dff g745(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2492), .Q(n4[62]));
    dff g746(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2491), .Q(n4[63]));
    or g747(n2541 ,n1692 ,n2280);
    or g748(n2540 ,n1521 ,n2348);
    or g749(n2539 ,n1700 ,n2284);
    or g750(n2538 ,n1537 ,n2283);
    or g751(n2537 ,n1698 ,n2347);
    or g752(n2536 ,n1590 ,n2281);
    or g753(n2535 ,n1697 ,n2346);
    or g754(n2534 ,n1610 ,n2345);
    or g755(n2533 ,n1693 ,n2344);
    or g756(n2532 ,n1690 ,n2343);
    or g757(n2531 ,n1464 ,n2279);
    or g758(n2530 ,n1689 ,n2342);
    or g759(n2529 ,n1688 ,n2341);
    or g760(n2528 ,n1687 ,n2340);
    or g761(n2527 ,n1701 ,n2282);
    or g762(n2526 ,n1685 ,n2339);
    or g763(n2525 ,n1699 ,n2349);
    or g764(n2524 ,n1684 ,n2338);
    or g765(n2523 ,n1548 ,n2278);
    or g766(n2522 ,n1681 ,n2337);
    or g767(n2521 ,n1679 ,n2336);
    or g768(n2520 ,n1676 ,n2335);
    or g769(n2519 ,n1675 ,n2334);
    or g770(n2518 ,n1650 ,n2277);
    or g771(n2517 ,n1674 ,n2333);
    or g772(n2516 ,n1691 ,n2276);
    or g773(n2515 ,n1683 ,n2332);
    or g774(n2514 ,n1696 ,n2331);
    or g775(n2513 ,n1669 ,n2275);
    or g776(n2512 ,n1672 ,n2330);
    or g777(n2511 ,n1671 ,n2329);
    or g778(n2510 ,n1670 ,n2328);
    or g779(n2509 ,n1499 ,n2242);
    or g780(n2508 ,n1664 ,n2326);
    or g781(n2507 ,n1552 ,n2325);
    or g782(n2506 ,n1657 ,n2274);
    or g783(n2505 ,n1661 ,n2324);
    or g784(n2504 ,n1658 ,n2323);
    or g785(n2503 ,n1655 ,n2322);
    or g786(n2502 ,n1647 ,n2273);
    or g787(n2501 ,n1652 ,n2321);
    or g788(n2500 ,n1649 ,n2320);
    or g789(n2499 ,n1645 ,n2319);
    or g790(n2498 ,n1636 ,n2272);
    or g791(n2497 ,n1601 ,n2318);
    or g792(n2496 ,n1644 ,n2269);
    or g793(n2495 ,n1653 ,n2316);
    or g794(n2494 ,n1694 ,n2271);
    or g795(n2493 ,n1663 ,n2315);
    or g796(n2492 ,n1654 ,n2314);
    or g797(n2491 ,n1695 ,n2313);
    or g798(n2490 ,n1630 ,n2317);
    or g799(n2489 ,n1635 ,n2270);
    or g800(n2488 ,n1627 ,n2268);
    or g801(n2487 ,n1622 ,n2267);
    or g802(n2486 ,n1609 ,n2265);
    or g803(n2485 ,n1616 ,n2266);
    or g804(n2484 ,n1605 ,n2264);
    or g805(n2483 ,n1598 ,n2263);
    or g806(n2482 ,n1597 ,n2262);
    or g807(n2481 ,n1591 ,n2261);
    or g808(n2480 ,n1588 ,n2260);
    or g809(n2479 ,n1576 ,n2258);
    or g810(n2478 ,n1571 ,n2257);
    or g811(n2477 ,n1582 ,n2259);
    or g812(n2476 ,n1567 ,n2256);
    or g813(n2475 ,n1563 ,n2255);
    or g814(n2474 ,n1559 ,n2254);
    or g815(n2473 ,n1556 ,n2253);
    or g816(n2472 ,n1550 ,n2251);
    or g817(n2471 ,n1541 ,n2228);
    or g818(n2470 ,n1546 ,n2252);
    or g819(n2469 ,n1533 ,n2249);
    or g820(n2468 ,n1539 ,n2250);
    or g821(n2467 ,n1524 ,n2247);
    or g822(n2466 ,n1529 ,n2248);
    or g823(n2465 ,n1519 ,n2246);
    or g824(n2464 ,n1514 ,n2245);
    or g825(n2463 ,n1508 ,n2244);
    or g826(n2462 ,n1506 ,n2243);
    or g827(n2461 ,n1667 ,n2327);
    or g828(n2460 ,n1491 ,n2241);
    or g829(n2459 ,n1490 ,n2240);
    or g830(n2458 ,n1487 ,n2239);
    or g831(n2457 ,n1486 ,n2238);
    or g832(n2456 ,n1488 ,n2312);
    or g833(n2455 ,n1485 ,n2311);
    or g834(n2454 ,n1482 ,n2237);
    or g835(n2453 ,n1484 ,n2310);
    or g836(n2452 ,n1481 ,n2236);
    or g837(n2451 ,n1483 ,n2309);
    or g838(n2450 ,n1478 ,n2235);
    or g839(n2449 ,n1480 ,n2308);
    or g840(n2448 ,n1479 ,n2307);
    or g841(n2447 ,n1680 ,n2285);
    or g842(n2446 ,n1477 ,n2306);
    or g843(n2445 ,n1474 ,n2234);
    or g844(n2444 ,n1476 ,n2305);
    or g845(n2443 ,n1473 ,n2304);
    or g846(n2442 ,n1471 ,n2303);
    or g847(n2441 ,n1472 ,n2233);
    or g848(n2440 ,n1470 ,n2302);
    or g849(n2439 ,n1469 ,n2232);
    or g850(n2438 ,n1468 ,n2301);
    or g851(n2437 ,n1467 ,n2231);
    or g852(n2436 ,n1466 ,n2300);
    or g853(n2435 ,n1465 ,n2299);
    or g854(n2434 ,n1641 ,n2230);
    or g855(n2433 ,n1463 ,n2298);
    or g856(n2432 ,n1462 ,n2297);
    or g857(n2431 ,n1457 ,n2229);
    or g858(n2430 ,n1460 ,n2296);
    or g859(n2429 ,n1459 ,n2227);
    or g860(n2428 ,n1458 ,n2295);
    or g861(n2427 ,n1455 ,n2226);
    or g862(n2426 ,n1456 ,n2294);
    or g863(n2425 ,n1453 ,n2293);
    or g864(n2424 ,n1452 ,n2292);
    or g865(n2423 ,n1449 ,n2291);
    or g866(n2422 ,n1448 ,n2290);
    or g867(n2421 ,n1447 ,n2224);
    or g868(n2420 ,n1450 ,n2225);
    or g869(n2419 ,n1446 ,n2289);
    or g870(n2418 ,n1500 ,n2223);
    or g871(n2417 ,n1475 ,n2288);
    or g872(n2416 ,n1619 ,n2222);
    or g873(n2415 ,n1579 ,n2287);
    or g874(n2414 ,n1662 ,n2286);
    or g875(n2413 ,n1534 ,n2066);
    or g876(n2412 ,n1682 ,n2128);
    or g877(n2411 ,n1624 ,n2126);
    or g878(n2410 ,n1665 ,n2123);
    or g879(n2409 ,n1686 ,n2119);
    or g880(n2408 ,n1531 ,n2117);
    or g881(n2407 ,n1668 ,n2114);
    or g882(n2406 ,n1632 ,n2111);
    or g883(n2405 ,n1660 ,n2108);
    or g884(n2404 ,n1651 ,n2104);
    or g885(n2403 ,n1646 ,n2102);
    or g886(n2402 ,n1643 ,n2099);
    or g887(n2401 ,n1642 ,n2096);
    or g888(n2400 ,n1640 ,n2156);
    or g889(n2399 ,n1638 ,n2092);
    or g890(n2398 ,n1634 ,n2091);
    or g891(n2397 ,n1631 ,n2155);
    or g892(n2396 ,n1628 ,n2090);
    or g893(n2395 ,n1625 ,n2154);
    or g894(n2394 ,n1621 ,n2153);
    or g895(n2393 ,n1618 ,n2089);
    or g896(n2392 ,n1615 ,n2152);
    or g897(n2391 ,n1613 ,n2151);
    or g898(n2390 ,n1611 ,n2088);
    or g899(n2389 ,n1606 ,n2087);
    or g900(n2388 ,n1603 ,n2086);
    or g901(n2387 ,n1600 ,n2085);
    or g902(n2386 ,n1596 ,n2150);
    or g903(n2385 ,n1594 ,n2149);
    or g904(n2384 ,n1592 ,n2084);
    or g905(n2383 ,n1587 ,n2148);
    or g906(n2382 ,n1584 ,n2083);
    or g907(n2381 ,n1581 ,n2082);
    or g908(n2380 ,n1578 ,n2081);
    or g909(n2379 ,n1575 ,n2080);
    or g910(n2378 ,n1573 ,n2079);
    or g911(n2377 ,n1570 ,n2078);
    or g912(n2376 ,n1568 ,n2125);
    or g913(n2375 ,n1565 ,n2076);
    or g914(n2374 ,n1562 ,n2075);
    or g915(n2373 ,n1560 ,n2074);
    or g916(n2372 ,n1557 ,n2073);
    or g917(n2371 ,n1554 ,n2072);
    or g918(n2370 ,n1551 ,n2071);
    or g919(n2369 ,n1547 ,n2070);
    or g920(n2368 ,n1544 ,n2069);
    or g921(n2367 ,n1542 ,n2068);
    or g922(n2366 ,n1538 ,n2067);
    or g923(n2365 ,n1461 ,n2157);
    or g924(n2364 ,n1530 ,n2147);
    or g925(n2363 ,n1527 ,n2146);
    or g926(n2362 ,n1525 ,n2065);
    or g927(n2361 ,n1522 ,n2064);
    or g928(n2360 ,n1518 ,n2063);
    or g929(n2359 ,n1516 ,n2062);
    or g930(n2358 ,n1513 ,n2061);
    or g931(n2357 ,n1511 ,n2060);
    or g932(n2356 ,n1507 ,n2059);
    or g933(n2355 ,n1504 ,n2145);
    or g934(n2354 ,n1502 ,n2058);
    or g935(n2353 ,n1498 ,n2144);
    or g936(n2352 ,n1496 ,n2057);
    or g937(n2351 ,n1493 ,n2056);
    or g938(n2350 ,n1454 ,n2143);
    or g939(n2349 ,n1883 ,n2141);
    or g940(n2348 ,n2028 ,n2140);
    or g941(n2347 ,n2027 ,n2139);
    or g942(n2346 ,n2026 ,n2138);
    or g943(n2345 ,n2024 ,n2137);
    or g944(n2344 ,n2023 ,n2136);
    or g945(n2343 ,n2022 ,n2135);
    or g946(n2342 ,n2021 ,n2134);
    or g947(n2341 ,n2020 ,n2133);
    or g948(n2340 ,n2018 ,n2132);
    or g949(n2339 ,n2017 ,n2131);
    or g950(n2338 ,n2016 ,n2130);
    or g951(n2337 ,n2015 ,n2129);
    or g952(n2336 ,n2013 ,n2127);
    or g953(n2335 ,n2012 ,n2077);
    or g954(n2334 ,n2011 ,n2124);
    or g955(n2333 ,n2010 ,n2122);
    or g956(n2332 ,n2019 ,n2121);
    or g957(n2331 ,n2009 ,n2120);
    or g958(n2330 ,n2008 ,n2118);
    or g959(n2329 ,n2007 ,n2116);
    or g960(n2328 ,n2006 ,n2115);
    or g961(n2327 ,n2005 ,n2113);
    or g962(n2326 ,n2004 ,n2112);
    or g963(n2325 ,n2003 ,n2110);
    or g964(n2324 ,n2002 ,n2109);
    or g965(n2323 ,n2001 ,n2107);
    or g966(n2322 ,n2000 ,n2106);
    or g967(n2321 ,n1992 ,n2105);
    or g968(n2320 ,n1999 ,n2103);
    or g969(n2319 ,n1998 ,n2101);
    or g970(n2318 ,n1997 ,n2100);
    or g971(n2317 ,n1797 ,n2205);
    or g972(n2316 ,n1995 ,n2097);
    or g973(n2315 ,n2014 ,n2095);
    or g974(n2314 ,n1994 ,n2094);
    or g975(n2313 ,n1993 ,n2093);
    or g976(n2312 ,n1991 ,n2055);
    or g977(n2311 ,n1990 ,n2054);
    or g978(n2310 ,n1989 ,n2053);
    or g979(n2309 ,n1988 ,n2052);
    or g980(n2308 ,n1987 ,n2051);
    or g981(n2307 ,n1986 ,n2050);
    or g982(n2306 ,n1985 ,n2049);
    or g983(n2305 ,n1984 ,n2048);
    or g984(n2304 ,n1983 ,n2047);
    or g985(n2303 ,n1982 ,n2046);
    or g986(n2302 ,n1981 ,n2045);
    or g987(n2301 ,n1980 ,n2044);
    or g988(n2300 ,n1979 ,n2043);
    or g989(n2299 ,n1978 ,n2042);
    or g990(n2298 ,n1977 ,n2041);
    or g991(n2297 ,n1976 ,n2040);
    or g992(n2296 ,n1975 ,n2039);
    or g993(n2295 ,n1974 ,n2038);
    or g994(n2294 ,n1973 ,n2037);
    or g995(n2293 ,n1972 ,n2036);
    or g996(n2292 ,n1971 ,n2035);
    or g997(n2291 ,n1970 ,n2034);
    or g998(n2290 ,n1969 ,n2033);
    or g999(n2289 ,n2025 ,n2032);
    or g1000(n2288 ,n1968 ,n2031);
    or g1001(n2287 ,n1967 ,n2030);
    or g1002(n2286 ,n1966 ,n2142);
    or g1003(n2285 ,n1805 ,n2218);
    or g1004(n2284 ,n1835 ,n2173);
    or g1005(n2283 ,n1832 ,n2220);
    or g1006(n2282 ,n1831 ,n2217);
    or g1007(n2281 ,n1828 ,n2219);
    or g1008(n2280 ,n1824 ,n2216);
    or g1009(n2279 ,n1822 ,n2215);
    or g1010(n2278 ,n1801 ,n2214);
    or g1011(n2277 ,n1816 ,n2213);
    or g1012(n2276 ,n1770 ,n2212);
    or g1013(n2275 ,n1807 ,n2211);
    or g1014(n2274 ,n1753 ,n2210);
    or g1015(n2273 ,n1795 ,n2209);
    or g1016(n2272 ,n1812 ,n2208);
    or g1017(n2271 ,n1799 ,n2207);
    or g1018(n2270 ,n1798 ,n2206);
    or g1019(n2269 ,n1996 ,n2098);
    or g1020(n2268 ,n1794 ,n2204);
    or g1021(n2267 ,n1790 ,n2203);
    or g1022(n2266 ,n1792 ,n2202);
    or g1023(n2265 ,n1789 ,n2201);
    or g1024(n2264 ,n1788 ,n2200);
    or g1025(n2263 ,n1786 ,n2199);
    or g1026(n2262 ,n1785 ,n2198);
    or g1027(n2261 ,n1784 ,n2197);
    or g1028(n2260 ,n1783 ,n2196);
    or g1029(n2259 ,n1782 ,n2195);
    or g1030(n2258 ,n1781 ,n2194);
    or g1031(n2257 ,n1780 ,n2193);
    or g1032(n2256 ,n1779 ,n2192);
    or g1033(n2255 ,n1777 ,n2191);
    or g1034(n2254 ,n1774 ,n2190);
    or g1035(n2253 ,n1773 ,n2189);
    or g1036(n2252 ,n1771 ,n2187);
    or g1037(n2251 ,n1772 ,n2188);
    or g1038(n2250 ,n1769 ,n2186);
    or g1039(n2249 ,n1767 ,n2185);
    or g1040(n2248 ,n1766 ,n2184);
    or g1041(n2247 ,n1764 ,n2183);
    or g1042(n2246 ,n1763 ,n2182);
    or g1043(n2245 ,n1761 ,n2181);
    or g1044(n2244 ,n1760 ,n2180);
    or g1045(n2243 ,n1759 ,n2179);
    or g1046(n2242 ,n1758 ,n2178);
    or g1047(n2241 ,n1755 ,n2177);
    or g1048(n2240 ,n1754 ,n2176);
    or g1049(n2239 ,n1752 ,n2175);
    or g1050(n2238 ,n1750 ,n2174);
    or g1051(n2237 ,n1747 ,n2221);
    or g1052(n2236 ,n1744 ,n2172);
    or g1053(n2235 ,n1742 ,n2171);
    or g1054(n2234 ,n1583 ,n2170);
    or g1055(n2233 ,n1724 ,n2169);
    or g1056(n2232 ,n1722 ,n2168);
    or g1057(n2231 ,n1720 ,n2167);
    or g1058(n2230 ,n1718 ,n2166);
    or g1059(n2229 ,n1715 ,n2165);
    or g1060(n2228 ,n1704 ,n2162);
    or g1061(n2227 ,n1712 ,n2164);
    or g1062(n2226 ,n1711 ,n2163);
    or g1063(n2225 ,n1707 ,n2161);
    or g1064(n2224 ,n1829 ,n2160);
    or g1065(n2223 ,n1703 ,n2159);
    or g1066(n2222 ,n1821 ,n2158);
    nor g1067(n2221 ,n638 ,n1735);
    nor g1068(n2220 ,n673 ,n1733);
    nor g1069(n2219 ,n681 ,n1733);
    nor g1070(n2218 ,n727 ,n1730);
    nor g1071(n2217 ,n649 ,n1730);
    nor g1072(n2216 ,n552 ,n1730);
    nor g1073(n2215 ,n709 ,n1730);
    nor g1074(n2214 ,n617 ,n1730);
    nor g1075(n2213 ,n675 ,n1730);
    nor g1076(n2212 ,n647 ,n1730);
    nor g1077(n2211 ,n628 ,n1731);
    nor g1078(n2210 ,n618 ,n1731);
    nor g1079(n2209 ,n703 ,n1731);
    nor g1080(n2208 ,n596 ,n1731);
    nor g1081(n2207 ,n598 ,n1731);
    nor g1082(n2206 ,n640 ,n1731);
    nor g1083(n2205 ,n713 ,n1731);
    nor g1084(n2204 ,n566 ,n1731);
    nor g1085(n2203 ,n563 ,n1732);
    nor g1086(n2202 ,n560 ,n1732);
    nor g1087(n2201 ,n593 ,n1732);
    nor g1088(n2200 ,n648 ,n1732);
    nor g1089(n2199 ,n733 ,n1732);
    nor g1090(n2198 ,n724 ,n1732);
    nor g1091(n2197 ,n607 ,n1732);
    nor g1092(n2196 ,n712 ,n1732);
    nor g1093(n2195 ,n627 ,n1737);
    nor g1094(n2194 ,n693 ,n1737);
    nor g1095(n2193 ,n683 ,n1737);
    nor g1096(n2192 ,n679 ,n1737);
    nor g1097(n2191 ,n650 ,n1737);
    nor g1098(n2190 ,n691 ,n1737);
    nor g1099(n2189 ,n664 ,n1737);
    nor g1100(n2188 ,n657 ,n1737);
    nor g1101(n2187 ,n653 ,n1734);
    nor g1102(n2186 ,n646 ,n1734);
    nor g1103(n2185 ,n698 ,n1734);
    nor g1104(n2184 ,n545 ,n1734);
    nor g1105(n2183 ,n685 ,n1734);
    nor g1106(n2182 ,n635 ,n1734);
    nor g1107(n2181 ,n601 ,n1734);
    nor g1108(n2180 ,n606 ,n1734);
    nor g1109(n2179 ,n599 ,n1735);
    nor g1110(n2178 ,n562 ,n1735);
    nor g1111(n2177 ,n699 ,n1735);
    nor g1112(n2176 ,n668 ,n1735);
    nor g1113(n2175 ,n642 ,n1735);
    nor g1114(n2174 ,n641 ,n1735);
    nor g1115(n2173 ,n729 ,n1733);
    nor g1116(n2172 ,n555 ,n1735);
    nor g1117(n2171 ,n626 ,n1736);
    nor g1118(n2170 ,n697 ,n1736);
    nor g1119(n2169 ,n549 ,n1736);
    nor g1120(n2168 ,n622 ,n1736);
    nor g1121(n2167 ,n717 ,n1736);
    nor g1122(n2166 ,n591 ,n1736);
    nor g1123(n2165 ,n660 ,n1736);
    nor g1124(n2164 ,n594 ,n1736);
    nor g1125(n2163 ,n623 ,n1733);
    nor g1126(n2162 ,n662 ,n1730);
    nor g1127(n2161 ,n571 ,n1733);
    nor g1128(n2160 ,n696 ,n1733);
    nor g1129(n2159 ,n694 ,n1733);
    nor g1130(n2158 ,n539 ,n1733);
    or g1131(n2157 ,n1495 ,n1954);
    or g1132(n2156 ,n1639 ,n1916);
    or g1133(n2155 ,n1629 ,n1913);
    or g1134(n2154 ,n1623 ,n1911);
    or g1135(n2153 ,n1620 ,n1910);
    or g1136(n2152 ,n1614 ,n1908);
    or g1137(n2151 ,n1612 ,n1907);
    or g1138(n2150 ,n1595 ,n1902);
    or g1139(n2149 ,n1593 ,n1901);
    or g1140(n2148 ,n1586 ,n1899);
    or g1141(n2147 ,n1528 ,n1878);
    or g1142(n2146 ,n1526 ,n1877);
    or g1143(n2145 ,n1503 ,n1869);
    or g1144(n2144 ,n1497 ,n1867);
    or g1145(n2143 ,n1489 ,n1864);
    or g1146(n2142 ,n1837 ,n1965);
    or g1147(n2141 ,n1836 ,n1964);
    or g1148(n2140 ,n1834 ,n1963);
    or g1149(n2139 ,n1775 ,n1962);
    or g1150(n2138 ,n1830 ,n1961);
    or g1151(n2137 ,n1827 ,n1960);
    or g1152(n2136 ,n1826 ,n1959);
    or g1153(n2135 ,n1706 ,n1958);
    or g1154(n2134 ,n1823 ,n1956);
    or g1155(n2133 ,n1727 ,n1955);
    or g1156(n2132 ,n1820 ,n1953);
    or g1157(n2131 ,n1756 ,n1952);
    or g1158(n2130 ,n1819 ,n1951);
    or g1159(n2129 ,n1793 ,n1949);
    or g1160(n2128 ,n1950 ,n1678);
    or g1161(n2127 ,n1818 ,n1947);
    or g1162(n2126 ,n1946 ,n1659);
    or g1163(n2125 ,n1891 ,n1566);
    or g1164(n2124 ,n1815 ,n1944);
    or g1165(n2123 ,n1943 ,n1673);
    or g1166(n2122 ,n1814 ,n1942);
    or g1167(n2121 ,n1708 ,n1941);
    or g1168(n2120 ,n1811 ,n1939);
    or g1169(n2119 ,n1940 ,n1510);
    or g1170(n2118 ,n1765 ,n1938);
    or g1171(n2117 ,n1937 ,n1607);
    or g1172(n2116 ,n1810 ,n1888);
    or g1173(n2115 ,n1809 ,n1936);
    or g1174(n2114 ,n1898 ,n1666);
    or g1175(n2113 ,n1808 ,n1934);
    or g1176(n2112 ,n1800 ,n1933);
    or g1177(n2111 ,n1932 ,n1535);
    or g1178(n2110 ,n1806 ,n1931);
    or g1179(n2109 ,n1709 ,n1930);
    or g1180(n2108 ,n1929 ,n1656);
    or g1181(n2107 ,n1804 ,n1928);
    or g1182(n2106 ,n1746 ,n1927);
    or g1183(n2105 ,n1757 ,n1926);
    or g1184(n2104 ,n1925 ,n1648);
    or g1185(n2103 ,n1762 ,n1924);
    or g1186(n2102 ,n1923 ,n1585);
    or g1187(n2101 ,n1791 ,n1922);
    or g1188(n2100 ,n1796 ,n1921);
    or g1189(n2099 ,n1919 ,n1451);
    or g1190(n2098 ,n1802 ,n1920);
    or g1191(n2097 ,n1813 ,n1935);
    or g1192(n2096 ,n1918 ,n1677);
    or g1193(n2095 ,n1825 ,n1948);
    or g1194(n2094 ,n1739 ,n1957);
    or g1195(n2093 ,n1833 ,n1917);
    or g1196(n2092 ,n1915 ,n1637);
    or g1197(n2091 ,n1914 ,n1633);
    or g1198(n2090 ,n1912 ,n1626);
    or g1199(n2089 ,n1909 ,n1617);
    or g1200(n2088 ,n1906 ,n1608);
    or g1201(n2087 ,n1905 ,n1604);
    or g1202(n2086 ,n1904 ,n1602);
    or g1203(n2085 ,n1903 ,n1599);
    or g1204(n2084 ,n1900 ,n1589);
    or g1205(n2083 ,n1897 ,n1729);
    or g1206(n2082 ,n1896 ,n1580);
    or g1207(n2081 ,n1895 ,n1577);
    or g1208(n2080 ,n1894 ,n1574);
    or g1209(n2079 ,n1893 ,n1572);
    or g1210(n2078 ,n1892 ,n1569);
    or g1211(n2077 ,n1817 ,n1945);
    or g1212(n2076 ,n1890 ,n1564);
    or g1213(n2075 ,n1889 ,n1561);
    or g1214(n2074 ,n1887 ,n1558);
    or g1215(n2073 ,n1886 ,n1555);
    or g1216(n2072 ,n1885 ,n1553);
    or g1217(n2071 ,n1884 ,n1549);
    or g1218(n2070 ,n2029 ,n1545);
    or g1219(n2069 ,n1882 ,n1543);
    or g1220(n2068 ,n1881 ,n1540);
    or g1221(n2067 ,n1880 ,n1536);
    or g1222(n2066 ,n1879 ,n1532);
    or g1223(n2065 ,n1876 ,n1523);
    or g1224(n2064 ,n1875 ,n1520);
    or g1225(n2063 ,n1874 ,n1517);
    or g1226(n2062 ,n1873 ,n1515);
    or g1227(n2061 ,n1872 ,n1512);
    or g1228(n2060 ,n1871 ,n1509);
    or g1229(n2059 ,n1870 ,n1505);
    or g1230(n2058 ,n1868 ,n1501);
    or g1231(n2057 ,n1866 ,n1494);
    or g1232(n2056 ,n1865 ,n1492);
    or g1233(n2055 ,n1751 ,n1863);
    or g1234(n2054 ,n1749 ,n1862);
    or g1235(n2053 ,n1748 ,n1861);
    or g1236(n2052 ,n1745 ,n1860);
    or g1237(n2051 ,n1743 ,n1859);
    or g1238(n2050 ,n1741 ,n1858);
    or g1239(n2049 ,n1740 ,n1857);
    or g1240(n2048 ,n1738 ,n1856);
    or g1241(n2047 ,n1728 ,n1855);
    or g1242(n2046 ,n1725 ,n1854);
    or g1243(n2045 ,n1723 ,n1853);
    or g1244(n2044 ,n1776 ,n1852);
    or g1245(n2043 ,n1721 ,n1851);
    or g1246(n2042 ,n1719 ,n1850);
    or g1247(n2041 ,n1717 ,n1849);
    or g1248(n2040 ,n1716 ,n1848);
    or g1249(n2039 ,n1714 ,n1847);
    or g1250(n2038 ,n1778 ,n1846);
    or g1251(n2037 ,n1787 ,n1845);
    or g1252(n2036 ,n1710 ,n1844);
    or g1253(n2035 ,n1768 ,n1843);
    or g1254(n2034 ,n1713 ,n1842);
    or g1255(n2033 ,n1726 ,n1841);
    or g1256(n2032 ,n1705 ,n1840);
    or g1257(n2031 ,n1803 ,n1839);
    or g1258(n2030 ,n1702 ,n1838);
    nor g1259(n2029 ,n736 ,n1226);
    nor g1260(n2028 ,n364 ,n1208);
    nor g1261(n2027 ,n455 ,n1208);
    nor g1262(n2026 ,n409 ,n1208);
    nor g1263(n2025 ,n472 ,n1219);
    nor g1264(n2024 ,n385 ,n1208);
    nor g1265(n2023 ,n456 ,n1217);
    nor g1266(n2022 ,n434 ,n1217);
    nor g1267(n2021 ,n407 ,n1217);
    nor g1268(n2020 ,n401 ,n1217);
    nor g1269(n2019 ,n405 ,n1210);
    nor g1270(n2018 ,n371 ,n1217);
    nor g1271(n2017 ,n367 ,n1217);
    nor g1272(n2016 ,n454 ,n1217);
    nor g1273(n2015 ,n362 ,n1217);
    nor g1274(n2014 ,n404 ,n1211);
    nor g1275(n2013 ,n373 ,n1210);
    nor g1276(n2012 ,n430 ,n1210);
    nor g1277(n2011 ,n374 ,n1210);
    nor g1278(n2010 ,n752 ,n1210);
    nor g1279(n2009 ,n363 ,n1210);
    nor g1280(n2008 ,n360 ,n1210);
    nor g1281(n2007 ,n749 ,n1210);
    nor g1282(n2006 ,n453 ,n1214);
    nor g1283(n2005 ,n381 ,n1214);
    nor g1284(n2004 ,n391 ,n1214);
    nor g1285(n2003 ,n390 ,n1214);
    nor g1286(n2002 ,n451 ,n1214);
    nor g1287(n2001 ,n410 ,n1214);
    nor g1288(n2000 ,n747 ,n1214);
    nor g1289(n1999 ,n408 ,n1211);
    nor g1290(n1998 ,n368 ,n1211);
    nor g1291(n1997 ,n375 ,n1211);
    nor g1292(n1996 ,n413 ,n1211);
    nor g1293(n1995 ,n389 ,n1211);
    nor g1294(n1994 ,n416 ,n1211);
    nor g1295(n1993 ,n429 ,n1211);
    nor g1296(n1992 ,n466 ,n1214);
    nor g1297(n1991 ,n402 ,n1220);
    nor g1298(n1990 ,n737 ,n1220);
    nor g1299(n1989 ,n452 ,n1220);
    nor g1300(n1988 ,n428 ,n1220);
    nor g1301(n1987 ,n411 ,n1220);
    nor g1302(n1986 ,n400 ,n1220);
    nor g1303(n1985 ,n379 ,n1220);
    nor g1304(n1984 ,n388 ,n1220);
    nor g1305(n1983 ,n739 ,n1221);
    nor g1306(n1982 ,n397 ,n1221);
    nor g1307(n1981 ,n421 ,n1221);
    nor g1308(n1980 ,n446 ,n1221);
    nor g1309(n1979 ,n743 ,n1221);
    nor g1310(n1978 ,n399 ,n1221);
    nor g1311(n1977 ,n365 ,n1221);
    nor g1312(n1976 ,n414 ,n1221);
    nor g1313(n1975 ,n465 ,n1219);
    nor g1314(n1974 ,n392 ,n1219);
    nor g1315(n1973 ,n398 ,n1219);
    nor g1316(n1972 ,n396 ,n1219);
    nor g1317(n1971 ,n461 ,n1219);
    nor g1318(n1970 ,n369 ,n1219);
    nor g1319(n1969 ,n382 ,n1219);
    nor g1320(n1968 ,n386 ,n1208);
    nor g1321(n1967 ,n463 ,n1208);
    nor g1322(n1966 ,n380 ,n1208);
    nor g1323(n1965 ,n582 ,n1222);
    nor g1324(n1964 ,n680 ,n1222);
    nor g1325(n1963 ,n701 ,n1222);
    nor g1326(n1962 ,n575 ,n1222);
    nor g1327(n1961 ,n636 ,n1222);
    nor g1328(n1960 ,n719 ,n1222);
    nor g1329(n1959 ,n605 ,n1231);
    nor g1330(n1958 ,n541 ,n1231);
    nor g1331(n1957 ,n612 ,n1224);
    nor g1332(n1956 ,n715 ,n1231);
    nor g1333(n1955 ,n665 ,n1231);
    nor g1334(n1954 ,n629 ,n1213);
    nor g1335(n1953 ,n687 ,n1231);
    nor g1336(n1952 ,n711 ,n1231);
    nor g1337(n1951 ,n588 ,n1231);
    nor g1338(n1950 ,n721 ,n1213);
    nor g1339(n1949 ,n716 ,n1231);
    nor g1340(n1948 ,n718 ,n1224);
    nor g1341(n1947 ,n587 ,n1225);
    nor g1342(n1946 ,n631 ,n1213);
    nor g1343(n1945 ,n602 ,n1225);
    nor g1344(n1944 ,n730 ,n1225);
    nor g1345(n1943 ,n565 ,n1213);
    nor g1346(n1942 ,n655 ,n1225);
    nor g1347(n1941 ,n568 ,n1225);
    nor g1348(n1940 ,n573 ,n1213);
    nor g1349(n1939 ,n684 ,n1225);
    nor g1350(n1938 ,n674 ,n1225);
    nor g1351(n1937 ,n700 ,n1213);
    nor g1352(n1936 ,n654 ,n1223);
    nor g1353(n1935 ,n645 ,n1224);
    nor g1354(n1934 ,n706 ,n1223);
    nor g1355(n1933 ,n630 ,n1223);
    nor g1356(n1932 ,n544 ,n1213);
    nor g1357(n1931 ,n619 ,n1223);
    nor g1358(n1930 ,n624 ,n1223);
    nor g1359(n1929 ,n558 ,n1216);
    nor g1360(n1928 ,n720 ,n1223);
    nor g1361(n1927 ,n678 ,n1223);
    nor g1362(n1926 ,n580 ,n1223);
    nor g1363(n1925 ,n548 ,n1216);
    nor g1364(n1924 ,n633 ,n1224);
    nor g1365(n1923 ,n600 ,n1216);
    nor g1366(n1922 ,n656 ,n1224);
    nor g1367(n1921 ,n669 ,n1224);
    nor g1368(n1920 ,n584 ,n1224);
    nor g1369(n1919 ,n604 ,n1216);
    nor g1370(n1918 ,n570 ,n1216);
    nor g1371(n1917 ,n722 ,n1224);
    nor g1372(n1916 ,n731 ,n1216);
    nor g1373(n1915 ,n652 ,n1216);
    nor g1374(n1914 ,n610 ,n1216);
    nor g1375(n1913 ,n603 ,n1227);
    nor g1376(n1912 ,n611 ,n1227);
    nor g1377(n1911 ,n643 ,n1227);
    nor g1378(n1910 ,n577 ,n1227);
    nor g1379(n1909 ,n553 ,n1227);
    nor g1380(n1908 ,n615 ,n1227);
    nor g1381(n1907 ,n616 ,n1227);
    nor g1382(n1906 ,n677 ,n1227);
    nor g1383(n1905 ,n734 ,n1228);
    nor g1384(n1904 ,n634 ,n1228);
    nor g1385(n1903 ,n621 ,n1228);
    nor g1386(n1902 ,n707 ,n1228);
    nor g1387(n1901 ,n726 ,n1228);
    nor g1388(n1900 ,n714 ,n1228);
    nor g1389(n1899 ,n557 ,n1228);
    nor g1390(n1898 ,n735 ,n1213);
    nor g1391(n1897 ,n659 ,n1228);
    nor g1392(n1896 ,n589 ,n1230);
    nor g1393(n1895 ,n609 ,n1230);
    nor g1394(n1894 ,n578 ,n1230);
    nor g1395(n1893 ,n540 ,n1230);
    nor g1396(n1892 ,n723 ,n1230);
    nor g1397(n1891 ,n690 ,n1230);
    nor g1398(n1890 ,n579 ,n1230);
    nor g1399(n1889 ,n688 ,n1230);
    nor g1400(n1888 ,n686 ,n1225);
    nor g1401(n1887 ,n581 ,n1226);
    nor g1402(n1886 ,n661 ,n1226);
    nor g1403(n1885 ,n682 ,n1226);
    nor g1404(n1884 ,n702 ,n1226);
    nor g1405(n1883 ,n403 ,n1208);
    nor g1406(n1882 ,n546 ,n1226);
    nor g1407(n1881 ,n608 ,n1226);
    nor g1408(n1880 ,n672 ,n1226);
    nor g1409(n1879 ,n576 ,n1229);
    nor g1410(n1878 ,n556 ,n1229);
    nor g1411(n1877 ,n644 ,n1229);
    nor g1412(n1876 ,n705 ,n1229);
    nor g1413(n1875 ,n639 ,n1229);
    nor g1414(n1874 ,n663 ,n1229);
    nor g1415(n1873 ,n689 ,n1229);
    nor g1416(n1872 ,n695 ,n1229);
    nor g1417(n1871 ,n572 ,n1209);
    nor g1418(n1870 ,n559 ,n1209);
    nor g1419(n1869 ,n567 ,n1209);
    nor g1420(n1868 ,n658 ,n1209);
    nor g1421(n1867 ,n676 ,n1209);
    nor g1422(n1866 ,n614 ,n1209);
    nor g1423(n1865 ,n569 ,n1209);
    nor g1424(n1864 ,n590 ,n1209);
    nor g1425(n1863 ,n551 ,n1218);
    nor g1426(n1862 ,n732 ,n1218);
    nor g1427(n1861 ,n670 ,n1218);
    nor g1428(n1860 ,n574 ,n1218);
    nor g1429(n1859 ,n710 ,n1218);
    nor g1430(n1858 ,n632 ,n1218);
    nor g1431(n1857 ,n667 ,n1218);
    nor g1432(n1856 ,n595 ,n1218);
    nor g1433(n1855 ,n625 ,n1212);
    nor g1434(n1854 ,n637 ,n1212);
    nor g1435(n1853 ,n725 ,n1212);
    nor g1436(n1852 ,n583 ,n1212);
    nor g1437(n1851 ,n585 ,n1212);
    nor g1438(n1850 ,n728 ,n1212);
    nor g1439(n1849 ,n671 ,n1212);
    nor g1440(n1848 ,n692 ,n1212);
    nor g1441(n1847 ,n651 ,n1215);
    nor g1442(n1846 ,n592 ,n1215);
    nor g1443(n1845 ,n708 ,n1215);
    nor g1444(n1844 ,n597 ,n1215);
    nor g1445(n1843 ,n620 ,n1215);
    nor g1446(n1842 ,n536 ,n1215);
    nor g1447(n1841 ,n550 ,n1215);
    nor g1448(n1840 ,n613 ,n1215);
    nor g1449(n1839 ,n586 ,n1222);
    nor g1450(n1838 ,n666 ,n1222);
    nor g1451(n1837 ,n2[90] ,n1440);
    nor g1452(n1836 ,n2[91] ,n1440);
    nor g1453(n1835 ,n5[61] ,n1441);
    nor g1454(n1834 ,n2[92] ,n1440);
    nor g1455(n1833 ,n2[127] ,n1436);
    nor g1456(n1832 ,n5[62] ,n1441);
    nor g1457(n1831 ,n5[2] ,n1439);
    nor g1458(n1830 ,n2[94] ,n1440);
    nor g1459(n1829 ,n5[58] ,n1441);
    nor g1460(n1828 ,n5[63] ,n1441);
    nor g1461(n1827 ,n2[95] ,n1440);
    nor g1462(n1826 ,n2[96] ,n1433);
    nor g1463(n1825 ,n2[125] ,n1436);
    nor g1464(n1824 ,n5[3] ,n1439);
    nor g1465(n1823 ,n2[98] ,n1433);
    nor g1466(n1822 ,n5[4] ,n1439);
    nor g1467(n1821 ,n5[60] ,n1441);
    nor g1468(n1820 ,n2[100] ,n1433);
    nor g1469(n1819 ,n2[102] ,n1433);
    nor g1470(n1818 ,n2[104] ,n1435);
    nor g1471(n1817 ,n2[105] ,n1435);
    nor g1472(n1816 ,n5[6] ,n1439);
    nor g1473(n1815 ,n2[106] ,n1435);
    nor g1474(n1814 ,n2[107] ,n1435);
    nor g1475(n1813 ,n2[124] ,n1436);
    nor g1476(n1812 ,n5[11] ,n1442);
    nor g1477(n1811 ,n2[109] ,n1435);
    nor g1478(n1810 ,n2[111] ,n1435);
    nor g1479(n1809 ,n2[112] ,n1434);
    nor g1480(n1808 ,n2[113] ,n1434);
    nor g1481(n1807 ,n5[8] ,n1442);
    nor g1482(n1806 ,n2[115] ,n1434);
    nor g1483(n1805 ,n5[1] ,n1439);
    nor g1484(n1804 ,n2[117] ,n1434);
    nor g1485(n1803 ,n2[88] ,n1440);
    nor g1486(n1802 ,n2[123] ,n1436);
    nor g1487(n1801 ,n5[5] ,n1439);
    nor g1488(n1800 ,n2[114] ,n1434);
    nor g1489(n1799 ,n5[12] ,n1442);
    nor g1490(n1798 ,n5[13] ,n1442);
    nor g1491(n1797 ,n5[14] ,n1442);
    nor g1492(n1796 ,n2[122] ,n1436);
    nor g1493(n1795 ,n5[10] ,n1442);
    nor g1494(n1794 ,n5[15] ,n1442);
    nor g1495(n1793 ,n2[103] ,n1433);
    nor g1496(n1792 ,n5[17] ,n1443);
    nor g1497(n1791 ,n2[121] ,n1436);
    nor g1498(n1790 ,n5[16] ,n1443);
    nor g1499(n1789 ,n5[18] ,n1443);
    nor g1500(n1788 ,n5[19] ,n1443);
    nor g1501(n1787 ,n2[82] ,n1437);
    nor g1502(n1786 ,n5[20] ,n1443);
    nor g1503(n1785 ,n5[21] ,n1443);
    nor g1504(n1784 ,n5[22] ,n1443);
    nor g1505(n1783 ,n5[23] ,n1443);
    nor g1506(n1782 ,n5[24] ,n1444);
    nor g1507(n1781 ,n5[25] ,n1444);
    nor g1508(n1780 ,n5[26] ,n1444);
    nor g1509(n1779 ,n5[27] ,n1444);
    nor g1510(n1778 ,n2[81] ,n1437);
    nor g1511(n1777 ,n5[28] ,n1444);
    nor g1512(n1776 ,n2[75] ,n1432);
    nor g1513(n1775 ,n2[93] ,n1440);
    nor g1514(n1774 ,n5[29] ,n1444);
    nor g1515(n1773 ,n5[30] ,n1444);
    nor g1516(n1772 ,n5[31] ,n1444);
    nor g1517(n1771 ,n5[32] ,n1445);
    nor g1518(n1770 ,n5[7] ,n1439);
    nor g1519(n1769 ,n5[33] ,n1445);
    nor g1520(n1768 ,n2[84] ,n1437);
    nor g1521(n1767 ,n5[34] ,n1445);
    nor g1522(n1766 ,n5[35] ,n1445);
    nor g1523(n1765 ,n2[110] ,n1435);
    nor g1524(n1764 ,n5[36] ,n1445);
    nor g1525(n1763 ,n5[37] ,n1445);
    nor g1526(n1762 ,n2[120] ,n1436);
    nor g1527(n1761 ,n5[38] ,n1445);
    nor g1528(n1760 ,n5[39] ,n1445);
    nor g1529(n1759 ,n5[40] ,n1430);
    nor g1530(n1758 ,n5[41] ,n1430);
    nor g1531(n1757 ,n2[119] ,n1434);
    nor g1532(n1756 ,n2[101] ,n1433);
    nor g1533(n1755 ,n5[42] ,n1430);
    nor g1534(n1754 ,n5[43] ,n1430);
    nor g1535(n1753 ,n5[9] ,n1442);
    nor g1536(n1752 ,n5[44] ,n1430);
    nor g1537(n1751 ,n2[64] ,n1438);
    nor g1538(n1750 ,n5[45] ,n1430);
    nor g1539(n1749 ,n2[65] ,n1438);
    nor g1540(n1748 ,n2[66] ,n1438);
    nor g1541(n1747 ,n5[46] ,n1430);
    nor g1542(n1746 ,n2[118] ,n1434);
    nor g1543(n1745 ,n2[67] ,n1438);
    nor g1544(n1744 ,n5[47] ,n1430);
    nor g1545(n1743 ,n2[68] ,n1438);
    nor g1546(n1742 ,n5[48] ,n1431);
    nor g1547(n1741 ,n2[69] ,n1438);
    nor g1548(n1740 ,n2[70] ,n1438);
    nor g1549(n1739 ,n2[126] ,n1436);
    nor g1550(n1738 ,n2[71] ,n1438);
    nor g1551(n1729 ,n1030 ,n1330);
    nor g1552(n1728 ,n2[72] ,n1432);
    nor g1553(n1727 ,n2[99] ,n1433);
    nor g1554(n1726 ,n2[86] ,n1437);
    nor g1555(n1725 ,n2[73] ,n1432);
    nor g1556(n1724 ,n5[50] ,n1431);
    nor g1557(n1723 ,n2[74] ,n1432);
    nor g1558(n1722 ,n5[51] ,n1431);
    nor g1559(n1721 ,n2[76] ,n1432);
    nor g1560(n1720 ,n5[52] ,n1431);
    nor g1561(n1719 ,n2[77] ,n1432);
    nor g1562(n1718 ,n5[53] ,n1431);
    nor g1563(n1717 ,n2[78] ,n1432);
    nor g1564(n1716 ,n2[79] ,n1432);
    nor g1565(n1715 ,n5[54] ,n1431);
    nor g1566(n1714 ,n2[80] ,n1437);
    nor g1567(n1713 ,n2[85] ,n1437);
    nor g1568(n1712 ,n5[55] ,n1431);
    nor g1569(n1711 ,n5[56] ,n1441);
    nor g1570(n1710 ,n2[83] ,n1437);
    nor g1571(n1709 ,n2[116] ,n1434);
    nor g1572(n1708 ,n2[108] ,n1435);
    nor g1573(n1707 ,n5[57] ,n1441);
    nor g1574(n1706 ,n2[97] ,n1433);
    nor g1575(n1705 ,n2[87] ,n1437);
    nor g1576(n1704 ,n5[0] ,n1439);
    nor g1577(n1703 ,n5[59] ,n1441);
    nor g1578(n1702 ,n2[89] ,n1440);
    or g1579(n1701 ,n1251 ,n1397);
    or g1580(n1700 ,n1282 ,n1372);
    or g1581(n1699 ,n831 ,n1067);
    or g1582(n1698 ,n864 ,n1122);
    or g1583(n1697 ,n887 ,n1195);
    or g1584(n1696 ,n870 ,n1181);
    or g1585(n1695 ,n947 ,n1158);
    or g1586(n1694 ,n1277 ,n1426);
    or g1587(n1693 ,n946 ,n1164);
    or g1588(n1692 ,n1279 ,n1421);
    or g1589(n1691 ,n1271 ,n1382);
    or g1590(n1690 ,n945 ,n1198);
    or g1591(n1689 ,n943 ,n1068);
    or g1592(n1688 ,n915 ,n1192);
    or g1593(n1687 ,n828 ,n1194);
    or g1594(n1686 ,n929 ,n1129);
    or g1595(n1685 ,n821 ,n1090);
    or g1596(n1684 ,n853 ,n1180);
    or g1597(n1683 ,n931 ,n1150);
    or g1598(n1682 ,n936 ,n1131);
    or g1599(n1681 ,n923 ,n1133);
    or g1600(n1680 ,n1281 ,n1425);
    or g1601(n1679 ,n890 ,n1126);
    nor g1602(n1678 ,n1031 ,n1342);
    nor g1603(n1677 ,n1052 ,n1347);
    or g1604(n1676 ,n917 ,n1185);
    or g1605(n1675 ,n930 ,n1184);
    or g1606(n1674 ,n924 ,n1182);
    nor g1607(n1673 ,n1061 ,n1345);
    or g1608(n1672 ,n842 ,n1097);
    or g1609(n1671 ,n818 ,n1178);
    or g1610(n1670 ,n858 ,n1124);
    or g1611(n1669 ,n1240 ,n1422);
    or g1612(n1668 ,n862 ,n1136);
    or g1613(n1667 ,n886 ,n1142);
    nor g1614(n1666 ,n1037 ,n1343);
    or g1615(n1665 ,n926 ,n1179);
    or g1616(n1664 ,n902 ,n1152);
    or g1617(n1663 ,n834 ,n1167);
    or g1618(n1662 ,n938 ,n1189);
    or g1619(n1661 ,n941 ,n1154);
    or g1620(n1660 ,n844 ,n1066);
    nor g1621(n1659 ,n1047 ,n1346);
    or g1622(n1658 ,n869 ,n1078);
    or g1623(n1657 ,n1269 ,n1359);
    nor g1624(n1656 ,n1036 ,n1332);
    or g1625(n1655 ,n920 ,n1076);
    or g1626(n1654 ,n944 ,n1165);
    or g1627(n1653 ,n868 ,n1168);
    or g1628(n1652 ,n827 ,n1085);
    or g1629(n1651 ,n840 ,n1102);
    or g1630(n1650 ,n1274 ,n1419);
    or g1631(n1649 ,n817 ,n1084);
    nor g1632(n1648 ,n1043 ,n1341);
    or g1633(n1647 ,n1292 ,n1393);
    or g1634(n1646 ,n860 ,n1079);
    or g1635(n1645 ,n933 ,n1172);
    or g1636(n1644 ,n932 ,n1170);
    or g1637(n1643 ,n912 ,n1166);
    or g1638(n1642 ,n850 ,n1175);
    or g1639(n1641 ,n1206 ,n1418);
    or g1640(n1640 ,n1266 ,n1389);
    or g1641(n1639 ,n909 ,n1161);
    or g1642(n1638 ,n907 ,n1160);
    nor g1643(n1637 ,n1042 ,n1340);
    or g1644(n1636 ,n1257 ,n1356);
    or g1645(n1635 ,n1264 ,n1414);
    or g1646(n1634 ,n905 ,n1159);
    nor g1647(n1633 ,n1041 ,n1339);
    or g1648(n1632 ,n916 ,n1174);
    or g1649(n1631 ,n1262 ,n1413);
    or g1650(n1630 ,n1263 ,n1412);
    or g1651(n1629 ,n904 ,n1157);
    or g1652(n1628 ,n903 ,n1156);
    or g1653(n1627 ,n1261 ,n1411);
    nor g1654(n1626 ,n1039 ,n1338);
    or g1655(n1625 ,n1260 ,n1410);
    or g1656(n1624 ,n839 ,n1186);
    or g1657(n1623 ,n863 ,n1153);
    or g1658(n1622 ,n1259 ,n1409);
    or g1659(n1621 ,n1258 ,n1408);
    or g1660(n1620 ,n900 ,n1151);
    or g1661(n1619 ,n1273 ,n1423);
    or g1662(n1618 ,n899 ,n1148);
    nor g1663(n1617 ,n1027 ,n1337);
    or g1664(n1616 ,n1254 ,n1406);
    or g1665(n1615 ,n1255 ,n1407);
    or g1666(n1614 ,n882 ,n1147);
    or g1667(n1613 ,n1253 ,n1405);
    or g1668(n1612 ,n895 ,n1145);
    or g1669(n1611 ,n894 ,n1144);
    or g1670(n1610 ,n891 ,n1146);
    or g1671(n1609 ,n1250 ,n1404);
    nor g1672(n1608 ,n1035 ,n1336);
    nor g1673(n1607 ,n1040 ,n1320);
    or g1674(n1606 ,n892 ,n1143);
    or g1675(n1605 ,n1249 ,n1403);
    nor g1676(n1604 ,n1033 ,n1335);
    or g1677(n1603 ,n906 ,n1141);
    nor g1678(n1602 ,n1032 ,n1334);
    or g1679(n1601 ,n884 ,n1171);
    or g1680(n1600 ,n889 ,n1163);
    nor g1681(n1599 ,n1048 ,n1333);
    or g1682(n1598 ,n1248 ,n1402);
    or g1683(n1597 ,n1246 ,n1400);
    or g1684(n1596 ,n1247 ,n1417);
    or g1685(n1595 ,n819 ,n1140);
    or g1686(n1594 ,n1270 ,n1399);
    or g1687(n1593 ,n885 ,n1139);
    or g1688(n1592 ,n883 ,n1138);
    or g1689(n1591 ,n1244 ,n1398);
    or g1690(n1590 ,n1245 ,n1401);
    nor g1691(n1589 ,n1056 ,n1331);
    or g1692(n1588 ,n1276 ,n1395);
    or g1693(n1587 ,n1243 ,n1396);
    or g1694(n1586 ,n939 ,n1188);
    nor g1695(n1585 ,n1060 ,n1301);
    or g1696(n1584 ,n942 ,n1137);
    nor g1697(n1583 ,n5[49] ,n1431);
    or g1698(n1582 ,n1239 ,n1394);
    or g1699(n1581 ,n872 ,n1135);
    nor g1700(n1580 ,n1028 ,n1329);
    or g1701(n1579 ,n927 ,n1064);
    or g1702(n1578 ,n820 ,n1134);
    nor g1703(n1577 ,n1025 ,n1328);
    or g1704(n1576 ,n1238 ,n1391);
    or g1705(n1575 ,n822 ,n1077);
    nor g1706(n1574 ,n1024 ,n1327);
    or g1707(n1573 ,n825 ,n1132);
    nor g1708(n1572 ,n1023 ,n1326);
    or g1709(n1571 ,n1297 ,n1390);
    or g1710(n1570 ,n837 ,n1130);
    nor g1711(n1569 ,n1022 ,n1325);
    or g1712(n1568 ,n851 ,n1128);
    or g1713(n1567 ,n1234 ,n1388);
    nor g1714(n1566 ,n1021 ,n1324);
    or g1715(n1565 ,n867 ,n1127);
    nor g1716(n1564 ,n1020 ,n1323);
    or g1717(n1563 ,n1256 ,n1387);
    or g1718(n1562 ,n865 ,n1125);
    nor g1719(n1561 ,n1019 ,n1322);
    or g1720(n1560 ,n866 ,n1123);
    or g1721(n1559 ,n1233 ,n1386);
    nor g1722(n1558 ,n1018 ,n1321);
    or g1723(n1557 ,n861 ,n1121);
    or g1724(n1556 ,n1272 ,n1385);
    nor g1725(n1555 ,n1055 ,n1319);
    or g1726(n1554 ,n859 ,n1120);
    nor g1727(n1553 ,n1016 ,n1318);
    or g1728(n1552 ,n913 ,n1176);
    or g1729(n1551 ,n857 ,n1193);
    or g1730(n1550 ,n1280 ,n1384);
    nor g1731(n1549 ,n1015 ,n1317);
    or g1732(n1548 ,n1237 ,n1416);
    or g1733(n1547 ,n855 ,n1119);
    or g1734(n1546 ,n1232 ,n1383);
    nor g1735(n1545 ,n1117 ,n1316);
    or g1736(n1544 ,n854 ,n1118);
    nor g1737(n1543 ,n1014 ,n1315);
    or g1738(n1542 ,n852 ,n1116);
    or g1739(n1541 ,n1201 ,n1353);
    nor g1740(n1540 ,n1029 ,n1314);
    or g1741(n1539 ,n1283 ,n1378);
    or g1742(n1538 ,n893 ,n1114);
    or g1743(n1537 ,n1236 ,n1424);
    nor g1744(n1536 ,n1050 ,n1313);
    nor g1745(n1535 ,n1173 ,n1311);
    or g1746(n1534 ,n832 ,n1113);
    or g1747(n1533 ,n1284 ,n1381);
    nor g1748(n1532 ,n1017 ,n1312);
    or g1749(n1531 ,n928 ,n1106);
    or g1750(n1530 ,n1235 ,n1392);
    or g1751(n1529 ,n1286 ,n1379);
    or g1752(n1528 ,n881 ,n1112);
    or g1753(n1527 ,n1252 ,n1380);
    or g1754(n1526 ,n914 ,n1111);
    or g1755(n1525 ,n908 ,n1110);
    or g1756(n1524 ,n1268 ,n1377);
    nor g1757(n1523 ,n1046 ,n1310);
    or g1758(n1522 ,n919 ,n1109);
    or g1759(n1521 ,n813 ,n1196);
    nor g1760(n1520 ,n1044 ,n1309);
    or g1761(n1519 ,n1287 ,n1376);
    or g1762(n1518 ,n925 ,n1108);
    nor g1763(n1517 ,n1045 ,n1308);
    or g1764(n1516 ,n849 ,n1107);
    nor g1765(n1515 ,n1057 ,n1307);
    or g1766(n1514 ,n1288 ,n1420);
    or g1767(n1513 ,n911 ,n1104);
    nor g1768(n1512 ,n1062 ,n1306);
    or g1769(n1511 ,n847 ,n1103);
    nor g1770(n1510 ,n1099 ,n1344);
    nor g1771(n1509 ,n1081 ,n1300);
    or g1772(n1508 ,n1290 ,n1375);
    or g1773(n1507 ,n845 ,n1101);
    or g1774(n1506 ,n1291 ,n1374);
    nor g1775(n1505 ,n1089 ,n1305);
    or g1776(n1504 ,n1289 ,n1373);
    or g1777(n1503 ,n843 ,n1100);
    or g1778(n1502 ,n948 ,n1207);
    nor g1779(n1501 ,n1053 ,n1304);
    or g1780(n1500 ,n1267 ,n1348);
    or g1781(n1499 ,n1294 ,n1370);
    or g1782(n1498 ,n1293 ,n1371);
    or g1783(n1497 ,n871 ,n1187);
    or g1784(n1496 ,n937 ,n1096);
    or g1785(n1495 ,n888 ,n1190);
    nor g1786(n1494 ,n1092 ,n1303);
    or g1787(n1493 ,n838 ,n1093);
    nor g1788(n1492 ,n1162 ,n1302);
    or g1789(n1491 ,n1296 ,n1369);
    or g1790(n1490 ,n1295 ,n1367);
    or g1791(n1489 ,n835 ,n1074);
    or g1792(n1488 ,n833 ,n1115);
    or g1793(n1487 ,n1275 ,n1366);
    or g1794(n1486 ,n1298 ,n1365);
    or g1795(n1485 ,n823 ,n1088);
    or g1796(n1484 ,n829 ,n1087);
    or g1797(n1483 ,n826 ,n1091);
    or g1798(n1482 ,n1265 ,n1415);
    or g1799(n1481 ,n1428 ,n1363);
    or g1800(n1480 ,n934 ,n1177);
    or g1801(n1479 ,n824 ,n1183);
    or g1802(n1478 ,n1429 ,n1362);
    or g1803(n1477 ,n940 ,n1083);
    or g1804(n1476 ,n856 ,n1094);
    or g1805(n1475 ,n841 ,n1169);
    or g1806(n1474 ,n1098 ,n1361);
    or g1807(n1473 ,n898 ,n1082);
    or g1808(n1472 ,n1427 ,n1360);
    or g1809(n1471 ,n816 ,n1080);
    or g1810(n1470 ,n836 ,n1095);
    or g1811(n1469 ,n1285 ,n1358);
    or g1812(n1468 ,n846 ,n1075);
    or g1813(n1467 ,n1242 ,n1357);
    or g1814(n1466 ,n897 ,n1073);
    or g1815(n1465 ,n901 ,n1072);
    or g1816(n1464 ,n1278 ,n1364);
    or g1817(n1463 ,n935 ,n1191);
    or g1818(n1462 ,n815 ,n1071);
    or g1819(n1461 ,n1204 ,n1355);
    or g1820(n1460 ,n918 ,n1070);
    or g1821(n1459 ,n1203 ,n1352);
    or g1822(n1458 ,n848 ,n1069);
    or g1823(n1457 ,n1205 ,n1354);
    or g1824(n1456 ,n921 ,n1149);
    or g1825(n1455 ,n1200 ,n1351);
    or g1826(n1454 ,n1202 ,n1368);
    or g1827(n1453 ,n910 ,n1155);
    or g1828(n1452 ,n922 ,n1197);
    nor g1829(n1451 ,n1105 ,n1299);
    or g1830(n1450 ,n1199 ,n1350);
    or g1831(n1449 ,n814 ,n1063);
    or g1832(n1448 ,n830 ,n1086);
    or g1833(n1447 ,n1241 ,n1349);
    or g1834(n1446 ,n896 ,n1065);
    nor g1835(n1737 ,n878 ,n1026);
    nor g1836(n1736 ,n878 ,n1054);
    nor g1837(n1735 ,n878 ,n1049);
    nor g1838(n1734 ,n878 ,n1034);
    nor g1839(n1733 ,n878 ,n1058);
    nor g1840(n1732 ,n878 ,n1038);
    nor g1841(n1731 ,n878 ,n1059);
    nor g1842(n1730 ,n878 ,n1051);
    nor g1843(n1429 ,n3072 ,n1012);
    nor g1844(n1428 ,n3071 ,n1013);
    nor g1845(n1427 ,n3074 ,n1012);
    nor g1846(n1426 ,n313 ,n959);
    nor g1847(n1425 ,n308 ,n965);
    nor g1848(n1424 ,n330 ,n968);
    nor g1849(n1423 ,n542 ,n968);
    nor g1850(n1422 ,n346 ,n959);
    nor g1851(n1421 ,n333 ,n965);
    nor g1852(n1420 ,n554 ,n971);
    nor g1853(n1419 ,n307 ,n965);
    nor g1854(n1418 ,n335 ,n972);
    nor g1855(n1417 ,n431 ,n960);
    nor g1856(n1416 ,n324 ,n965);
    nor g1857(n1415 ,n304 ,n953);
    nor g1858(n1414 ,n352 ,n959);
    nor g1859(n1413 ,n469 ,n963);
    nor g1860(n1412 ,n321 ,n959);
    nor g1861(n1411 ,n316 ,n959);
    nor g1862(n1410 ,n440 ,n963);
    nor g1863(n1409 ,n704 ,n962);
    nor g1864(n1408 ,n422 ,n963);
    nor g1865(n1407 ,n433 ,n963);
    nor g1866(n1406 ,n354 ,n962);
    nor g1867(n1405 ,n756 ,n963);
    nor g1868(n1404 ,n344 ,n962);
    nor g1869(n1403 ,n357 ,n962);
    nor g1870(n1402 ,n305 ,n962);
    nor g1871(n1401 ,n331 ,n968);
    nor g1872(n1400 ,n334 ,n962);
    nor g1873(n1399 ,n427 ,n960);
    nor g1874(n1398 ,n306 ,n962);
    nor g1875(n1397 ,n350 ,n965);
    nor g1876(n1396 ,n393 ,n960);
    nor g1877(n1395 ,n547 ,n962);
    nor g1878(n1394 ,n543 ,n958);
    nor g1879(n1393 ,n318 ,n959);
    nor g1880(n1392 ,n361 ,n954);
    nor g1881(n1391 ,n342 ,n958);
    nor g1882(n1390 ,n353 ,n958);
    nor g1883(n1389 ,n376 ,n990);
    nor g1884(n1388 ,n358 ,n958);
    nor g1885(n1387 ,n340 ,n958);
    nor g1886(n1386 ,n319 ,n958);
    nor g1887(n1385 ,n338 ,n958);
    nor g1888(n1384 ,n317 ,n958);
    nor g1889(n1383 ,n314 ,n971);
    nor g1890(n1382 ,n332 ,n965);
    nor g1891(n1381 ,n327 ,n971);
    nor g1892(n1380 ,n432 ,n954);
    nor g1893(n1379 ,n325 ,n971);
    nor g1894(n1378 ,n351 ,n971);
    nor g1895(n1377 ,n322 ,n971);
    nor g1896(n1376 ,n356 ,n971);
    nor g1897(n1375 ,n359 ,n971);
    nor g1898(n1374 ,n337 ,n953);
    nor g1899(n1373 ,n412 ,n966);
    nor g1900(n1372 ,n538 ,n968);
    nor g1901(n1371 ,n464 ,n966);
    nor g1902(n1370 ,n310 ,n953);
    nor g1903(n1369 ,n345 ,n953);
    nor g1904(n1368 ,n419 ,n966);
    nor g1905(n1367 ,n343 ,n953);
    nor g1906(n1366 ,n326 ,n953);
    nor g1907(n1365 ,n336 ,n953);
    nor g1908(n1364 ,n349 ,n965);
    nor g1909(n1363 ,n537 ,n953);
    nor g1910(n1362 ,n320 ,n972);
    nor g1911(n1361 ,n312 ,n972);
    nor g1912(n1360 ,n347 ,n972);
    nor g1913(n1359 ,n315 ,n959);
    nor g1914(n1358 ,n323 ,n972);
    nor g1915(n1357 ,n328 ,n972);
    nor g1916(n1356 ,n311 ,n959);
    nor g1917(n1355 ,n439 ,n969);
    nor g1918(n1354 ,n341 ,n972);
    nor g1919(n1353 ,n348 ,n965);
    nor g1920(n1352 ,n309 ,n972);
    nor g1921(n1351 ,n564 ,n968);
    nor g1922(n1350 ,n355 ,n968);
    nor g1923(n1349 ,n329 ,n968);
    nor g1924(n1348 ,n339 ,n968);
    nor g1925(n1347 ,n370 ,n991);
    nor g1926(n1346 ,n751 ,n970);
    nor g1927(n1345 ,n746 ,n970);
    nor g1928(n1344 ,n417 ,n970);
    nor g1929(n1343 ,n441 ,n970);
    nor g1930(n1342 ,n448 ,n970);
    nor g1931(n1341 ,n740 ,n991);
    nor g1932(n1340 ,n387 ,n991);
    nor g1933(n1339 ,n754 ,n991);
    nor g1934(n1338 ,n435 ,n964);
    nor g1935(n1337 ,n418 ,n964);
    nor g1936(n1336 ,n366 ,n964);
    nor g1937(n1335 ,n444 ,n961);
    nor g1938(n1334 ,n750 ,n961);
    nor g1939(n1333 ,n755 ,n961);
    nor g1940(n1332 ,n449 ,n991);
    nor g1941(n1331 ,n471 ,n961);
    nor g1942(n1330 ,n460 ,n961);
    nor g1943(n1329 ,n450 ,n957);
    nor g1944(n1328 ,n457 ,n957);
    nor g1945(n1327 ,n437 ,n957);
    nor g1946(n1326 ,n468 ,n957);
    nor g1947(n1325 ,n394 ,n957);
    nor g1948(n1324 ,n425 ,n957);
    nor g1949(n1323 ,n462 ,n957);
    nor g1950(n1322 ,n420 ,n957);
    nor g1951(n1321 ,n378 ,n956);
    nor g1952(n1320 ,n395 ,n970);
    nor g1953(n1319 ,n406 ,n956);
    nor g1954(n1318 ,n423 ,n956);
    nor g1955(n1317 ,n377 ,n956);
    nor g1956(n1316 ,n384 ,n956);
    nor g1957(n1315 ,n438 ,n956);
    nor g1958(n1314 ,n474 ,n956);
    nor g1959(n1313 ,n415 ,n956);
    nor g1960(n1312 ,n436 ,n955);
    nor g1961(n1311 ,n467 ,n970);
    nor g1962(n1310 ,n383 ,n955);
    nor g1963(n1309 ,n458 ,n955);
    nor g1964(n1308 ,n447 ,n955);
    nor g1965(n1307 ,n459 ,n955);
    nor g1966(n1306 ,n445 ,n955);
    nor g1967(n1305 ,n424 ,n967);
    nor g1968(n1304 ,n470 ,n967);
    nor g1969(n1303 ,n473 ,n967);
    nor g1970(n1302 ,n372 ,n967);
    nor g1971(n1301 ,n426 ,n991);
    nor g1972(n1300 ,n442 ,n967);
    nor g1973(n1299 ,n443 ,n991);
    nor g1974(n1298 ,n3069 ,n1013);
    nor g1975(n1297 ,n3050 ,n992);
    nor g1976(n1296 ,n3066 ,n1013);
    nor g1977(n1295 ,n3067 ,n1013);
    nor g1978(n1294 ,n3065 ,n1013);
    nor g1979(n1293 ,n2[60] ,n1008);
    nor g1980(n1292 ,n3034 ,n1005);
    nor g1981(n1291 ,n3064 ,n1013);
    nor g1982(n1290 ,n3063 ,n998);
    nor g1983(n1289 ,n2[58] ,n1008);
    nor g1984(n1288 ,n3062 ,n998);
    nor g1985(n1287 ,n3061 ,n998);
    nor g1986(n1286 ,n3059 ,n998);
    nor g1987(n1285 ,n3075 ,n1012);
    nor g1988(n1284 ,n3058 ,n998);
    nor g1989(n1283 ,n3057 ,n998);
    nor g1990(n1282 ,n3085 ,n1004);
    nor g1991(n1281 ,n3025 ,n997);
    nor g1992(n1280 ,n3055 ,n992);
    nor g1993(n1279 ,n3027 ,n997);
    nor g1994(n1278 ,n3028 ,n997);
    nor g1995(n1277 ,n3036 ,n1005);
    nor g1996(n1276 ,n3047 ,n1000);
    nor g1997(n1275 ,n3068 ,n1013);
    nor g1998(n1274 ,n3030 ,n997);
    nor g1999(n1273 ,n3084 ,n1004);
    nor g2000(n1272 ,n3054 ,n992);
    nor g2001(n1271 ,n3031 ,n997);
    nor g2002(n1270 ,n2[28] ,n1001);
    nor g2003(n1269 ,n3033 ,n1005);
    nor g2004(n1268 ,n3060 ,n998);
    nor g2005(n1267 ,n3083 ,n1004);
    nor g2006(n1266 ,n2[13] ,n993);
    nor g2007(n1265 ,n3070 ,n1013);
    nor g2008(n1264 ,n3037 ,n1005);
    nor g2009(n1263 ,n3038 ,n1005);
    nor g2010(n1262 ,n2[16] ,n1010);
    nor g2011(n1261 ,n3039 ,n1005);
    nor g2012(n1260 ,n2[18] ,n1010);
    nor g2013(n1259 ,n3040 ,n1000);
    nor g2014(n1258 ,n2[19] ,n1010);
    nor g2015(n1257 ,n3035 ,n1005);
    nor g2016(n1256 ,n3052 ,n992);
    nor g2017(n1255 ,n2[21] ,n1010);
    nor g2018(n1254 ,n3041 ,n1000);
    nor g2019(n1253 ,n2[22] ,n1010);
    nor g2020(n1252 ,n2[50] ,n1006);
    nor g2021(n1251 ,n3026 ,n997);
    nor g2022(n1250 ,n3042 ,n1000);
    nor g2023(n1249 ,n3043 ,n1000);
    nor g2024(n1248 ,n3044 ,n1000);
    nor g2025(n1247 ,n2[27] ,n1001);
    nor g2026(n1246 ,n3045 ,n1000);
    nor g2027(n1245 ,n3087 ,n1004);
    nor g2028(n1244 ,n3046 ,n1000);
    nor g2029(n1243 ,n2[30] ,n1001);
    nor g2030(n1242 ,n3076 ,n1012);
    nor g2031(n1241 ,n3082 ,n1004);
    nor g2032(n1240 ,n3032 ,n1005);
    nor g2033(n1239 ,n3048 ,n992);
    nor g2034(n1238 ,n3049 ,n992);
    nor g2035(n1237 ,n3029 ,n997);
    nor g2036(n1236 ,n3086 ,n1004);
    nor g2037(n1235 ,n2[49] ,n1006);
    nor g2038(n1234 ,n3051 ,n992);
    nor g2039(n1233 ,n3053 ,n992);
    nor g2040(n1232 ,n3056 ,n998);
    or g2041(n1445 ,n298 ,n952);
    or g2042(n1444 ,n300 ,n952);
    or g2043(n1443 ,n301 ,n952);
    or g2044(n1442 ,n297 ,n952);
    or g2045(n1441 ,n302 ,n952);
    or g2046(n1440 ,n300 ,n983);
    or g2047(n1439 ,n534 ,n952);
    or g2048(n1438 ,n534 ,n983);
    or g2049(n1437 ,n301 ,n983);
    or g2050(n1436 ,n302 ,n983);
    or g2051(n1435 ,n299 ,n983);
    or g2052(n1434 ,n303 ,n983);
    or g2053(n1433 ,n298 ,n983);
    or g2054(n1432 ,n297 ,n983);
    or g2055(n1431 ,n303 ,n952);
    or g2056(n1430 ,n299 ,n952);
    nor g2057(n1207 ,n3[59] ,n984);
    nor g2058(n1206 ,n3077 ,n1012);
    nor g2059(n1205 ,n3078 ,n1012);
    nor g2060(n1204 ,n2[0] ,n995);
    nor g2061(n1203 ,n3079 ,n1012);
    nor g2062(n1202 ,n2[63] ,n1008);
    nor g2063(n1201 ,n3024 ,n997);
    nor g2064(n1200 ,n3080 ,n1004);
    nor g2065(n1199 ,n3081 ,n1004);
    nor g2066(n1198 ,n4[33] ,n988);
    nor g2067(n1197 ,n4[20] ,n989);
    nor g2068(n1196 ,n4[28] ,n981);
    nor g2069(n1195 ,n4[30] ,n981);
    nor g2070(n1194 ,n4[36] ,n988);
    nor g2071(n1193 ,n3[43] ,n982);
    nor g2072(n1192 ,n4[35] ,n988);
    nor g2073(n1191 ,n4[14] ,n985);
    nor g2074(n1190 ,n3[0] ,n986);
    nor g2075(n1189 ,n4[26] ,n981);
    nor g2076(n1188 ,n3[30] ,n981);
    nor g2077(n1187 ,n3[60] ,n984);
    nor g2078(n1186 ,n3[2] ,n986);
    nor g2079(n1185 ,n4[41] ,n982);
    nor g2080(n1184 ,n4[42] ,n982);
    nor g2081(n1183 ,n4[5] ,n986);
    nor g2082(n1182 ,n4[43] ,n982);
    nor g2083(n1181 ,n4[45] ,n982);
    nor g2084(n1180 ,n4[38] ,n988);
    nor g2085(n1179 ,n3[3] ,n986);
    nor g2086(n1178 ,n4[47] ,n982);
    nor g2087(n1177 ,n4[4] ,n986);
    nor g2088(n1176 ,n4[51] ,n987);
    nor g2089(n1175 ,n3[12] ,n985);
    nor g2090(n1174 ,n3[7] ,n986);
    nor g2091(n1173 ,n2[7] ,n996);
    nor g2092(n1172 ,n4[57] ,n984);
    nor g2093(n1171 ,n4[58] ,n984);
    nor g2094(n1170 ,n4[59] ,n984);
    nor g2095(n1169 ,n4[24] ,n981);
    nor g2096(n1168 ,n4[60] ,n984);
    nor g2097(n1167 ,n4[61] ,n984);
    nor g2098(n1166 ,n3[11] ,n985);
    nor g2099(n1165 ,n4[62] ,n984);
    nor g2100(n1164 ,n4[32] ,n988);
    nor g2101(n1163 ,n3[26] ,n981);
    nor g2102(n1162 ,n2[62] ,n1009);
    nor g2103(n1161 ,n3[13] ,n985);
    nor g2104(n1160 ,n3[14] ,n985);
    nor g2105(n1159 ,n3[15] ,n985);
    nor g2106(n1158 ,n4[63] ,n984);
    nor g2107(n1157 ,n3[16] ,n989);
    nor g2108(n1156 ,n3[17] ,n989);
    nor g2109(n1155 ,n4[19] ,n989);
    nor g2110(n1154 ,n4[52] ,n987);
    nor g2111(n1153 ,n3[18] ,n989);
    nor g2112(n1152 ,n4[50] ,n987);
    nor g2113(n1151 ,n3[19] ,n989);
    nor g2114(n1150 ,n4[44] ,n982);
    nor g2115(n1149 ,n4[18] ,n989);
    nor g2116(n1148 ,n3[20] ,n989);
    nor g2117(n1147 ,n3[21] ,n989);
    nor g2118(n1146 ,n4[31] ,n981);
    nor g2119(n1145 ,n3[22] ,n989);
    nor g2120(n1144 ,n3[23] ,n989);
    nor g2121(n1143 ,n3[24] ,n981);
    nor g2122(n1142 ,n4[49] ,n987);
    nor g2123(n1141 ,n3[25] ,n981);
    nor g2124(n1140 ,n3[27] ,n981);
    nor g2125(n1139 ,n3[28] ,n981);
    nor g2126(n1138 ,n3[29] ,n981);
    nor g2127(n1137 ,n3[31] ,n981);
    nor g2128(n1136 ,n3[6] ,n986);
    nor g2129(n1135 ,n3[32] ,n988);
    nor g2130(n1134 ,n3[33] ,n988);
    nor g2131(n1133 ,n4[39] ,n988);
    nor g2132(n1132 ,n3[35] ,n988);
    nor g2133(n1131 ,n3[1] ,n986);
    nor g2134(n1130 ,n3[36] ,n988);
    nor g2135(n1129 ,n3[4] ,n986);
    nor g2136(n1128 ,n3[37] ,n988);
    nor g2137(n1127 ,n3[38] ,n988);
    nor g2138(n1126 ,n4[40] ,n982);
    nor g2139(n1125 ,n3[39] ,n988);
    nor g2140(n1124 ,n4[48] ,n987);
    nor g2141(n1123 ,n3[40] ,n982);
    nor g2142(n1122 ,n4[29] ,n981);
    nor g2143(n1121 ,n3[41] ,n982);
    nor g2144(n1120 ,n3[42] ,n982);
    nor g2145(n1119 ,n3[44] ,n982);
    nor g2146(n1118 ,n3[45] ,n982);
    nor g2147(n1117 ,n2[44] ,n999);
    nor g2148(n1116 ,n3[46] ,n982);
    nor g2149(n1115 ,n4[0] ,n986);
    nor g2150(n1114 ,n3[47] ,n982);
    nor g2151(n1113 ,n3[48] ,n987);
    nor g2152(n1112 ,n3[49] ,n987);
    nor g2153(n1111 ,n3[50] ,n987);
    nor g2154(n1110 ,n3[51] ,n987);
    nor g2155(n1109 ,n3[52] ,n987);
    nor g2156(n1108 ,n3[53] ,n987);
    nor g2157(n1107 ,n3[54] ,n987);
    nor g2158(n1106 ,n3[5] ,n986);
    nor g2159(n1105 ,n2[11] ,n994);
    nor g2160(n1104 ,n3[55] ,n987);
    nor g2161(n1103 ,n3[56] ,n984);
    nor g2162(n1102 ,n3[9] ,n985);
    nor g2163(n1101 ,n3[57] ,n984);
    nor g2164(n1100 ,n3[58] ,n984);
    nor g2165(n1099 ,n2[4] ,n996);
    nor g2166(n1098 ,n3073 ,n1012);
    nor g2167(n1097 ,n4[46] ,n982);
    nor g2168(n1096 ,n3[61] ,n984);
    nor g2169(n1095 ,n4[10] ,n985);
    nor g2170(n1094 ,n4[7] ,n986);
    nor g2171(n1093 ,n3[62] ,n984);
    nor g2172(n1092 ,n2[61] ,n1009);
    nor g2173(n1091 ,n4[3] ,n986);
    nor g2174(n1090 ,n4[37] ,n988);
    nor g2175(n1089 ,n2[57] ,n1009);
    nor g2176(n1088 ,n4[1] ,n986);
    nor g2177(n1087 ,n4[2] ,n986);
    nor g2178(n1086 ,n4[22] ,n989);
    nor g2179(n1085 ,n4[55] ,n987);
    nor g2180(n1084 ,n4[56] ,n984);
    nor g2181(n1083 ,n4[6] ,n986);
    nor g2182(n1082 ,n4[8] ,n985);
    nor g2183(n1081 ,n2[56] ,n1009);
    nor g2184(n1080 ,n4[9] ,n985);
    nor g2185(n1079 ,n3[10] ,n985);
    nor g2186(n1078 ,n4[53] ,n987);
    nor g2187(n1077 ,n3[34] ,n988);
    nor g2188(n1076 ,n4[54] ,n987);
    nor g2189(n1075 ,n4[11] ,n985);
    nor g2190(n1074 ,n3[63] ,n984);
    nor g2191(n1073 ,n4[12] ,n985);
    nor g2192(n1072 ,n4[13] ,n985);
    nor g2193(n1071 ,n4[15] ,n985);
    nor g2194(n1070 ,n4[16] ,n989);
    nor g2195(n1069 ,n4[17] ,n989);
    nor g2196(n1068 ,n4[34] ,n988);
    nor g2197(n1067 ,n4[27] ,n981);
    nor g2198(n1066 ,n3[8] ,n985);
    nor g2199(n1065 ,n4[23] ,n989);
    nor g2200(n1064 ,n4[25] ,n981);
    nor g2201(n1063 ,n4[21] ,n989);
    nor g2202(n1062 ,n2[55] ,n1007);
    nor g2203(n1061 ,n2[3] ,n996);
    nor g2204(n1060 ,n2[10] ,n994);
    nor g2205(n1059 ,n7[15] ,n952);
    nor g2206(n1058 ,n7[63] ,n952);
    nor g2207(n1057 ,n2[54] ,n1007);
    nor g2208(n1056 ,n2[29] ,n1002);
    nor g2209(n1055 ,n2[41] ,n999);
    nor g2210(n1054 ,n7[55] ,n952);
    nor g2211(n1053 ,n2[59] ,n1009);
    nor g2212(n1052 ,n2[12] ,n994);
    nor g2213(n1051 ,n7[7] ,n952);
    nor g2214(n1050 ,n2[47] ,n999);
    nor g2215(n1049 ,n7[47] ,n952);
    nor g2216(n1048 ,n2[26] ,n1002);
    nor g2217(n1047 ,n2[2] ,n996);
    nor g2218(n1046 ,n2[51] ,n1007);
    nor g2219(n1045 ,n2[53] ,n1007);
    nor g2220(n1044 ,n2[52] ,n1007);
    nor g2221(n1043 ,n2[9] ,n994);
    nor g2222(n1042 ,n2[14] ,n994);
    nor g2223(n1041 ,n2[15] ,n994);
    nor g2224(n1040 ,n2[5] ,n996);
    nor g2225(n1039 ,n2[17] ,n1011);
    nor g2226(n1038 ,n7[23] ,n952);
    nor g2227(n1037 ,n2[6] ,n996);
    nor g2228(n1036 ,n2[8] ,n994);
    nor g2229(n1035 ,n2[23] ,n1011);
    nor g2230(n1034 ,n7[39] ,n952);
    nor g2231(n1033 ,n2[24] ,n1002);
    nor g2232(n1032 ,n2[25] ,n1002);
    nor g2233(n1031 ,n2[1] ,n996);
    nor g2234(n1030 ,n2[31] ,n1002);
    nor g2235(n1029 ,n2[46] ,n999);
    nor g2236(n1028 ,n2[32] ,n1003);
    nor g2237(n1027 ,n2[20] ,n1011);
    nor g2238(n1026 ,n7[31] ,n952);
    nor g2239(n1025 ,n2[33] ,n1003);
    nor g2240(n1024 ,n2[34] ,n1003);
    nor g2241(n1023 ,n2[35] ,n1003);
    nor g2242(n1022 ,n2[36] ,n1003);
    nor g2243(n1021 ,n2[37] ,n1003);
    nor g2244(n1020 ,n2[38] ,n1003);
    nor g2245(n1019 ,n2[39] ,n1003);
    nor g2246(n1018 ,n2[40] ,n999);
    nor g2247(n1017 ,n2[48] ,n1007);
    nor g2248(n1016 ,n2[42] ,n999);
    nor g2249(n1015 ,n2[43] ,n999);
    nor g2250(n1014 ,n2[45] ,n999);
    nor g2251(n1231 ,n976 ,n880);
    nor g2252(n1230 ,n976 ,n879);
    nor g2253(n1229 ,n978 ,n879);
    nor g2254(n1228 ,n973 ,n879);
    nor g2255(n1227 ,n974 ,n879);
    nor g2256(n1226 ,n979 ,n879);
    nor g2257(n1225 ,n979 ,n880);
    nor g2258(n1224 ,n975 ,n880);
    nor g2259(n1223 ,n978 ,n880);
    nor g2260(n1222 ,n973 ,n880);
    or g2261(n1221 ,n7[15] ,n983);
    or g2262(n1220 ,n7[7] ,n983);
    or g2263(n1219 ,n7[23] ,n983);
    nor g2264(n1218 ,n977 ,n880);
    or g2265(n1217 ,n7[39] ,n983);
    nor g2266(n1216 ,n980 ,n879);
    nor g2267(n1215 ,n974 ,n880);
    or g2268(n1214 ,n7[55] ,n983);
    nor g2269(n1213 ,n977 ,n879);
    nor g2270(n1212 ,n980 ,n880);
    or g2271(n1211 ,n7[63] ,n983);
    or g2272(n1210 ,n7[47] ,n983);
    nor g2273(n1209 ,n975 ,n879);
    or g2274(n1208 ,n7[31] ,n983);
    not g2275(n1010 ,n1011);
    not g2276(n1008 ,n1009);
    not g2277(n1006 ,n1007);
    not g2278(n1001 ,n1002);
    not g2279(n995 ,n996);
    not g2280(n993 ,n994);
    not g2281(n990 ,n991);
    or g2282(n1013 ,n299 ,n876);
    or g2283(n1012 ,n303 ,n876);
    nor g2284(n1011 ,n301 ,n875);
    nor g2285(n1009 ,n302 ,n875);
    nor g2286(n1007 ,n303 ,n875);
    or g2287(n1005 ,n297 ,n876);
    or g2288(n1004 ,n302 ,n876);
    nor g2289(n1003 ,n298 ,n875);
    nor g2290(n1002 ,n300 ,n875);
    or g2291(n1000 ,n301 ,n876);
    nor g2292(n999 ,n299 ,n875);
    or g2293(n998 ,n298 ,n876);
    or g2294(n997 ,n534 ,n876);
    nor g2295(n996 ,n534 ,n875);
    nor g2296(n994 ,n297 ,n875);
    or g2297(n992 ,n300 ,n876);
    nor g2298(n991 ,n7[15] ,n875);
    or g2299(n989 ,n301 ,n874);
    or g2300(n988 ,n298 ,n874);
    or g2301(n987 ,n303 ,n874);
    or g2302(n986 ,n534 ,n874);
    or g2303(n985 ,n297 ,n874);
    or g2304(n984 ,n302 ,n874);
    or g2305(n983 ,n796 ,n877);
    or g2306(n982 ,n299 ,n874);
    or g2307(n981 ,n300 ,n874);
    not g2308(n969 ,n970);
    not g2309(n966 ,n967);
    not g2310(n963 ,n964);
    not g2311(n960 ,n961);
    not g2312(n954 ,n955);
    nor g2313(n951 ,n1 ,n810);
    nor g2314(n950 ,n1 ,n812);
    nor g2315(n949 ,n1 ,n811);
    nor g2316(n980 ,n7[15] ,n874);
    nor g2317(n979 ,n7[47] ,n874);
    nor g2318(n978 ,n7[55] ,n874);
    nor g2319(n977 ,n7[7] ,n874);
    nor g2320(n976 ,n7[39] ,n874);
    nor g2321(n975 ,n7[63] ,n874);
    nor g2322(n974 ,n7[23] ,n874);
    nor g2323(n973 ,n7[31] ,n874);
    or g2324(n972 ,n7[55] ,n876);
    or g2325(n971 ,n7[39] ,n876);
    nor g2326(n970 ,n7[7] ,n875);
    or g2327(n968 ,n7[63] ,n876);
    nor g2328(n967 ,n7[63] ,n875);
    or g2329(n965 ,n7[7] ,n876);
    nor g2330(n964 ,n7[23] ,n875);
    or g2331(n962 ,n7[23] ,n876);
    nor g2332(n961 ,n7[31] ,n875);
    or g2333(n959 ,n7[15] ,n876);
    or g2334(n958 ,n7[31] ,n876);
    nor g2335(n957 ,n7[39] ,n875);
    nor g2336(n956 ,n7[47] ,n875);
    nor g2337(n955 ,n7[55] ,n875);
    or g2338(n953 ,n7[47] ,n876);
    nor g2339(n952 ,n873 ,n295);
    nor g2340(n948 ,n339 ,n293);
    nor g2341(n947 ,n522 ,n293);
    nor g2342(n946 ,n768 ,n296);
    nor g2343(n945 ,n503 ,n296);
    nor g2344(n944 ,n498 ,n293);
    nor g2345(n943 ,n527 ,n294);
    nor g2346(n942 ,n317 ,n296);
    nor g2347(n941 ,n501 ,n293);
    nor g2348(n940 ,n758 ,n293);
    nor g2349(n939 ,n338 ,n293);
    nor g2350(n938 ,n509 ,n296);
    nor g2351(n937 ,n538 ,n293);
    nor g2352(n936 ,n308 ,n294);
    nor g2353(n935 ,n505 ,n293);
    nor g2354(n934 ,n485 ,n293);
    nor g2355(n933 ,n484 ,n296);
    nor g2356(n932 ,n529 ,n296);
    nor g2357(n931 ,n524 ,n296);
    nor g2358(n930 ,n514 ,n293);
    nor g2359(n929 ,n349 ,n296);
    nor g2360(n928 ,n324 ,n296);
    nor g2361(n927 ,n481 ,n296);
    nor g2362(n926 ,n333 ,n293);
    nor g2363(n925 ,n335 ,n296);
    nor g2364(n924 ,n518 ,n296);
    nor g2365(n923 ,n500 ,n296);
    nor g2366(n922 ,n763 ,n296);
    nor g2367(n921 ,n496 ,n293);
    nor g2368(n920 ,n486 ,n294);
    nor g2369(n919 ,n328 ,n293);
    nor g2370(n918 ,n525 ,n293);
    nor g2371(n917 ,n530 ,n294);
    nor g2372(n916 ,n332 ,n294);
    nor g2373(n915 ,n516 ,n294);
    nor g2374(n914 ,n347 ,n294);
    nor g2375(n913 ,n764 ,n294);
    nor g2376(n912 ,n311 ,n294);
    nor g2377(n911 ,n309 ,n293);
    nor g2378(n910 ,n491 ,n293);
    nor g2379(n909 ,n352 ,n293);
    nor g2380(n908 ,n323 ,n293);
    nor g2381(n907 ,n321 ,n294);
    nor g2382(n906 ,n342 ,n294);
    nor g2383(n905 ,n316 ,n294);
    nor g2384(n904 ,n704 ,n294);
    nor g2385(n903 ,n354 ,n293);
    nor g2386(n902 ,n766 ,n293);
    nor g2387(n901 ,n531 ,n294);
    nor g2388(n900 ,n357 ,n294);
    nor g2389(n899 ,n305 ,n293);
    nor g2390(n898 ,n521 ,n293);
    nor g2391(n897 ,n511 ,n293);
    nor g2392(n896 ,n519 ,n296);
    nor g2393(n895 ,n306 ,n296);
    nor g2394(n894 ,n547 ,n293);
    nor g2395(n893 ,n537 ,n296);
    nor g2396(n892 ,n543 ,n296);
    nor g2397(n891 ,n523 ,n296);
    nor g2398(n890 ,n492 ,n293);
    nor g2399(n889 ,n353 ,n294);
    nor g2400(n888 ,n348 ,n293);
    nor g2401(n887 ,n515 ,n293);
    nor g2402(n886 ,n493 ,n293);
    nor g2403(n885 ,n340 ,n294);
    nor g2404(n884 ,n507 ,n296);
    nor g2405(n883 ,n319 ,n293);
    nor g2406(n882 ,n334 ,n293);
    nor g2407(n881 ,n312 ,n296);
    not g2408(n877 ,n878);
    not g2409(n874 ,n873);
    nor g2410(n872 ,n314 ,n294);
    nor g2411(n871 ,n542 ,n293);
    nor g2412(n870 ,n479 ,n296);
    nor g2413(n869 ,n761 ,n296);
    nor g2414(n868 ,n497 ,n296);
    nor g2415(n867 ,n554 ,n293);
    nor g2416(n866 ,n337 ,n296);
    nor g2417(n865 ,n359 ,n296);
    nor g2418(n864 ,n487 ,n296);
    nor g2419(n863 ,n344 ,n296);
    nor g2420(n862 ,n307 ,n296);
    nor g2421(n861 ,n310 ,n293);
    nor g2422(n860 ,n318 ,n296);
    nor g2423(n859 ,n345 ,n296);
    nor g2424(n858 ,n478 ,n294);
    nor g2425(n857 ,n343 ,n293);
    nor g2426(n856 ,n502 ,n293);
    nor g2427(n855 ,n326 ,n294);
    nor g2428(n854 ,n336 ,n294);
    nor g2429(n853 ,n494 ,n293);
    nor g2430(n852 ,n304 ,n294);
    nor g2431(n851 ,n356 ,n294);
    nor g2432(n850 ,n313 ,n296);
    nor g2433(n849 ,n341 ,n296);
    nor g2434(n848 ,n528 ,n293);
    nor g2435(n847 ,n564 ,n293);
    nor g2436(n846 ,n757 ,n296);
    nor g2437(n845 ,n355 ,n296);
    nor g2438(n844 ,n346 ,n296);
    nor g2439(n843 ,n329 ,n296);
    nor g2440(n842 ,n508 ,n294);
    nor g2441(n841 ,n499 ,n296);
    nor g2442(n840 ,n315 ,n294);
    nor g2443(n839 ,n350 ,n296);
    nor g2444(n838 ,n330 ,n293);
    nor g2445(n837 ,n322 ,n293);
    nor g2446(n836 ,n517 ,n296);
    nor g2447(n835 ,n331 ,n294);
    nor g2448(n834 ,n762 ,n296);
    nor g2449(n833 ,n520 ,n293);
    nor g2450(n832 ,n320 ,n294);
    nor g2451(n831 ,n488 ,n296);
    nor g2452(n830 ,n767 ,n296);
    nor g2453(n829 ,n760 ,n293);
    nor g2454(n828 ,n475 ,n293);
    nor g2455(n827 ,n490 ,n293);
    nor g2456(n826 ,n489 ,n294);
    nor g2457(n825 ,n325 ,n293);
    nor g2458(n824 ,n532 ,n293);
    nor g2459(n823 ,n477 ,n296);
    nor g2460(n822 ,n327 ,n294);
    nor g2461(n821 ,n759 ,n296);
    nor g2462(n820 ,n351 ,n294);
    nor g2463(n819 ,n358 ,n293);
    nor g2464(n818 ,n506 ,n293);
    nor g2465(n817 ,n533 ,n294);
    nor g2466(n816 ,n765 ,n294);
    nor g2467(n815 ,n510 ,n296);
    nor g2468(n814 ,n480 ,n296);
    nor g2469(n813 ,n476 ,n296);
    nor g2470(n812 ,n806 ,n802);
    nor g2471(n811 ,n808 ,n805);
    nor g2472(n810 ,n807 ,n803);
    nor g2473(n880 ,n795 ,n804);
    nor g2474(n879 ,n1 ,n801);
    nor g2475(n878 ,n797 ,n804);
    or g2476(n876 ,n6[0] ,n809);
    or g2477(n875 ,n792 ,n804);
    nor g2478(n873 ,n535 ,n809);
    nor g2479(n808 ,n535 ,n793);
    nor g2480(n807 ,n291 ,n793);
    nor g2481(n806 ,n292 ,n793);
    nor g2482(n805 ,n772 ,n794);
    or g2483(n809 ,n1 ,n798);
    not g2484(n293 ,n295);
    not g2485(n294 ,n295);
    not g2486(n295 ,n296);
    nor g2487(n803 ,n770 ,n794);
    nor g2488(n802 ,n785 ,n794);
    nor g2489(n801 ,n786 ,n794);
    or g2490(n804 ,n1 ,n799);
    or g2491(n296 ,n1 ,n800);
    not g2492(n800 ,n799);
    not g2493(n798 ,n797);
    nor g2494(n799 ,n291 ,n792);
    nor g2495(n797 ,n292 ,n790);
    not g2496(n796 ,n795);
    not g2497(n793 ,n794);
    nor g2498(n795 ,n535 ,n790);
    nor g2499(n794 ,n789 ,n791);
    not g2500(n792 ,n791);
    nor g2501(n791 ,n769 ,n788);
    not g2502(n790 ,n789);
    nor g2503(n789 ,n2543 ,n788);
    or g2504(n788 ,n781 ,n787);
    or g2505(n787 ,n780 ,n784);
    not g2506(n786 ,n785);
    or g2507(n784 ,n782 ,n777);
    xnor g2508(n785 ,n292 ,n535);
    nor g2509(n783 ,n482 ,n1);
    or g2510(n782 ,n561 ,n741);
    or g2511(n781 ,n744 ,n748);
    or g2512(n780 ,n742 ,n745);
    nor g2513(n779 ,n526 ,n1);
    nor g2514(n778 ,n512 ,n1);
    or g2515(n777 ,n738 ,n753);
    nor g2516(n776 ,n513 ,n1);
    nor g2517(n775 ,n495 ,n1);
    nor g2518(n774 ,n504 ,n1);
    nor g2519(n773 ,n483 ,n1);
    or g2520(n772 ,n6[0] ,n2543);
    nor g2521(n771 ,n8[0] ,n1);
    or g2522(n770 ,n535 ,n292);
    or g2523(n769 ,n6[0] ,n2542);
    not g2524(n768 ,n2992);
    not g2525(n767 ,n2982);
    not g2526(n766 ,n3010);
    not g2527(n765 ,n2969);
    not g2528(n764 ,n3011);
    not g2529(n763 ,n2980);
    not g2530(n762 ,n3021);
    not g2531(n761 ,n3013);
    not g2532(n760 ,n2962);
    not g2533(n759 ,n2997);
    not g2534(n758 ,n2966);
    not g2535(n757 ,n2971);
    not g2536(n756 ,n2[22]);
    not g2537(n755 ,n2[26]);
    not g2538(n754 ,n2[15]);
    not g2539(n753 ,n8[3]);
    not g2540(n752 ,n2[107]);
    not g2541(n751 ,n2[2]);
    not g2542(n750 ,n2[25]);
    not g2543(n749 ,n2[111]);
    not g2544(n748 ,n8[7]);
    not g2545(n747 ,n2[118]);
    not g2546(n746 ,n2[3]);
    not g2547(n745 ,n8[5]);
    not g2548(n744 ,n8[6]);
    not g2549(n743 ,n2[76]);
    not g2550(n742 ,n8[4]);
    not g2551(n741 ,n8[1]);
    not g2552(n740 ,n2[9]);
    not g2553(n739 ,n2[72]);
    not g2554(n738 ,n8[2]);
    not g2555(n737 ,n2[65]);
    not g2556(n736 ,n3[44]);
    not g2557(n735 ,n3[6]);
    not g2558(n734 ,n3[24]);
    not g2559(n733 ,n5[20]);
    not g2560(n732 ,n4[1]);
    not g2561(n731 ,n3[13]);
    not g2562(n730 ,n4[42]);
    not g2563(n729 ,n5[61]);
    not g2564(n728 ,n4[13]);
    not g2565(n727 ,n5[1]);
    not g2566(n726 ,n3[28]);
    not g2567(n725 ,n4[10]);
    not g2568(n724 ,n5[21]);
    not g2569(n723 ,n3[36]);
    not g2570(n722 ,n4[63]);
    not g2571(n721 ,n3[1]);
    not g2572(n720 ,n4[53]);
    not g2573(n719 ,n4[31]);
    not g2574(n718 ,n4[61]);
    not g2575(n717 ,n5[52]);
    not g2576(n716 ,n4[39]);
    not g2577(n715 ,n4[34]);
    not g2578(n714 ,n3[29]);
    not g2579(n713 ,n5[14]);
    not g2580(n712 ,n5[23]);
    not g2581(n711 ,n4[37]);
    not g2582(n710 ,n4[4]);
    not g2583(n709 ,n5[4]);
    not g2584(n708 ,n4[18]);
    not g2585(n707 ,n3[27]);
    not g2586(n706 ,n4[49]);
    not g2587(n705 ,n3[51]);
    not g2588(n704 ,n3040);
    not g2589(n703 ,n5[10]);
    not g2590(n702 ,n3[43]);
    not g2591(n701 ,n4[28]);
    not g2592(n700 ,n3[5]);
    not g2593(n699 ,n5[42]);
    not g2594(n698 ,n5[34]);
    not g2595(n697 ,n5[49]);
    not g2596(n696 ,n5[58]);
    not g2597(n695 ,n3[55]);
    not g2598(n694 ,n5[59]);
    not g2599(n693 ,n5[25]);
    not g2600(n692 ,n4[15]);
    not g2601(n691 ,n5[29]);
    not g2602(n690 ,n3[37]);
    not g2603(n689 ,n3[54]);
    not g2604(n688 ,n3[39]);
    not g2605(n687 ,n4[36]);
    not g2606(n686 ,n4[47]);
    not g2607(n685 ,n5[36]);
    not g2608(n684 ,n4[45]);
    not g2609(n683 ,n5[26]);
    not g2610(n682 ,n3[42]);
    not g2611(n681 ,n5[63]);
    not g2612(n680 ,n4[27]);
    not g2613(n679 ,n5[27]);
    not g2614(n678 ,n4[54]);
    not g2615(n677 ,n3[23]);
    not g2616(n676 ,n3[60]);
    not g2617(n675 ,n5[6]);
    not g2618(n674 ,n4[46]);
    not g2619(n673 ,n5[62]);
    not g2620(n672 ,n3[47]);
    not g2621(n671 ,n4[14]);
    not g2622(n670 ,n4[2]);
    not g2623(n669 ,n4[58]);
    not g2624(n668 ,n5[43]);
    not g2625(n667 ,n4[6]);
    not g2626(n666 ,n4[25]);
    not g2627(n665 ,n4[35]);
    not g2628(n664 ,n5[30]);
    not g2629(n663 ,n3[53]);
    not g2630(n662 ,n5[0]);
    not g2631(n661 ,n3[41]);
    not g2632(n660 ,n5[54]);
    not g2633(n659 ,n3[31]);
    not g2634(n658 ,n3[59]);
    not g2635(n657 ,n5[31]);
    not g2636(n656 ,n4[57]);
    not g2637(n655 ,n4[43]);
    not g2638(n654 ,n4[48]);
    not g2639(n653 ,n5[32]);
    not g2640(n652 ,n3[14]);
    not g2641(n651 ,n4[16]);
    not g2642(n650 ,n5[28]);
    not g2643(n649 ,n5[2]);
    not g2644(n648 ,n5[19]);
    not g2645(n647 ,n5[7]);
    not g2646(n646 ,n5[33]);
    not g2647(n645 ,n4[60]);
    not g2648(n644 ,n3[50]);
    not g2649(n643 ,n3[18]);
    not g2650(n642 ,n5[44]);
    not g2651(n641 ,n5[45]);
    not g2652(n640 ,n5[13]);
    not g2653(n639 ,n3[52]);
    not g2654(n638 ,n5[46]);
    not g2655(n637 ,n4[9]);
    not g2656(n636 ,n4[30]);
    not g2657(n635 ,n5[37]);
    not g2658(n634 ,n3[25]);
    not g2659(n633 ,n4[56]);
    not g2660(n632 ,n4[5]);
    not g2661(n631 ,n3[2]);
    not g2662(n630 ,n4[50]);
    not g2663(n629 ,n3[0]);
    not g2664(n628 ,n5[8]);
    not g2665(n627 ,n5[24]);
    not g2666(n626 ,n5[48]);
    not g2667(n625 ,n4[8]);
    not g2668(n624 ,n4[52]);
    not g2669(n623 ,n5[56]);
    not g2670(n622 ,n5[51]);
    not g2671(n621 ,n3[26]);
    not g2672(n620 ,n4[20]);
    not g2673(n619 ,n4[51]);
    not g2674(n618 ,n5[9]);
    not g2675(n617 ,n5[5]);
    not g2676(n616 ,n3[22]);
    not g2677(n615 ,n3[21]);
    not g2678(n614 ,n3[61]);
    not g2679(n613 ,n4[23]);
    not g2680(n612 ,n4[62]);
    not g2681(n611 ,n3[17]);
    not g2682(n610 ,n3[15]);
    not g2683(n609 ,n3[33]);
    not g2684(n608 ,n3[46]);
    not g2685(n607 ,n5[22]);
    not g2686(n606 ,n5[39]);
    not g2687(n605 ,n4[32]);
    not g2688(n604 ,n3[11]);
    not g2689(n603 ,n3[16]);
    not g2690(n602 ,n4[41]);
    not g2691(n601 ,n5[38]);
    not g2692(n600 ,n3[10]);
    not g2693(n599 ,n5[40]);
    not g2694(n598 ,n5[12]);
    not g2695(n597 ,n4[19]);
    not g2696(n596 ,n5[11]);
    not g2697(n595 ,n4[7]);
    not g2698(n594 ,n5[55]);
    not g2699(n593 ,n5[18]);
    not g2700(n592 ,n4[17]);
    not g2701(n591 ,n5[53]);
    not g2702(n590 ,n3[63]);
    not g2703(n589 ,n3[32]);
    not g2704(n588 ,n4[38]);
    not g2705(n587 ,n4[40]);
    not g2706(n586 ,n4[24]);
    not g2707(n585 ,n4[12]);
    not g2708(n584 ,n4[59]);
    not g2709(n583 ,n4[11]);
    not g2710(n582 ,n4[26]);
    not g2711(n581 ,n3[40]);
    not g2712(n580 ,n4[55]);
    not g2713(n579 ,n3[38]);
    not g2714(n578 ,n3[34]);
    not g2715(n577 ,n3[19]);
    not g2716(n576 ,n3[48]);
    not g2717(n575 ,n4[29]);
    not g2718(n574 ,n4[3]);
    not g2719(n573 ,n3[4]);
    not g2720(n572 ,n3[56]);
    not g2721(n571 ,n5[57]);
    not g2722(n570 ,n3[12]);
    not g2723(n569 ,n3[62]);
    not g2724(n568 ,n4[44]);
    not g2725(n567 ,n3[58]);
    not g2726(n566 ,n5[15]);
    not g2727(n565 ,n3[3]);
    not g2728(n564 ,n3080);
    not g2729(n563 ,n5[16]);
    not g2730(n562 ,n5[41]);
    not g2731(n561 ,n8[0]);
    not g2732(n560 ,n5[17]);
    not g2733(n559 ,n3[57]);
    not g2734(n558 ,n3[8]);
    not g2735(n557 ,n3[30]);
    not g2736(n556 ,n3[49]);
    not g2737(n555 ,n5[47]);
    not g2738(n554 ,n3062);
    not g2739(n553 ,n3[20]);
    not g2740(n552 ,n5[3]);
    not g2741(n551 ,n4[0]);
    not g2742(n550 ,n4[22]);
    not g2743(n549 ,n5[50]);
    not g2744(n548 ,n3[9]);
    not g2745(n547 ,n3047);
    not g2746(n546 ,n3[45]);
    not g2747(n545 ,n5[35]);
    not g2748(n544 ,n3[7]);
    not g2749(n543 ,n3048);
    not g2750(n542 ,n3084);
    not g2751(n541 ,n4[33]);
    not g2752(n540 ,n3[35]);
    not g2753(n539 ,n5[60]);
    not g2754(n538 ,n3085);
    not g2755(n537 ,n3071);
    not g2756(n536 ,n4[21]);
    not g2757(n292 ,n2542);
    buf g2758(n6[1] ,n2542);
    not g2759(n291 ,n2543);
    buf g2760(n6[2] ,n2543);
    not g2761(n535 ,n6[0]);
    not g2762(n534 ,n7[7]);
    not g2763(n533 ,n3016);
    not g2764(n532 ,n2965);
    not g2765(n531 ,n2973);
    not g2766(n530 ,n3001);
    not g2767(n529 ,n3019);
    not g2768(n528 ,n2977);
    not g2769(n527 ,n2994);
    not g2770(n526 ,n3220);
    not g2771(n525 ,n2976);
    not g2772(n524 ,n3004);
    not g2773(n523 ,n2991);
    not g2774(n522 ,n3023);
    not g2775(n521 ,n2968);
    not g2776(n520 ,n2960);
    not g2777(n519 ,n2983);
    not g2778(n518 ,n3003);
    not g2779(n517 ,n2970);
    not g2780(n516 ,n2995);
    not g2781(n515 ,n2990);
    not g2782(n514 ,n3002);
    not g2783(n513 ,n3216);
    not g2784(n512 ,n3219);
    not g2785(n511 ,n2972);
    not g2786(n510 ,n2975);
    not g2787(n509 ,n2986);
    not g2788(n508 ,n3006);
    not g2789(n507 ,n3018);
    not g2790(n506 ,n3007);
    not g2791(n505 ,n2974);
    not g2792(n504 ,n3221);
    not g2793(n503 ,n2993);
    not g2794(n502 ,n2967);
    not g2795(n501 ,n3012);
    not g2796(n500 ,n2999);
    not g2797(n499 ,n2984);
    not g2798(n498 ,n3022);
    not g2799(n497 ,n3020);
    not g2800(n496 ,n2978);
    not g2801(n495 ,n3222);
    not g2802(n494 ,n2998);
    not g2803(n493 ,n3009);
    not g2804(n492 ,n3000);
    not g2805(n491 ,n2979);
    not g2806(n490 ,n3015);
    not g2807(n489 ,n2963);
    not g2808(n488 ,n2987);
    not g2809(n487 ,n2989);
    not g2810(n486 ,n3014);
    not g2811(n485 ,n2964);
    not g2812(n484 ,n3017);
    not g2813(n483 ,n3217);
    not g2814(n482 ,n3218);
    not g2815(n481 ,n2985);
    not g2816(n480 ,n2981);
    not g2817(n479 ,n3005);
    not g2818(n478 ,n3008);
    not g2819(n477 ,n2961);
    not g2820(n476 ,n2988);
    not g2821(n475 ,n2996);
    not g2822(n474 ,n2[46]);
    not g2823(n473 ,n2[61]);
    not g2824(n472 ,n2[87]);
    not g2825(n471 ,n2[29]);
    not g2826(n470 ,n2[59]);
    not g2827(n469 ,n2[16]);
    not g2828(n468 ,n2[35]);
    not g2829(n467 ,n2[7]);
    not g2830(n466 ,n2[119]);
    not g2831(n465 ,n2[80]);
    not g2832(n464 ,n2[60]);
    not g2833(n463 ,n2[89]);
    not g2834(n462 ,n2[38]);
    not g2835(n461 ,n2[84]);
    not g2836(n460 ,n2[31]);
    not g2837(n459 ,n2[54]);
    not g2838(n458 ,n2[52]);
    not g2839(n457 ,n2[33]);
    not g2840(n456 ,n2[96]);
    not g2841(n455 ,n2[93]);
    not g2842(n454 ,n2[102]);
    not g2843(n453 ,n2[112]);
    not g2844(n452 ,n2[66]);
    not g2845(n451 ,n2[116]);
    not g2846(n450 ,n2[32]);
    not g2847(n449 ,n2[8]);
    not g2848(n448 ,n2[1]);
    not g2849(n447 ,n2[53]);
    not g2850(n446 ,n2[75]);
    not g2851(n445 ,n2[55]);
    not g2852(n444 ,n2[24]);
    not g2853(n443 ,n2[11]);
    not g2854(n442 ,n2[56]);
    not g2855(n441 ,n2[6]);
    not g2856(n440 ,n2[18]);
    not g2857(n439 ,n2[0]);
    not g2858(n438 ,n2[45]);
    not g2859(n437 ,n2[34]);
    not g2860(n436 ,n2[48]);
    not g2861(n435 ,n2[17]);
    not g2862(n434 ,n2[97]);
    not g2863(n433 ,n2[21]);
    not g2864(n432 ,n2[50]);
    not g2865(n431 ,n2[27]);
    not g2866(n430 ,n2[105]);
    not g2867(n429 ,n2[127]);
    not g2868(n428 ,n2[67]);
    not g2869(n427 ,n2[28]);
    not g2870(n426 ,n2[10]);
    not g2871(n425 ,n2[37]);
    not g2872(n424 ,n2[57]);
    not g2873(n423 ,n2[42]);
    not g2874(n422 ,n2[19]);
    not g2875(n421 ,n2[74]);
    not g2876(n420 ,n2[39]);
    not g2877(n419 ,n2[63]);
    not g2878(n418 ,n2[20]);
    not g2879(n417 ,n2[4]);
    not g2880(n416 ,n2[126]);
    not g2881(n415 ,n2[47]);
    not g2882(n414 ,n2[79]);
    not g2883(n413 ,n2[123]);
    not g2884(n412 ,n2[58]);
    not g2885(n411 ,n2[68]);
    not g2886(n410 ,n2[117]);
    not g2887(n409 ,n2[94]);
    not g2888(n408 ,n2[120]);
    not g2889(n407 ,n2[98]);
    not g2890(n406 ,n2[41]);
    not g2891(n405 ,n2[108]);
    not g2892(n404 ,n2[125]);
    not g2893(n403 ,n2[91]);
    not g2894(n402 ,n2[64]);
    not g2895(n401 ,n2[99]);
    not g2896(n400 ,n2[69]);
    not g2897(n399 ,n2[77]);
    not g2898(n398 ,n2[82]);
    not g2899(n397 ,n2[73]);
    not g2900(n396 ,n2[83]);
    not g2901(n395 ,n2[5]);
    not g2902(n394 ,n2[36]);
    not g2903(n393 ,n2[30]);
    not g2904(n392 ,n2[81]);
    not g2905(n391 ,n2[114]);
    not g2906(n390 ,n2[115]);
    not g2907(n389 ,n2[124]);
    not g2908(n388 ,n2[71]);
    not g2909(n387 ,n2[14]);
    not g2910(n386 ,n2[88]);
    not g2911(n385 ,n2[95]);
    not g2912(n384 ,n2[44]);
    not g2913(n383 ,n2[51]);
    not g2914(n382 ,n2[86]);
    not g2915(n381 ,n2[113]);
    not g2916(n380 ,n2[90]);
    not g2917(n379 ,n2[70]);
    not g2918(n378 ,n2[40]);
    not g2919(n377 ,n2[43]);
    not g2920(n376 ,n2[13]);
    not g2921(n375 ,n2[122]);
    not g2922(n374 ,n2[106]);
    not g2923(n373 ,n2[104]);
    not g2924(n372 ,n2[62]);
    not g2925(n371 ,n2[100]);
    not g2926(n370 ,n2[12]);
    not g2927(n369 ,n2[85]);
    not g2928(n368 ,n2[121]);
    not g2929(n367 ,n2[101]);
    not g2930(n366 ,n2[23]);
    not g2931(n365 ,n2[78]);
    not g2932(n364 ,n2[92]);
    not g2933(n363 ,n2[109]);
    not g2934(n362 ,n2[103]);
    not g2935(n361 ,n2[49]);
    not g2936(n360 ,n2[110]);
    not g2937(n359 ,n3063);
    not g2938(n358 ,n3051);
    not g2939(n357 ,n3043);
    not g2940(n356 ,n3061);
    not g2941(n355 ,n3081);
    not g2942(n354 ,n3041);
    not g2943(n353 ,n3050);
    not g2944(n352 ,n3037);
    not g2945(n351 ,n3057);
    not g2946(n350 ,n3026);
    not g2947(n349 ,n3028);
    not g2948(n348 ,n3024);
    not g2949(n347 ,n3074);
    not g2950(n346 ,n3032);
    not g2951(n345 ,n3066);
    not g2952(n344 ,n3042);
    not g2953(n343 ,n3067);
    not g2954(n342 ,n3049);
    not g2955(n341 ,n3078);
    not g2956(n340 ,n3052);
    not g2957(n339 ,n3083);
    not g2958(n338 ,n3054);
    not g2959(n337 ,n3064);
    not g2960(n336 ,n3069);
    not g2961(n335 ,n3077);
    not g2962(n334 ,n3045);
    not g2963(n333 ,n3027);
    not g2964(n332 ,n3031);
    not g2965(n331 ,n3087);
    not g2966(n330 ,n3086);
    not g2967(n329 ,n3082);
    not g2968(n328 ,n3076);
    not g2969(n327 ,n3058);
    not g2970(n326 ,n3068);
    not g2971(n325 ,n3059);
    not g2972(n324 ,n3029);
    not g2973(n323 ,n3075);
    not g2974(n322 ,n3060);
    not g2975(n321 ,n3038);
    not g2976(n320 ,n3072);
    not g2977(n319 ,n3053);
    not g2978(n318 ,n3034);
    not g2979(n317 ,n3055);
    not g2980(n316 ,n3039);
    not g2981(n315 ,n3033);
    not g2982(n314 ,n3056);
    not g2983(n313 ,n3036);
    not g2984(n312 ,n3073);
    not g2985(n311 ,n3035);
    not g2986(n310 ,n3065);
    not g2987(n309 ,n3079);
    not g2988(n308 ,n3025);
    not g2989(n307 ,n3030);
    not g2990(n306 ,n3046);
    not g2991(n305 ,n3044);
    not g2992(n304 ,n3070);
    not g2993(n303 ,n7[55]);
    not g2994(n302 ,n7[63]);
    not g2995(n301 ,n7[23]);
    not g2996(n300 ,n7[31]);
    not g2997(n299 ,n7[47]);
    not g2998(n298 ,n7[39]);
    not g2999(n297 ,n7[15]);
    xnor g3000(n3087 ,n78 ,n266);
    nor g3001(n266 ,n51 ,n265);
    xnor g3002(n3086 ,n94 ,n264);
    nor g3003(n265 ,n94 ,n264);
    nor g3004(n264 ,n40 ,n263);
    xnor g3005(n3085 ,n115 ,n262);
    nor g3006(n263 ,n115 ,n262);
    nor g3007(n262 ,n69 ,n261);
    xnor g3008(n3084 ,n97 ,n260);
    nor g3009(n261 ,n97 ,n260);
    nor g3010(n260 ,n43 ,n259);
    xnor g3011(n3083 ,n102 ,n258);
    nor g3012(n259 ,n102 ,n258);
    nor g3013(n258 ,n55 ,n257);
    xnor g3014(n3082 ,n124 ,n256);
    nor g3015(n257 ,n124 ,n256);
    nor g3016(n256 ,n36 ,n255);
    xnor g3017(n3081 ,n107 ,n254);
    nor g3018(n255 ,n107 ,n254);
    nor g3019(n254 ,n70 ,n253);
    xnor g3020(n3080 ,n96 ,n252);
    nor g3021(n253 ,n96 ,n252);
    nor g3022(n252 ,n16 ,n251);
    xnor g3023(n3079 ,n135 ,n250);
    nor g3024(n251 ,n135 ,n250);
    nor g3025(n250 ,n35 ,n249);
    xnor g3026(n3078 ,n89 ,n248);
    nor g3027(n249 ,n89 ,n248);
    nor g3028(n248 ,n62 ,n247);
    xnor g3029(n3077 ,n130 ,n246);
    nor g3030(n247 ,n130 ,n246);
    nor g3031(n246 ,n47 ,n245);
    xnor g3032(n3076 ,n125 ,n244);
    nor g3033(n245 ,n125 ,n244);
    nor g3034(n244 ,n39 ,n243);
    xnor g3035(n3075 ,n119 ,n242);
    nor g3036(n243 ,n119 ,n242);
    nor g3037(n242 ,n31 ,n241);
    xnor g3038(n3074 ,n111 ,n240);
    nor g3039(n241 ,n111 ,n240);
    nor g3040(n240 ,n27 ,n239);
    xnor g3041(n3073 ,n100 ,n238);
    nor g3042(n239 ,n100 ,n238);
    nor g3043(n238 ,n21 ,n237);
    xnor g3044(n3072 ,n109 ,n236);
    nor g3045(n237 ,n109 ,n236);
    nor g3046(n236 ,n14 ,n235);
    xnor g3047(n3071 ,n85 ,n234);
    nor g3048(n235 ,n85 ,n234);
    nor g3049(n234 ,n57 ,n233);
    xnor g3050(n3070 ,n80 ,n232);
    nor g3051(n233 ,n80 ,n232);
    nor g3052(n232 ,n75 ,n231);
    xnor g3053(n3069 ,n82 ,n230);
    nor g3054(n231 ,n82 ,n230);
    nor g3055(n230 ,n56 ,n229);
    xnor g3056(n3068 ,n88 ,n228);
    nor g3057(n229 ,n88 ,n228);
    nor g3058(n228 ,n63 ,n227);
    xnor g3059(n3067 ,n137 ,n226);
    nor g3060(n227 ,n137 ,n226);
    nor g3061(n226 ,n30 ,n225);
    xnor g3062(n3066 ,n133 ,n224);
    nor g3063(n225 ,n133 ,n224);
    nor g3064(n224 ,n49 ,n223);
    xnor g3065(n3065 ,n128 ,n222);
    nor g3066(n223 ,n128 ,n222);
    nor g3067(n222 ,n25 ,n221);
    xnor g3068(n3064 ,n98 ,n220);
    nor g3069(n221 ,n98 ,n220);
    nor g3070(n220 ,n41 ,n219);
    xnor g3071(n3063 ,n122 ,n218);
    nor g3072(n219 ,n122 ,n218);
    nor g3073(n218 ,n66 ,n217);
    xnor g3074(n3062 ,n118 ,n216);
    nor g3075(n217 ,n118 ,n216);
    nor g3076(n216 ,n33 ,n215);
    xnor g3077(n3061 ,n113 ,n214);
    nor g3078(n215 ,n113 ,n214);
    nor g3079(n214 ,n38 ,n213);
    xnor g3080(n3060 ,n110 ,n212);
    nor g3081(n213 ,n110 ,n212);
    nor g3082(n212 ,n53 ,n211);
    xnor g3083(n3059 ,n108 ,n210);
    nor g3084(n211 ,n108 ,n210);
    nor g3085(n210 ,n17 ,n209);
    xnor g3086(n3058 ,n104 ,n208);
    nor g3087(n209 ,n104 ,n208);
    nor g3088(n208 ,n23 ,n207);
    xnor g3089(n3057 ,n99 ,n206);
    nor g3090(n207 ,n99 ,n206);
    nor g3091(n206 ,n46 ,n205);
    xnor g3092(n3056 ,n92 ,n204);
    nor g3093(n205 ,n92 ,n204);
    nor g3094(n204 ,n72 ,n203);
    xnor g3095(n3055 ,n87 ,n202);
    nor g3096(n203 ,n87 ,n202);
    nor g3097(n202 ,n73 ,n201);
    xnor g3098(n3054 ,n84 ,n200);
    nor g3099(n201 ,n84 ,n200);
    nor g3100(n200 ,n15 ,n199);
    xnor g3101(n3053 ,n79 ,n198);
    nor g3102(n199 ,n79 ,n198);
    nor g3103(n198 ,n52 ,n197);
    xnor g3104(n3052 ,n81 ,n196);
    nor g3105(n197 ,n81 ,n196);
    nor g3106(n196 ,n67 ,n195);
    xnor g3107(n3051 ,n83 ,n194);
    nor g3108(n195 ,n83 ,n194);
    nor g3109(n194 ,n64 ,n193);
    xnor g3110(n3050 ,n86 ,n192);
    nor g3111(n193 ,n86 ,n192);
    nor g3112(n192 ,n44 ,n191);
    xnor g3113(n3049 ,n91 ,n190);
    nor g3114(n191 ,n91 ,n190);
    nor g3115(n190 ,n42 ,n189);
    xnor g3116(n3048 ,n90 ,n188);
    nor g3117(n189 ,n90 ,n188);
    nor g3118(n188 ,n18 ,n187);
    xnor g3119(n3047 ,n139 ,n186);
    nor g3120(n187 ,n139 ,n186);
    nor g3121(n186 ,n61 ,n185);
    xnor g3122(n3046 ,n136 ,n184);
    nor g3123(n185 ,n136 ,n184);
    nor g3124(n184 ,n58 ,n183);
    xnor g3125(n3045 ,n134 ,n182);
    nor g3126(n183 ,n134 ,n182);
    nor g3127(n182 ,n54 ,n181);
    xnor g3128(n3044 ,n132 ,n180);
    nor g3129(n181 ,n132 ,n180);
    nor g3130(n180 ,n50 ,n179);
    xnor g3131(n3043 ,n131 ,n178);
    nor g3132(n179 ,n131 ,n178);
    nor g3133(n178 ,n48 ,n177);
    xnor g3134(n3042 ,n129 ,n176);
    nor g3135(n177 ,n129 ,n176);
    nor g3136(n176 ,n29 ,n175);
    xnor g3137(n3041 ,n126 ,n174);
    nor g3138(n175 ,n126 ,n174);
    nor g3139(n174 ,n20 ,n173);
    xnor g3140(n3040 ,n105 ,n172);
    nor g3141(n173 ,n105 ,n172);
    nor g3142(n172 ,n22 ,n171);
    xnor g3143(n3039 ,n123 ,n170);
    nor g3144(n171 ,n123 ,n170);
    nor g3145(n170 ,n65 ,n169);
    xnor g3146(n3038 ,n121 ,n168);
    nor g3147(n169 ,n121 ,n168);
    nor g3148(n168 ,n37 ,n167);
    xnor g3149(n3037 ,n120 ,n166);
    nor g3150(n167 ,n120 ,n166);
    nor g3151(n166 ,n34 ,n165);
    xnor g3152(n3036 ,n117 ,n164);
    nor g3153(n165 ,n117 ,n164);
    nor g3154(n164 ,n68 ,n163);
    xnor g3155(n3035 ,n116 ,n162);
    nor g3156(n163 ,n116 ,n162);
    nor g3157(n162 ,n32 ,n161);
    xnor g3158(n3034 ,n114 ,n160);
    nor g3159(n161 ,n114 ,n160);
    nor g3160(n160 ,n45 ,n159);
    xnor g3161(n3033 ,n112 ,n158);
    nor g3162(n159 ,n112 ,n158);
    nor g3163(n158 ,n28 ,n157);
    xnor g3164(n3032 ,n127 ,n156);
    nor g3165(n157 ,n127 ,n156);
    nor g3166(n156 ,n59 ,n155);
    xnor g3167(n3031 ,n93 ,n154);
    nor g3168(n155 ,n93 ,n154);
    nor g3169(n154 ,n26 ,n153);
    xnor g3170(n3030 ,n138 ,n152);
    nor g3171(n153 ,n138 ,n152);
    nor g3172(n152 ,n24 ,n151);
    xnor g3173(n3029 ,n106 ,n150);
    nor g3174(n151 ,n106 ,n150);
    nor g3175(n150 ,n74 ,n149);
    xnor g3176(n3028 ,n103 ,n148);
    nor g3177(n149 ,n103 ,n148);
    nor g3178(n148 ,n71 ,n147);
    xor g3179(n3027 ,n101 ,n145);
    nor g3180(n147 ,n101 ,n146);
    not g3181(n146 ,n145);
    nor g3182(n145 ,n60 ,n144);
    xnor g3183(n3026 ,n140 ,n142);
    nor g3184(n144 ,n140 ,n143);
    not g3185(n143 ,n142);
    nor g3186(n142 ,n19 ,n141);
    xnor g3187(n3025 ,n95 ,n77);
    nor g3188(n141 ,n77 ,n95);
    nor g3189(n3024 ,n77 ,n76);
    xnor g3190(n140 ,n3154 ,n3090);
    xnor g3191(n139 ,n3175 ,n3111);
    xnor g3192(n138 ,n3158 ,n3094);
    xnor g3193(n137 ,n3195 ,n3131);
    xnor g3194(n136 ,n3174 ,n3110);
    xnor g3195(n135 ,n3207 ,n3143);
    xnor g3196(n134 ,n3173 ,n3109);
    xnor g3197(n133 ,n3194 ,n3130);
    xnor g3198(n132 ,n3172 ,n3108);
    xnor g3199(n131 ,n3171 ,n3107);
    xnor g3200(n130 ,n3205 ,n3141);
    xnor g3201(n129 ,n3170 ,n3106);
    xnor g3202(n128 ,n3193 ,n3129);
    xnor g3203(n127 ,n3160 ,n3096);
    xnor g3204(n126 ,n3169 ,n3105);
    xnor g3205(n125 ,n3204 ,n3140);
    xnor g3206(n124 ,n3210 ,n3146);
    xnor g3207(n123 ,n3167 ,n3103);
    xnor g3208(n122 ,n3191 ,n3127);
    xnor g3209(n121 ,n3166 ,n3102);
    xnor g3210(n120 ,n3165 ,n3101);
    xnor g3211(n119 ,n3203 ,n3139);
    xnor g3212(n118 ,n3190 ,n3126);
    xnor g3213(n117 ,n3164 ,n3100);
    xnor g3214(n116 ,n3163 ,n3099);
    xnor g3215(n115 ,n3213 ,n3149);
    xnor g3216(n114 ,n3162 ,n3098);
    xnor g3217(n113 ,n3189 ,n3125);
    xnor g3218(n112 ,n3161 ,n3097);
    xnor g3219(n111 ,n3202 ,n3138);
    xnor g3220(n110 ,n3188 ,n3124);
    xnor g3221(n109 ,n3200 ,n3136);
    xnor g3222(n108 ,n3187 ,n3123);
    xnor g3223(n107 ,n3209 ,n3145);
    xnor g3224(n106 ,n3157 ,n3093);
    xnor g3225(n105 ,n3168 ,n3104);
    xnor g3226(n104 ,n3186 ,n3122);
    xnor g3227(n103 ,n3156 ,n3092);
    xnor g3228(n102 ,n3211 ,n3147);
    xnor g3229(n101 ,n3155 ,n3091);
    xnor g3230(n100 ,n3201 ,n3137);
    xnor g3231(n99 ,n3185 ,n3121);
    xnor g3232(n98 ,n3192 ,n3128);
    xnor g3233(n97 ,n3212 ,n3148);
    xnor g3234(n96 ,n3208 ,n3144);
    xnor g3235(n95 ,n3153 ,n3089);
    xnor g3236(n94 ,n3214 ,n3150);
    xnor g3237(n93 ,n3159 ,n3095);
    xnor g3238(n92 ,n3184 ,n3120);
    xnor g3239(n91 ,n3177 ,n3113);
    xnor g3240(n90 ,n3176 ,n3112);
    xnor g3241(n89 ,n3206 ,n3142);
    xnor g3242(n88 ,n3196 ,n3132);
    xnor g3243(n87 ,n3183 ,n3119);
    xnor g3244(n86 ,n3178 ,n3114);
    xnor g3245(n85 ,n3199 ,n3135);
    xnor g3246(n84 ,n3182 ,n3118);
    xnor g3247(n83 ,n3179 ,n3115);
    xnor g3248(n82 ,n3197 ,n3133);
    xnor g3249(n81 ,n3180 ,n3116);
    xnor g3250(n80 ,n3198 ,n3134);
    xnor g3251(n79 ,n3181 ,n3117);
    xnor g3252(n78 ,n3215 ,n3151);
    nor g3253(n76 ,n3152 ,n3088);
    nor g3254(n75 ,n3197 ,n3133);
    nor g3255(n74 ,n3156 ,n3092);
    nor g3256(n73 ,n3182 ,n3118);
    nor g3257(n72 ,n3183 ,n3119);
    nor g3258(n71 ,n3155 ,n3091);
    nor g3259(n70 ,n3208 ,n3144);
    nor g3260(n69 ,n3212 ,n3148);
    nor g3261(n68 ,n3163 ,n3099);
    nor g3262(n67 ,n3179 ,n3115);
    nor g3263(n66 ,n3190 ,n3126);
    nor g3264(n65 ,n3166 ,n3102);
    nor g3265(n64 ,n3178 ,n3114);
    nor g3266(n63 ,n3195 ,n3131);
    nor g3267(n62 ,n3205 ,n3141);
    nor g3268(n61 ,n3174 ,n3110);
    nor g3269(n60 ,n12 ,n11);
    nor g3270(n59 ,n3159 ,n3095);
    nor g3271(n58 ,n3173 ,n3109);
    nor g3272(n57 ,n3198 ,n3134);
    nor g3273(n56 ,n3196 ,n3132);
    nor g3274(n55 ,n3210 ,n3146);
    nor g3275(n54 ,n3172 ,n3108);
    nor g3276(n53 ,n3187 ,n3123);
    nor g3277(n52 ,n3180 ,n3116);
    nor g3278(n51 ,n3214 ,n3150);
    nor g3279(n50 ,n3171 ,n3107);
    nor g3280(n49 ,n3193 ,n3129);
    nor g3281(n48 ,n3170 ,n3106);
    nor g3282(n47 ,n3204 ,n3140);
    nor g3283(n46 ,n3184 ,n3120);
    nor g3284(n77 ,n13 ,n10);
    nor g3285(n45 ,n3161 ,n3097);
    nor g3286(n44 ,n3177 ,n3113);
    nor g3287(n43 ,n3211 ,n3147);
    nor g3288(n42 ,n3176 ,n3112);
    nor g3289(n41 ,n3191 ,n3127);
    nor g3290(n40 ,n3213 ,n3149);
    nor g3291(n39 ,n3203 ,n3139);
    nor g3292(n38 ,n3188 ,n3124);
    nor g3293(n37 ,n3165 ,n3101);
    nor g3294(n36 ,n3209 ,n3145);
    nor g3295(n35 ,n3206 ,n3142);
    nor g3296(n34 ,n3164 ,n3100);
    nor g3297(n33 ,n3189 ,n3125);
    nor g3298(n32 ,n3162 ,n3098);
    nor g3299(n31 ,n3202 ,n3138);
    nor g3300(n30 ,n3194 ,n3130);
    nor g3301(n29 ,n3169 ,n3105);
    nor g3302(n28 ,n3160 ,n3096);
    nor g3303(n27 ,n3201 ,n3137);
    nor g3304(n26 ,n3158 ,n3094);
    nor g3305(n25 ,n3192 ,n3128);
    nor g3306(n24 ,n3157 ,n3093);
    nor g3307(n23 ,n3185 ,n3121);
    nor g3308(n22 ,n3167 ,n3103);
    nor g3309(n21 ,n3200 ,n3136);
    nor g3310(n20 ,n3168 ,n3104);
    nor g3311(n19 ,n3153 ,n3089);
    nor g3312(n18 ,n3175 ,n3111);
    nor g3313(n17 ,n3186 ,n3122);
    nor g3314(n16 ,n3207 ,n3143);
    nor g3315(n15 ,n3181 ,n3117);
    nor g3316(n14 ,n3199 ,n3135);
    not g3317(n13 ,n3152);
    not g3318(n12 ,n3154);
    not g3319(n11 ,n3090);
    not g3320(n10 ,n3088);
    xor g3321(n3216 ,n8[7] ,n290);
    nor g3322(n3217 ,n289 ,n290);
    nor g3323(n290 ,n267 ,n288);
    nor g3324(n289 ,n8[6] ,n287);
    nor g3325(n3218 ,n286 ,n287);
    not g3326(n288 ,n287);
    nor g3327(n287 ,n272 ,n285);
    nor g3328(n286 ,n8[5] ,n284);
    nor g3329(n3219 ,n283 ,n284);
    not g3330(n285 ,n284);
    nor g3331(n284 ,n269 ,n282);
    nor g3332(n283 ,n8[4] ,n281);
    nor g3333(n3220 ,n280 ,n281);
    not g3334(n282 ,n281);
    nor g3335(n281 ,n270 ,n279);
    nor g3336(n280 ,n8[3] ,n278);
    nor g3337(n3221 ,n277 ,n278);
    not g3338(n279 ,n278);
    nor g3339(n278 ,n273 ,n276);
    nor g3340(n277 ,n8[2] ,n275);
    nor g3341(n3222 ,n275 ,n274);
    not g3342(n276 ,n275);
    nor g3343(n275 ,n271 ,n268);
    nor g3344(n274 ,n8[1] ,n8[0]);
    not g3345(n273 ,n8[2]);
    not g3346(n272 ,n8[5]);
    not g3347(n271 ,n8[1]);
    not g3348(n270 ,n8[3]);
    not g3349(n269 ,n8[4]);
    not g3350(n268 ,n8[0]);
    not g3351(n267 ,n8[6]);
    xor g3352(n3023 ,n3589 ,n4[63]);
    xor g3353(n3022 ,n4[62] ,n3587);
    xor g3354(n3021 ,n4[61] ,n3586);
    nor g3355(n3589 ,n3316 ,n3588);
    not g3356(n3588 ,n3587);
    nor g3357(n3587 ,n3320 ,n3585);
    nor g3358(n3586 ,n3296 ,n3585);
    xnor g3359(n3020 ,n4[60] ,n3584);
    or g3360(n3585 ,n3299 ,n3584);
    xnor g3361(n3019 ,n4[59] ,n3581);
    nor g3362(n3584 ,n3583 ,n3582);
    xnor g3363(n3018 ,n4[58] ,n3576);
    nor g3364(n3583 ,n3271 ,n3580);
    nor g3365(n3582 ,n4[59] ,n3578);
    nor g3366(n3581 ,n3579 ,n3577);
    xnor g3367(n3017 ,n4[57] ,n3571);
    not g3368(n3580 ,n3579);
    nor g3369(n3579 ,n3267 ,n3575);
    not g3370(n3578 ,n3577);
    nor g3371(n3577 ,n4[58] ,n3573);
    nor g3372(n3576 ,n3574 ,n3572);
    not g3373(n3575 ,n3574);
    nor g3374(n3574 ,n3268 ,n3570);
    not g3375(n3573 ,n3572);
    nor g3376(n3572 ,n4[57] ,n3568);
    nor g3377(n3571 ,n3569 ,n3567);
    xnor g3378(n3016 ,n3319 ,n3565);
    not g3379(n3570 ,n3569);
    nor g3380(n3569 ,n3304 ,n3566);
    not g3381(n3568 ,n3567);
    nor g3382(n3567 ,n3290 ,n3565);
    not g3383(n3566 ,n3565);
    nor g3384(n3565 ,n3563 ,n3564);
    xnor g3385(n3015 ,n4[55] ,n3561);
    nor g3386(n3564 ,n3225 ,n3562);
    nor g3387(n3563 ,n4[55] ,n3561);
    xnor g3388(n3014 ,n4[54] ,n3557);
    xor g3389(n3013 ,n4[53] ,n3559);
    not g3390(n3562 ,n3561);
    nor g3391(n3561 ,n3560 ,n3558);
    xor g3392(n3012 ,n4[52] ,n3550);
    nor g3393(n3560 ,n3231 ,n3556);
    nor g3394(n3559 ,n3322 ,n3551);
    nor g3395(n3558 ,n4[54] ,n3553);
    nor g3396(n3557 ,n3555 ,n3552);
    or g3397(n3011 ,n3554 ,n3549);
    not g3398(n3556 ,n3555);
    nor g3399(n3555 ,n3303 ,n3548);
    nor g3400(n3554 ,n3539 ,n3547);
    not g3401(n3553 ,n3552);
    nor g3402(n3552 ,n4[53] ,n3545);
    not g3403(n3551 ,n3550);
    nor g3404(n3550 ,n3546 ,n3544);
    nor g3405(n3549 ,n4[51] ,n3543);
    xnor g3406(n3010 ,n4[50] ,n3538);
    or g3407(n3548 ,n3235 ,n3542);
    not g3408(n3547 ,n3546);
    nor g3409(n3546 ,n3259 ,n3541);
    or g3410(n3545 ,n3289 ,n3540);
    nor g3411(n3544 ,n4[51] ,n3539);
    nor g3412(n3543 ,n3541 ,n3539);
    xnor g3413(n3009 ,n4[49] ,n3533);
    not g3414(n3542 ,n3541);
    nor g3415(n3541 ,n3263 ,n3537);
    not g3416(n3540 ,n3539);
    nor g3417(n3539 ,n4[50] ,n3535);
    nor g3418(n3538 ,n3536 ,n3534);
    xnor g3419(n3008 ,n7[55] ,n3528);
    not g3420(n3537 ,n3536);
    nor g3421(n3536 ,n3266 ,n3532);
    not g3422(n3535 ,n3534);
    nor g3423(n3534 ,n4[49] ,n3530);
    nor g3424(n3533 ,n3531 ,n3529);
    not g3425(n3532 ,n3531);
    nor g3426(n3531 ,n3225 ,n3527);
    not g3427(n3530 ,n3529);
    nor g3428(n3529 ,n7[55] ,n3526);
    xor g3429(n3528 ,n4[48] ,n3524);
    or g3430(n3527 ,n3252 ,n3525);
    or g3431(n3526 ,n4[48] ,n3524);
    xor g3432(n3007 ,n4[47] ,n3522);
    not g3433(n3525 ,n3524);
    nor g3434(n3524 ,n3523 ,n3521);
    nor g3435(n3523 ,n3254 ,n3520);
    nor g3436(n3522 ,n3298 ,n3519);
    nor g3437(n3521 ,n4[47] ,n3519);
    xnor g3438(n3006 ,n4[46] ,n3518);
    nor g3439(n3520 ,n3262 ,n3518);
    or g3440(n3519 ,n3306 ,n3518);
    xnor g3441(n3005 ,n4[45] ,n3515);
    nor g3442(n3518 ,n3517 ,n3516);
    xnor g3443(n3004 ,n4[44] ,n3510);
    nor g3444(n3517 ,n3239 ,n3514);
    nor g3445(n3516 ,n4[45] ,n3512);
    nor g3446(n3515 ,n3513 ,n3511);
    xnor g3447(n3003 ,n4[43] ,n3505);
    not g3448(n3514 ,n3513);
    nor g3449(n3513 ,n3265 ,n3509);
    not g3450(n3512 ,n3511);
    nor g3451(n3511 ,n4[44] ,n3507);
    nor g3452(n3510 ,n3508 ,n3506);
    xnor g3453(n3002 ,n4[42] ,n3500);
    not g3454(n3509 ,n3508);
    nor g3455(n3508 ,n3272 ,n3504);
    not g3456(n3507 ,n3506);
    nor g3457(n3506 ,n4[43] ,n3502);
    nor g3458(n3505 ,n3503 ,n3501);
    xnor g3459(n3001 ,n4[41] ,n3495);
    not g3460(n3504 ,n3503);
    nor g3461(n3503 ,n3228 ,n3499);
    not g3462(n3502 ,n3501);
    nor g3463(n3501 ,n4[42] ,n3497);
    nor g3464(n3500 ,n3498 ,n3496);
    xnor g3465(n3000 ,n7[47] ,n3490);
    not g3466(n3499 ,n3498);
    nor g3467(n3498 ,n3270 ,n3494);
    not g3468(n3497 ,n3496);
    nor g3469(n3496 ,n4[41] ,n3492);
    nor g3470(n3495 ,n3493 ,n3491);
    not g3471(n3494 ,n3493);
    nor g3472(n3493 ,n3254 ,n3489);
    not g3473(n3492 ,n3491);
    nor g3474(n3491 ,n7[47] ,n3488);
    xor g3475(n3490 ,n4[40] ,n3484);
    or g3476(n3489 ,n3282 ,n3485);
    or g3477(n2999 ,n3487 ,n3486);
    or g3478(n3488 ,n4[40] ,n3484);
    nor g3479(n3487 ,n3287 ,n3482);
    nor g3480(n3486 ,n3312 ,n3481);
    not g3481(n3485 ,n3484);
    nor g3482(n3484 ,n3483 ,n3480);
    nor g3483(n3483 ,n3257 ,n3479);
    nor g3484(n3482 ,n3312 ,n3478);
    not g3485(n3481 ,n3480);
    nor g3486(n3480 ,n4[39] ,n3478);
    xnor g3487(n2998 ,n4[38] ,n3477);
    nor g3488(n3479 ,n3234 ,n3477);
    or g3489(n3478 ,n3309 ,n3477);
    xnor g3490(n2997 ,n4[37] ,n3474);
    nor g3491(n3477 ,n3476 ,n3475);
    xnor g3492(n2996 ,n4[36] ,n3469);
    nor g3493(n3476 ,n3240 ,n3473);
    nor g3494(n3475 ,n4[37] ,n3471);
    nor g3495(n3474 ,n3472 ,n3470);
    xnor g3496(n2995 ,n4[35] ,n3464);
    not g3497(n3473 ,n3472);
    nor g3498(n3472 ,n3274 ,n3468);
    not g3499(n3471 ,n3470);
    nor g3500(n3470 ,n4[36] ,n3466);
    nor g3501(n3469 ,n3467 ,n3465);
    xnor g3502(n2994 ,n4[34] ,n3459);
    not g3503(n3468 ,n3467);
    nor g3504(n3467 ,n3236 ,n3463);
    not g3505(n3466 ,n3465);
    nor g3506(n3465 ,n4[35] ,n3461);
    nor g3507(n3464 ,n3462 ,n3460);
    xnor g3508(n2993 ,n4[33] ,n3454);
    not g3509(n3463 ,n3462);
    nor g3510(n3462 ,n3233 ,n3458);
    not g3511(n3461 ,n3460);
    nor g3512(n3460 ,n4[34] ,n3456);
    nor g3513(n3459 ,n3457 ,n3455);
    not g3514(n3458 ,n3457);
    nor g3515(n3457 ,n3277 ,n3453);
    not g3516(n3456 ,n3455);
    nor g3517(n3455 ,n4[33] ,n3451);
    nor g3518(n3454 ,n3452 ,n3450);
    xnor g3519(n2992 ,n3313 ,n3448);
    not g3520(n3453 ,n3452);
    nor g3521(n3452 ,n3302 ,n3449);
    not g3522(n3451 ,n3450);
    nor g3523(n3450 ,n3293 ,n3448);
    not g3524(n3449 ,n3448);
    nor g3525(n3448 ,n3447 ,n3446);
    xor g3526(n2991 ,n4[31] ,n3443);
    nor g3527(n3447 ,n3224 ,n3445);
    nor g3528(n3446 ,n4[31] ,n3444);
    xnor g3529(n2990 ,n4[30] ,n3442);
    nor g3530(n3445 ,n3264 ,n3442);
    not g3531(n3444 ,n3443);
    nor g3532(n3443 ,n3318 ,n3442);
    xnor g3533(n2989 ,n4[29] ,n3439);
    nor g3534(n3442 ,n3441 ,n3440);
    xnor g3535(n2988 ,n4[28] ,n3434);
    nor g3536(n3441 ,n3243 ,n3438);
    nor g3537(n3440 ,n4[29] ,n3436);
    nor g3538(n3439 ,n3437 ,n3435);
    xnor g3539(n2987 ,n4[27] ,n3429);
    not g3540(n3438 ,n3437);
    nor g3541(n3437 ,n3280 ,n3433);
    not g3542(n3436 ,n3435);
    nor g3543(n3435 ,n4[28] ,n3431);
    nor g3544(n3434 ,n3432 ,n3430);
    xnor g3545(n2986 ,n4[26] ,n3424);
    not g3546(n3433 ,n3432);
    nor g3547(n3432 ,n3232 ,n3428);
    not g3548(n3431 ,n3430);
    nor g3549(n3430 ,n4[27] ,n3426);
    nor g3550(n3429 ,n3427 ,n3425);
    xnor g3551(n2985 ,n4[25] ,n3419);
    not g3552(n3428 ,n3427);
    nor g3553(n3427 ,n3261 ,n3423);
    not g3554(n3426 ,n3425);
    nor g3555(n3425 ,n4[26] ,n3421);
    nor g3556(n3424 ,n3422 ,n3420);
    not g3557(n3423 ,n3422);
    nor g3558(n3422 ,n3237 ,n3418);
    not g3559(n3421 ,n3420);
    nor g3560(n3420 ,n4[25] ,n3416);
    nor g3561(n3419 ,n3417 ,n3415);
    xnor g3562(n2984 ,n3314 ,n3413);
    not g3563(n3418 ,n3417);
    nor g3564(n3417 ,n3301 ,n3414);
    not g3565(n3416 ,n3415);
    nor g3566(n3415 ,n3292 ,n3413);
    not g3567(n3414 ,n3413);
    nor g3568(n3413 ,n3411 ,n3412);
    xnor g3569(n2983 ,n4[23] ,n3409);
    nor g3570(n3412 ,n3260 ,n3410);
    nor g3571(n3411 ,n4[23] ,n3409);
    xnor g3572(n2981 ,n3405 ,n3399);
    xnor g3573(n2982 ,n4[22] ,n3406);
    not g3574(n3410 ,n3409);
    nor g3575(n3409 ,n3408 ,n3407);
    nor g3576(n3408 ,n3241 ,n3404);
    nor g3577(n3407 ,n4[22] ,n3402);
    nor g3578(n3406 ,n3403 ,n3401);
    xnor g3579(n3405 ,n4[21] ,n3397);
    xnor g3580(n2980 ,n4[20] ,n3396);
    not g3581(n3404 ,n3403);
    nor g3582(n3403 ,n3244 ,n3400);
    not g3583(n3402 ,n3401);
    nor g3584(n3401 ,n4[21] ,n3398);
    xnor g3585(n2979 ,n4[19] ,n3391);
    not g3586(n3400 ,n3399);
    nor g3587(n3399 ,n3273 ,n3395);
    not g3588(n3398 ,n3397);
    nor g3589(n3397 ,n4[20] ,n3393);
    nor g3590(n3396 ,n3394 ,n3392);
    xnor g3591(n2978 ,n4[18] ,n3386);
    not g3592(n3395 ,n3394);
    nor g3593(n3394 ,n3230 ,n3390);
    not g3594(n3393 ,n3392);
    nor g3595(n3392 ,n4[19] ,n3388);
    nor g3596(n3391 ,n3389 ,n3387);
    xnor g3597(n2977 ,n4[17] ,n3381);
    not g3598(n3390 ,n3389);
    nor g3599(n3389 ,n3227 ,n3385);
    not g3600(n3388 ,n3387);
    nor g3601(n3387 ,n4[18] ,n3383);
    nor g3602(n3386 ,n3384 ,n3382);
    xnor g3603(n2976 ,n7[23] ,n3376);
    not g3604(n3385 ,n3384);
    nor g3605(n3384 ,n3275 ,n3380);
    not g3606(n3383 ,n3382);
    nor g3607(n3382 ,n4[17] ,n3378);
    nor g3608(n3381 ,n3379 ,n3377);
    not g3609(n3380 ,n3379);
    nor g3610(n3379 ,n3260 ,n3375);
    not g3611(n3378 ,n3377);
    nor g3612(n3377 ,n7[23] ,n3374);
    xor g3613(n3376 ,n4[16] ,n3372);
    or g3614(n3375 ,n3246 ,n3373);
    or g3615(n3374 ,n4[16] ,n3372);
    not g3616(n3373 ,n3372);
    nor g3617(n3372 ,n3368 ,n3371);
    xor g3618(n2975 ,n4[15] ,n3369);
    nor g3619(n3371 ,n3223 ,n3370);
    xor g3620(n2974 ,n4[14] ,n3364);
    nor g3621(n3370 ,n3305 ,n3367);
    nor g3622(n3369 ,n3323 ,n3365);
    nor g3623(n3368 ,n4[15] ,n3366);
    xor g3624(n2973 ,n3362 ,n4[13]);
    xor g3625(n2972 ,n4[12] ,n3361);
    or g3626(n3367 ,n3238 ,n3363);
    or g3627(n3366 ,n3291 ,n3363);
    not g3628(n3365 ,n3364);
    nor g3629(n3364 ,n3315 ,n3363);
    not g3630(n3363 ,n3362);
    nor g3631(n3362 ,n3321 ,n3360);
    nor g3632(n3361 ,n3294 ,n3360);
    xnor g3633(n2971 ,n4[11] ,n3359);
    or g3634(n3360 ,n3297 ,n3359);
    xnor g3635(n2970 ,n4[10] ,n3356);
    nor g3636(n3359 ,n3358 ,n3357);
    xnor g3637(n2969 ,n4[9] ,n3351);
    nor g3638(n3358 ,n3269 ,n3355);
    nor g3639(n3357 ,n4[10] ,n3353);
    nor g3640(n3356 ,n3354 ,n3352);
    xnor g3641(n2968 ,n7[15] ,n3346);
    not g3642(n3355 ,n3354);
    nor g3643(n3354 ,n3279 ,n3350);
    not g3644(n3353 ,n3352);
    nor g3645(n3352 ,n4[9] ,n3348);
    nor g3646(n3351 ,n3349 ,n3347);
    not g3647(n3350 ,n3349);
    nor g3648(n3349 ,n3223 ,n3345);
    not g3649(n3348 ,n3347);
    nor g3650(n3347 ,n7[15] ,n3344);
    xnor g3651(n3346 ,n4[8] ,n3342);
    or g3652(n3345 ,n3288 ,n3342);
    or g3653(n3344 ,n4[8] ,n3343);
    not g3654(n3343 ,n3342);
    nor g3655(n3342 ,n3281 ,n3341);
    xor g3656(n2967 ,n4[7] ,n3339);
    nor g3657(n3341 ,n3249 ,n3340);
    nor g3658(n2966 ,n3338 ,n3339);
    not g3659(n3340 ,n3339);
    nor g3660(n3339 ,n3253 ,n3337);
    nor g3661(n3338 ,n4[6] ,n3336);
    nor g3662(n2965 ,n3335 ,n3336);
    not g3663(n3337 ,n3336);
    nor g3664(n3336 ,n3286 ,n3334);
    nor g3665(n3335 ,n4[5] ,n3333);
    nor g3666(n2964 ,n3332 ,n3333);
    not g3667(n3334 ,n3333);
    nor g3668(n3333 ,n3250 ,n3331);
    nor g3669(n3332 ,n4[4] ,n3330);
    nor g3670(n2963 ,n3329 ,n3330);
    not g3671(n3331 ,n3330);
    nor g3672(n3330 ,n3285 ,n3328);
    nor g3673(n3329 ,n4[3] ,n3327);
    nor g3674(n2962 ,n3326 ,n3327);
    not g3675(n3328 ,n3327);
    nor g3676(n3327 ,n3248 ,n3325);
    nor g3677(n3326 ,n4[2] ,n3324);
    nor g3678(n2961 ,n3317 ,n3324);
    not g3679(n3325 ,n3324);
    xor g3680(n3323 ,n4[13] ,n4[14]);
    xnor g3681(n3322 ,n3259 ,n4[52]);
    nor g3682(n3321 ,n3308 ,n3295);
    nor g3683(n3320 ,n3307 ,n3300);
    xor g3684(n3319 ,n7[63] ,n4[56]);
    nor g3685(n3324 ,n3284 ,n3311);
    xnor g3686(n3318 ,n3264 ,n7[31]);
    nor g3687(n3317 ,n4[1] ,n3310);
    xor g3688(n3316 ,n7[63] ,n4[62]);
    xnor g3689(n2960 ,n3281 ,n4[0]);
    xnor g3690(n3315 ,n3223 ,n4[13]);
    xnor g3691(n3314 ,n3224 ,n4[24]);
    xnor g3692(n3313 ,n3257 ,n4[32]);
    not g3693(n3311 ,n3310);
    nor g3694(n3309 ,n3234 ,n7[39]);
    nor g3695(n3308 ,n3242 ,n3223);
    nor g3696(n3307 ,n3276 ,n3255);
    nor g3697(n3306 ,n3262 ,n7[47]);
    or g3698(n3305 ,n3229 ,n3256);
    nor g3699(n3312 ,n3257 ,n4[38]);
    or g3700(n3304 ,n3245 ,n3255);
    or g3701(n3303 ,n3278 ,n3259);
    or g3702(n3302 ,n3283 ,n3257);
    or g3703(n3301 ,n3251 ,n3224);
    nor g3704(n3310 ,n3247 ,n3281);
    nor g3705(n3300 ,n4[61] ,n4[60]);
    nor g3706(n3299 ,n3255 ,n4[60]);
    nor g3707(n3298 ,n3254 ,n4[46]);
    nor g3708(n3297 ,n3223 ,n4[11]);
    nor g3709(n3296 ,n3226 ,n7[63]);
    nor g3710(n3295 ,n4[12] ,n4[11]);
    nor g3711(n3294 ,n3258 ,n7[15]);
    or g3712(n3293 ,n4[32] ,n7[39]);
    or g3713(n3292 ,n4[24] ,n7[31]);
    or g3714(n3291 ,n4[14] ,n4[13]);
    or g3715(n3290 ,n4[56] ,n7[63]);
    or g3716(n3289 ,n4[52] ,n4[51]);
    not g3717(n3288 ,n4[8]);
    not g3718(n3287 ,n4[39]);
    not g3719(n3286 ,n4[5]);
    not g3720(n3285 ,n4[3]);
    not g3721(n3284 ,n4[1]);
    not g3722(n3283 ,n4[32]);
    not g3723(n3282 ,n4[40]);
    not g3724(n3281 ,n7[7]);
    not g3725(n3280 ,n4[28]);
    not g3726(n3279 ,n4[9]);
    not g3727(n3278 ,n4[52]);
    not g3728(n3277 ,n4[33]);
    not g3729(n3276 ,n4[61]);
    not g3730(n3275 ,n4[17]);
    not g3731(n3274 ,n4[36]);
    not g3732(n3273 ,n4[20]);
    not g3733(n3272 ,n4[43]);
    not g3734(n3271 ,n4[59]);
    not g3735(n3270 ,n4[41]);
    not g3736(n3269 ,n4[10]);
    not g3737(n3268 ,n4[57]);
    not g3738(n3267 ,n4[58]);
    not g3739(n3266 ,n4[49]);
    not g3740(n3265 ,n4[44]);
    not g3741(n3264 ,n4[30]);
    not g3742(n3263 ,n4[50]);
    not g3743(n3262 ,n4[46]);
    not g3744(n3261 ,n4[26]);
    not g3745(n3260 ,n7[23]);
    not g3746(n3259 ,n4[51]);
    not g3747(n3258 ,n4[11]);
    not g3748(n3257 ,n7[39]);
    not g3749(n3256 ,n4[13]);
    not g3750(n3255 ,n7[63]);
    not g3751(n3254 ,n7[47]);
    not g3752(n3253 ,n4[6]);
    not g3753(n3252 ,n4[48]);
    not g3754(n3251 ,n4[24]);
    not g3755(n3250 ,n4[4]);
    not g3756(n3249 ,n4[7]);
    not g3757(n3248 ,n4[2]);
    not g3758(n3247 ,n4[0]);
    not g3759(n3246 ,n4[16]);
    not g3760(n3245 ,n4[56]);
    not g3761(n3244 ,n4[21]);
    not g3762(n3243 ,n4[29]);
    not g3763(n3242 ,n4[12]);
    not g3764(n3241 ,n4[22]);
    not g3765(n3240 ,n4[37]);
    not g3766(n3239 ,n4[45]);
    not g3767(n3238 ,n4[15]);
    not g3768(n3237 ,n4[25]);
    not g3769(n3236 ,n4[35]);
    not g3770(n3235 ,n4[53]);
    not g3771(n3234 ,n4[38]);
    not g3772(n3233 ,n4[34]);
    not g3773(n3232 ,n4[27]);
    not g3774(n3231 ,n4[54]);
    not g3775(n3230 ,n4[19]);
    not g3776(n3229 ,n4[14]);
    not g3777(n3228 ,n4[42]);
    not g3778(n3227 ,n4[18]);
    not g3779(n3226 ,n4[60]);
    not g3780(n3225 ,n7[55]);
    not g3781(n3224 ,n7[31]);
    not g3782(n3223 ,n7[15]);
    dff g3783(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3630), .Q(n9[19]));
    or g3784(n3630 ,n1 ,n3629);
    xor g3785(n3629 ,n3619 ,n3620);
    dff g3786(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3623), .Q(n7[23]));
    dff g3787(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3624), .Q(n7[15]));
    dff g3788(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3625), .Q(n7[7]));
    dff g3789(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3622), .Q(n7[31]));
    dff g3790(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3628), .Q(n7[55]));
    dff g3791(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3627), .Q(n7[47]));
    dff g3792(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3621), .Q(n7[39]));
    dff g3793(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3626), .Q(n7[63]));
    dff g3794(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3605), .Q(n9[16]));
    dff g3795(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3617), .Q(n9[18]));
    dff g3796(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3602), .Q(n9[8]));
    dff g3797(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3600), .Q(n9[12]));
    dff g3798(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3618), .Q(n9[14]));
    dff g3799(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3610), .Q(n9[17]));
    dff g3800(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3609), .Q(n9[6]));
    dff g3801(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3604), .Q(n9[11]));
    dff g3802(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3601), .Q(n9[3]));
    dff g3803(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3606), .Q(n9[4]));
    dff g3804(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3607), .Q(n9[15]));
    dff g3805(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3616), .Q(n9[5]));
    dff g3806(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3608), .Q(n9[0]));
    dff g3807(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3603), .Q(n9[7]));
    dff g3808(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3612), .Q(n9[9]));
    xor g3809(n3628 ,n9[6] ,n2[6]);
    xor g3810(n3627 ,n9[5] ,n2[5]);
    dff g3811(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3611), .Q(n9[13]));
    xor g3812(n3626 ,n9[7] ,n2[7]);
    dff g3813(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3614), .Q(n9[10]));
    xor g3814(n3625 ,n9[0] ,n2[0]);
    xor g3815(n3624 ,n9[1] ,n2[1]);
    xor g3816(n3623 ,n9[2] ,n2[2]);
    xor g3817(n3622 ,n9[3] ,n2[3]);
    xor g3818(n3621 ,n9[4] ,n2[4]);
    xnor g3819(n3620 ,n9[7] ,n9[0]);
    xnor g3820(n3619 ,n9[11] ,n9[15]);
    dff g3821(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3613), .Q(n9[2]));
    dff g3822(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3615), .Q(n9[1]));
    nor g3823(n3618 ,n3591 ,n1);
    nor g3824(n3617 ,n3599 ,n1);
    nor g3825(n3616 ,n3596 ,n1);
    nor g3826(n3615 ,n3592 ,n1);
    nor g3827(n3614 ,n3595 ,n1);
    nor g3828(n3613 ,n3594 ,n1);
    nor g3829(n3612 ,n3597 ,n1);
    nor g3830(n3611 ,n3593 ,n1);
    nor g3831(n3610 ,n3598 ,n1);
    nor g3832(n3609 ,n3590 ,n1);
    or g3833(n3608 ,n9[1] ,n1);
    or g3834(n3607 ,n9[16] ,n1);
    or g3835(n3606 ,n9[5] ,n1);
    or g3836(n3605 ,n9[17] ,n1);
    or g3837(n3604 ,n9[12] ,n1);
    or g3838(n3603 ,n9[8] ,n1);
    or g3839(n3602 ,n9[9] ,n1);
    or g3840(n3601 ,n9[4] ,n1);
    or g3841(n3600 ,n9[13] ,n1);
    not g3842(n3599 ,n9[19]);
    not g3843(n3598 ,n9[18]);
    not g3844(n3597 ,n9[10]);
    not g3845(n3596 ,n9[6]);
    not g3846(n3595 ,n9[11]);
    not g3847(n3594 ,n9[3]);
    not g3848(n3593 ,n9[14]);
    not g3849(n3592 ,n9[2]);
    not g3850(n3591 ,n9[15]);
    not g3851(n3590 ,n9[7]);
endmodule
