module top(n0, n1, n2, n3, n4, n5, n6);
    input n0, n1;
    input [13:0] n2;
    input [12:0] n3;
    output [12:0] n4, n5, n6;
    wire n0, n1;
    wire [13:0] n2;
    wire [12:0] n3;
    wire [12:0] n4, n5, n6;
    wire [12:0] n7;
    wire [12:0] n8;
    wire [12:0] n9;
    wire [12:0] n10;
    wire [12:0] n11;
    wire [12:0] n12;
    wire [2:0] n13;
    wire [3:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848;
    not g0(n706 ,n7[11]);
    not g1(n705 ,n7[5]);
    not g2(n704 ,n7[10]);
    not g3(n703 ,n7[8]);
    not g4(n702 ,n7[2]);
    not g5(n701 ,n7[9]);
    not g6(n700 ,n7[4]);
    not g7(n699 ,n7[1]);
    not g8(n698 ,n7[7]);
    not g9(n697 ,n7[0]);
    not g10(n696 ,n7[12]);
    not g11(n695 ,n7[6]);
    not g12(n694 ,n7[3]);
    xnor g13(n5[3] ,n688 ,n8[3]);
    xnor g14(n4[10] ,n687 ,n9[10]);
    xnor g15(n4[9] ,n692 ,n9[9]);
    xnor g16(n4[6] ,n691 ,n9[6]);
    xnor g17(n4[5] ,n693 ,n9[5]);
    xnor g18(n5[11] ,n686 ,n8[11]);
    xnor g19(n5[10] ,n687 ,n8[10]);
    xnor g20(n5[9] ,n692 ,n8[9]);
    xnor g21(n5[8] ,n689 ,n8[8]);
    xnor g22(n4[8] ,n689 ,n9[8]);
    xnor g23(n5[7] ,n684 ,n8[7]);
    xnor g24(n5[6] ,n691 ,n8[6]);
    xnor g25(n5[5] ,n693 ,n8[5]);
    xnor g26(n5[4] ,n690 ,n8[4]);
    xnor g27(n4[4] ,n690 ,n9[4]);
    xnor g28(n4[11] ,n686 ,n9[11]);
    xnor g29(n5[2] ,n685 ,n8[2]);
    xnor g30(n5[1] ,n683 ,n8[1]);
    xnor g31(n4[7] ,n684 ,n9[7]);
    xnor g32(n4[3] ,n688 ,n9[3]);
    xnor g33(n6[11] ,n686 ,n10[11]);
    xnor g34(n6[10] ,n687 ,n10[10]);
    xnor g35(n6[9] ,n692 ,n10[9]);
    xnor g36(n4[2] ,n685 ,n9[2]);
    xnor g37(n6[8] ,n689 ,n10[8]);
    xnor g38(n6[7] ,n684 ,n10[7]);
    xnor g39(n6[6] ,n691 ,n10[6]);
    xnor g40(n6[5] ,n693 ,n10[5]);
    xnor g41(n4[1] ,n683 ,n9[1]);
    xnor g42(n6[4] ,n690 ,n10[4]);
    xnor g43(n6[3] ,n688 ,n10[3]);
    xnor g44(n6[2] ,n685 ,n10[2]);
    xnor g45(n6[1] ,n683 ,n10[1]);
    xnor g46(n4[0] ,n681 ,n9[0]);
    xnor g47(n5[12] ,n682 ,n8[12]);
    xnor g48(n5[0] ,n681 ,n8[0]);
    xnor g49(n6[12] ,n682 ,n10[12]);
    xnor g50(n4[12] ,n682 ,n9[12]);
    xnor g51(n6[0] ,n681 ,n10[0]);
    xnor g52(n693 ,n11[5] ,n679);
    xnor g53(n692 ,n11[9] ,n680);
    xnor g54(n691 ,n11[6] ,n670);
    xnor g55(n690 ,n11[4] ,n678);
    xnor g56(n689 ,n11[8] ,n677);
    xnor g57(n688 ,n11[3] ,n676);
    xnor g58(n687 ,n11[10] ,n675);
    xnor g59(n686 ,n11[11] ,n671);
    xnor g60(n685 ,n11[2] ,n674);
    xnor g61(n684 ,n11[7] ,n673);
    xnor g62(n683 ,n11[1] ,n672);
    xnor g63(n682 ,n11[12] ,n664);
    xnor g64(n681 ,n3[0] ,n665);
    xor g65(n764 ,n11[9] ,n3[9]);
    xor g66(n763 ,n11[8] ,n3[8]);
    xor g67(n762 ,n11[7] ,n3[7]);
    xor g68(n761 ,n11[6] ,n3[6]);
    xor g69(n759 ,n11[4] ,n3[4]);
    xor g70(n758 ,n11[3] ,n3[3]);
    xor g71(n757 ,n11[2] ,n3[2]);
    xor g72(n756 ,n11[1] ,n3[1]);
    xor g73(n789 ,n11[8] ,n2[8]);
    xor g74(n788 ,n11[7] ,n2[7]);
    xor g75(n740 ,n11[11] ,n741);
    xor g76(n738 ,n11[10] ,n739);
    xor g77(n736 ,n11[9] ,n737);
    nor g78(n680 ,n701 ,n666);
    nor g79(n679 ,n705 ,n657);
    nor g80(n678 ,n700 ,n662);
    nor g81(n677 ,n703 ,n661);
    nor g82(n676 ,n694 ,n660);
    nor g83(n675 ,n704 ,n658);
    nor g84(n674 ,n702 ,n659);
    nor g85(n673 ,n698 ,n663);
    nor g86(n672 ,n699 ,n669);
    nor g87(n671 ,n706 ,n668);
    nor g88(n670 ,n695 ,n667);
    xor g89(n734 ,n11[8] ,n735);
    xor g90(n732 ,n11[7] ,n733);
    xor g91(n730 ,n11[6] ,n731);
    xor g92(n728 ,n11[5] ,n729);
    xor g93(n726 ,n11[4] ,n727);
    xor g94(n724 ,n11[3] ,n725);
    xor g95(n722 ,n11[2] ,n723);
    xor g96(n720 ,n11[1] ,n721);
    xor g97(n792 ,n11[11] ,n2[11]);
    xor g98(n791 ,n11[10] ,n2[10]);
    xor g99(n790 ,n11[9] ,n2[9]);
    xor g100(n783 ,n11[2] ,n2[2]);
    xor g101(n787 ,n11[6] ,n2[6]);
    xor g102(n785 ,n11[4] ,n2[4]);
    xor g103(n784 ,n11[3] ,n2[3]);
    xor g104(n782 ,n11[1] ,n2[1]);
    xor g105(n786 ,n11[5] ,n2[5]);
    xor g106(n760 ,n11[5] ,n3[5]);
    xor g107(n766 ,n11[11] ,n3[11]);
    xor g108(n765 ,n11[10] ,n3[10]);
    xor g109(n742 ,n11[12] ,n743);
    xor g110(n793 ,n11[12] ,n2[12]);
    xor g111(n767 ,n11[12] ,n3[12]);
    xor g112(n781 ,n2[0] ,n3[0]);
    not g113(n12[1] ,n669);
    not g114(n12[11] ,n668);
    not g115(n12[6] ,n667);
    not g116(n12[9] ,n666);
    nor g117(n665 ,n656 ,n697);
    nor g118(n664 ,n655 ,n696);
    nor g119(n669 ,n3[0] ,n11[2]);
    nor g120(n668 ,n11[12] ,n11[10]);
    nor g121(n667 ,n11[7] ,n11[5]);
    nor g122(n666 ,n11[10] ,n11[8]);
    not g123(n12[7] ,n663);
    not g124(n12[4] ,n662);
    not g125(n12[8] ,n661);
    not g126(n12[3] ,n660);
    not g127(n12[2] ,n659);
    not g128(n12[10] ,n658);
    not g129(n12[5] ,n657);
    nor g130(n663 ,n11[8] ,n11[6]);
    nor g131(n662 ,n11[5] ,n11[3]);
    nor g132(n661 ,n11[9] ,n11[7]);
    nor g133(n660 ,n11[4] ,n11[2]);
    nor g134(n659 ,n11[3] ,n11[1]);
    nor g135(n658 ,n11[11] ,n11[9]);
    nor g136(n657 ,n11[6] ,n11[4]);
    not g137(n656 ,n11[1]);
    not g138(n655 ,n11[11]);
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n594), .Q(n9[0]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n570), .Q(n9[1]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n603), .Q(n9[2]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n597), .Q(n9[3]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n596), .Q(n9[4]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n587), .Q(n9[5]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n586), .Q(n9[6]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n581), .Q(n9[7]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n580), .Q(n9[8]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n579), .Q(n9[9]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n9[10]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n578), .Q(n9[11]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n577), .Q(n9[12]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n576), .Q(n8[0]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n601), .Q(n8[1]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n574), .Q(n8[2]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n573), .Q(n8[3]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n572), .Q(n8[4]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n571), .Q(n8[5]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n602), .Q(n8[6]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n616), .Q(n8[7]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n631), .Q(n8[8]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n567), .Q(n8[9]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n600), .Q(n8[10]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n599), .Q(n8[11]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n598), .Q(n8[12]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n640), .Q(n10[0]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n568), .Q(n10[1]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n595), .Q(n10[2]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n593), .Q(n10[3]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n592), .Q(n10[4]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n591), .Q(n10[5]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n590), .Q(n10[6]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n589), .Q(n10[7]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n588), .Q(n10[8]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n585), .Q(n10[9]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n584), .Q(n10[10]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n583), .Q(n10[11]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n582), .Q(n10[12]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n646), .Q(n7[0]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n645), .Q(n7[1]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n644), .Q(n7[2]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n643), .Q(n7[3]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n642), .Q(n7[4]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n641), .Q(n7[5]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n647), .Q(n7[6]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n639), .Q(n7[7]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n638), .Q(n7[8]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n637), .Q(n7[9]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n636), .Q(n7[10]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n635), .Q(n7[11]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n634), .Q(n7[12]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n496), .Q(n13[0]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n495), .Q(n13[1]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n13[2]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n654), .Q(n14[0]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n653), .Q(n14[1]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n652), .Q(n14[2]));
    nor g197(n654 ,n1 ,n651);
    nor g198(n653 ,n1 ,n650);
    nor g199(n652 ,n1 ,n648);
    or g200(n651 ,n364 ,n649);
    or g201(n650 ,n373 ,n649);
    not g202(n648 ,n649);
    nor g203(n649 ,n369 ,n633);
    or g204(n647 ,n618 ,n617);
    or g205(n646 ,n629 ,n628);
    or g206(n645 ,n626 ,n627);
    or g207(n644 ,n625 ,n624);
    or g208(n643 ,n622 ,n623);
    or g209(n642 ,n619 ,n621);
    or g210(n641 ,n630 ,n620);
    or g211(n640 ,n557 ,n569);
    or g212(n639 ,n615 ,n632);
    or g213(n638 ,n614 ,n613);
    or g214(n637 ,n611 ,n612);
    or g215(n636 ,n610 ,n609);
    or g216(n635 ,n607 ,n608);
    or g217(n634 ,n605 ,n606);
    nor g218(n633 ,n14[0] ,n604);
    nor g219(n632 ,n259 ,n566);
    or g220(n631 ,n563 ,n523);
    nor g221(n630 ,n307 ,n526);
    nor g222(n629 ,n317 ,n526);
    nor g223(n628 ,n251 ,n566);
    nor g224(n627 ,n262 ,n566);
    nor g225(n626 ,n313 ,n526);
    nor g226(n625 ,n319 ,n526);
    nor g227(n624 ,n257 ,n566);
    nor g228(n623 ,n254 ,n566);
    nor g229(n622 ,n312 ,n526);
    nor g230(n621 ,n255 ,n566);
    nor g231(n620 ,n264 ,n566);
    nor g232(n619 ,n315 ,n526);
    nor g233(n618 ,n309 ,n526);
    nor g234(n617 ,n252 ,n566);
    or g235(n616 ,n564 ,n524);
    nor g236(n615 ,n318 ,n526);
    nor g237(n614 ,n310 ,n526);
    nor g238(n613 ,n260 ,n566);
    nor g239(n612 ,n258 ,n566);
    nor g240(n611 ,n311 ,n526);
    nor g241(n610 ,n316 ,n526);
    nor g242(n609 ,n253 ,n566);
    nor g243(n608 ,n261 ,n566);
    nor g244(n607 ,n314 ,n526);
    nor g245(n606 ,n265 ,n566);
    nor g246(n605 ,n306 ,n526);
    nor g247(n604 ,n360 ,n529);
    or g248(n603 ,n560 ,n517);
    or g249(n602 ,n545 ,n527);
    or g250(n601 ,n427 ,n489);
    or g251(n600 ,n561 ,n519);
    or g252(n599 ,n559 ,n518);
    or g253(n598 ,n558 ,n516);
    or g254(n597 ,n556 ,n515);
    or g255(n596 ,n553 ,n511);
    or g256(n595 ,n555 ,n513);
    or g257(n594 ,n538 ,n491);
    or g258(n593 ,n554 ,n512);
    or g259(n592 ,n552 ,n490);
    or g260(n591 ,n551 ,n510);
    or g261(n590 ,n549 ,n509);
    or g262(n589 ,n548 ,n507);
    or g263(n588 ,n547 ,n506);
    or g264(n587 ,n550 ,n508);
    or g265(n586 ,n565 ,n504);
    or g266(n585 ,n546 ,n505);
    or g267(n584 ,n544 ,n522);
    or g268(n583 ,n543 ,n503);
    or g269(n582 ,n542 ,n502);
    or g270(n581 ,n541 ,n500);
    or g271(n580 ,n540 ,n498);
    or g272(n579 ,n539 ,n497);
    or g273(n578 ,n536 ,n494);
    or g274(n577 ,n535 ,n493);
    or g275(n576 ,n534 ,n492);
    or g276(n575 ,n537 ,n499);
    or g277(n574 ,n533 ,n488);
    or g278(n573 ,n532 ,n487);
    or g279(n572 ,n531 ,n486);
    or g280(n571 ,n530 ,n501);
    or g281(n570 ,n459 ,n521);
    or g282(n569 ,n479 ,n528);
    or g283(n568 ,n452 ,n514);
    or g284(n567 ,n562 ,n520);
    nor g285(n565 ,n323 ,n435);
    nor g286(n564 ,n357 ,n447);
    nor g287(n563 ,n352 ,n446);
    nor g288(n562 ,n356 ,n442);
    nor g289(n561 ,n333 ,n443);
    nor g290(n560 ,n343 ,n440);
    nor g291(n559 ,n263 ,n441);
    nor g292(n558 ,n331 ,n439);
    nor g293(n557 ,n346 ,n436);
    nor g294(n556 ,n341 ,n438);
    nor g295(n555 ,n340 ,n440);
    nor g296(n554 ,n332 ,n438);
    nor g297(n553 ,n335 ,n444);
    nor g298(n552 ,n349 ,n444);
    nor g299(n551 ,n324 ,n445);
    nor g300(n550 ,n344 ,n445);
    nor g301(n549 ,n327 ,n435);
    nor g302(n548 ,n330 ,n447);
    nor g303(n547 ,n338 ,n446);
    nor g304(n546 ,n348 ,n442);
    nor g305(n545 ,n325 ,n435);
    nor g306(n544 ,n326 ,n443);
    nor g307(n543 ,n353 ,n441);
    nor g308(n542 ,n350 ,n439);
    nor g309(n541 ,n329 ,n447);
    nor g310(n540 ,n334 ,n446);
    nor g311(n539 ,n355 ,n442);
    nor g312(n538 ,n347 ,n436);
    nor g313(n537 ,n336 ,n443);
    nor g314(n536 ,n342 ,n441);
    nor g315(n535 ,n328 ,n439);
    nor g316(n534 ,n339 ,n436);
    nor g317(n533 ,n351 ,n440);
    nor g318(n532 ,n354 ,n438);
    nor g319(n531 ,n345 ,n444);
    nor g320(n530 ,n337 ,n445);
    or g321(n529 ,n377 ,n420);
    nor g322(n528 ,n367 ,n419);
    or g323(n527 ,n461 ,n478);
    or g324(n566 ,n1 ,n449);
    nor g325(n525 ,n1 ,n415);
    or g326(n524 ,n460 ,n485);
    or g327(n523 ,n458 ,n480);
    or g328(n522 ,n473 ,n482);
    nor g329(n521 ,n418 ,n437);
    or g330(n520 ,n467 ,n481);
    or g331(n519 ,n456 ,n482);
    or g332(n518 ,n430 ,n483);
    or g333(n517 ,n453 ,n474);
    or g334(n516 ,n454 ,n484);
    or g335(n515 ,n450 ,n476);
    nor g336(n514 ,n416 ,n437);
    or g337(n513 ,n457 ,n474);
    or g338(n512 ,n455 ,n476);
    or g339(n511 ,n464 ,n477);
    or g340(n510 ,n465 ,n475);
    or g341(n509 ,n466 ,n478);
    or g342(n508 ,n462 ,n475);
    or g343(n507 ,n469 ,n485);
    or g344(n506 ,n468 ,n480);
    or g345(n505 ,n451 ,n481);
    or g346(n504 ,n471 ,n478);
    or g347(n503 ,n470 ,n483);
    or g348(n502 ,n472 ,n484);
    or g349(n501 ,n422 ,n475);
    or g350(n500 ,n417 ,n485);
    or g351(n499 ,n433 ,n482);
    or g352(n498 ,n421 ,n480);
    or g353(n497 ,n432 ,n481);
    nor g354(n496 ,n1 ,n434);
    nor g355(n495 ,n1 ,n413);
    or g356(n494 ,n431 ,n483);
    or g357(n493 ,n429 ,n484);
    or g358(n492 ,n428 ,n479);
    or g359(n491 ,n426 ,n479);
    or g360(n490 ,n463 ,n477);
    nor g361(n489 ,n414 ,n437);
    or g362(n488 ,n425 ,n474);
    or g363(n487 ,n424 ,n476);
    or g364(n486 ,n423 ,n477);
    or g365(n526 ,n1 ,n448);
    nor g366(n473 ,n289 ,n384);
    nor g367(n472 ,n272 ,n384);
    nor g368(n471 ,n275 ,n384);
    nor g369(n470 ,n271 ,n384);
    nor g370(n469 ,n305 ,n384);
    nor g371(n468 ,n287 ,n384);
    nor g372(n467 ,n297 ,n384);
    nor g373(n466 ,n288 ,n384);
    nor g374(n465 ,n293 ,n384);
    nor g375(n464 ,n302 ,n384);
    nor g376(n463 ,n266 ,n384);
    nor g377(n462 ,n279 ,n384);
    nor g378(n461 ,n301 ,n384);
    nor g379(n460 ,n283 ,n384);
    nor g380(n459 ,n277 ,n384);
    nor g381(n458 ,n280 ,n384);
    nor g382(n457 ,n273 ,n384);
    nor g383(n456 ,n285 ,n384);
    nor g384(n455 ,n284 ,n384);
    nor g385(n454 ,n303 ,n384);
    nor g386(n453 ,n300 ,n384);
    nor g387(n452 ,n270 ,n384);
    nor g388(n451 ,n299 ,n384);
    nor g389(n450 ,n268 ,n384);
    nor g390(n485 ,n318 ,n408);
    nor g391(n484 ,n306 ,n394);
    nor g392(n483 ,n314 ,n406);
    nor g393(n482 ,n316 ,n404);
    nor g394(n481 ,n311 ,n396);
    nor g395(n480 ,n310 ,n390);
    nor g396(n479 ,n317 ,n388);
    nor g397(n478 ,n309 ,n392);
    nor g398(n477 ,n315 ,n386);
    nor g399(n476 ,n312 ,n412);
    nor g400(n475 ,n307 ,n410);
    nor g401(n474 ,n319 ,n402);
    not g402(n449 ,n448);
    xnor g403(n434 ,n376 ,n13[0]);
    nor g404(n433 ,n304 ,n384);
    nor g405(n432 ,n276 ,n384);
    nor g406(n431 ,n274 ,n384);
    nor g407(n430 ,n278 ,n384);
    nor g408(n429 ,n295 ,n384);
    nor g409(n428 ,n290 ,n384);
    nor g410(n427 ,n282 ,n384);
    nor g411(n426 ,n269 ,n384);
    nor g412(n425 ,n267 ,n384);
    nor g413(n424 ,n281 ,n384);
    nor g414(n423 ,n291 ,n384);
    nor g415(n422 ,n292 ,n384);
    nor g416(n421 ,n298 ,n384);
    or g417(n420 ,n365 ,n383);
    or g418(n419 ,n362 ,n384);
    nor g419(n418 ,n9[1] ,n400);
    nor g420(n417 ,n286 ,n384);
    nor g421(n416 ,n10[1] ,n400);
    nor g422(n415 ,n381 ,n398);
    nor g423(n414 ,n8[1] ,n400);
    nor g424(n413 ,n382 ,n399);
    nor g425(n448 ,n361 ,n380);
    nor g426(n447 ,n374 ,n407);
    nor g427(n446 ,n374 ,n389);
    nor g428(n445 ,n374 ,n409);
    nor g429(n444 ,n374 ,n385);
    nor g430(n443 ,n374 ,n403);
    nor g431(n442 ,n374 ,n395);
    nor g432(n441 ,n374 ,n405);
    nor g433(n440 ,n374 ,n401);
    nor g434(n439 ,n374 ,n393);
    nor g435(n438 ,n374 ,n411);
    nor g436(n437 ,n374 ,n397);
    nor g437(n436 ,n374 ,n387);
    nor g438(n435 ,n374 ,n391);
    not g439(n412 ,n411);
    not g440(n410 ,n409);
    not g441(n408 ,n407);
    not g442(n406 ,n405);
    not g443(n404 ,n403);
    not g444(n402 ,n401);
    nor g445(n399 ,n296 ,n375);
    nor g446(n398 ,n294 ,n375);
    nor g447(n397 ,n262 ,n379);
    nor g448(n411 ,n254 ,n379);
    nor g449(n409 ,n264 ,n379);
    nor g450(n407 ,n259 ,n379);
    nor g451(n405 ,n261 ,n379);
    nor g452(n403 ,n253 ,n379);
    nor g453(n401 ,n257 ,n379);
    nor g454(n400 ,n313 ,n379);
    not g455(n396 ,n395);
    not g456(n394 ,n393);
    not g457(n392 ,n391);
    not g458(n390 ,n389);
    not g459(n388 ,n387);
    not g460(n386 ,n385);
    or g461(n383 ,n7[12] ,n378);
    nor g462(n382 ,n320 ,n376);
    nor g463(n381 ,n321 ,n376);
    or g464(n380 ,n13[2] ,n375);
    nor g465(n395 ,n258 ,n379);
    nor g466(n393 ,n265 ,n379);
    nor g467(n391 ,n252 ,n379);
    nor g468(n389 ,n260 ,n379);
    nor g469(n387 ,n251 ,n379);
    nor g470(n385 ,n255 ,n379);
    or g471(n384 ,n14[2] ,n372);
    or g472(n378 ,n366 ,n359);
    or g473(n377 ,n358 ,n363);
    or g474(n379 ,n369 ,n370);
    not g475(n375 ,n376);
    nor g476(n373 ,n371 ,n368);
    or g477(n372 ,n14[1] ,n370);
    nor g478(n376 ,n14[1] ,n364);
    nor g479(n374 ,n1 ,n371);
    not g480(n369 ,n368);
    nor g481(n367 ,n251 ,n256);
    or g482(n366 ,n7[6] ,n7[7]);
    or g483(n365 ,n7[10] ,n7[11]);
    nor g484(n371 ,n308 ,n14[2]);
    or g485(n370 ,n308 ,n1);
    nor g486(n368 ,n322 ,n14[2]);
    or g487(n363 ,n7[4] ,n7[5]);
    nor g488(n362 ,n3[0] ,n707);
    or g489(n361 ,n13[0] ,n13[1]);
    or g490(n360 ,n7[0] ,n7[1]);
    or g491(n359 ,n7[8] ,n7[9]);
    or g492(n358 ,n7[2] ,n7[3]);
    or g493(n364 ,n14[0] ,n14[2]);
    not g494(n357 ,n8[7]);
    not g495(n356 ,n8[9]);
    not g496(n355 ,n9[9]);
    not g497(n354 ,n8[3]);
    not g498(n353 ,n10[11]);
    not g499(n352 ,n8[8]);
    not g500(n351 ,n8[2]);
    not g501(n350 ,n10[12]);
    not g502(n349 ,n10[4]);
    not g503(n348 ,n10[9]);
    not g504(n347 ,n9[0]);
    not g505(n346 ,n10[0]);
    not g506(n345 ,n8[4]);
    not g507(n344 ,n9[5]);
    not g508(n343 ,n9[2]);
    not g509(n342 ,n9[11]);
    not g510(n341 ,n9[3]);
    not g511(n340 ,n10[2]);
    not g512(n339 ,n8[0]);
    not g513(n338 ,n10[8]);
    not g514(n337 ,n8[5]);
    not g515(n336 ,n9[10]);
    not g516(n335 ,n9[4]);
    not g517(n334 ,n9[8]);
    not g518(n333 ,n8[10]);
    not g519(n332 ,n10[3]);
    not g520(n331 ,n8[12]);
    not g521(n330 ,n10[7]);
    not g522(n329 ,n9[7]);
    not g523(n328 ,n9[12]);
    not g524(n327 ,n10[6]);
    not g525(n326 ,n10[10]);
    not g526(n325 ,n8[6]);
    not g527(n324 ,n10[5]);
    not g528(n323 ,n9[6]);
    not g529(n322 ,n14[1]);
    not g530(n321 ,n13[2]);
    not g531(n320 ,n13[1]);
    not g532(n319 ,n7[2]);
    not g533(n318 ,n7[7]);
    not g534(n317 ,n7[0]);
    not g535(n316 ,n7[10]);
    not g536(n315 ,n7[4]);
    not g537(n314 ,n7[11]);
    not g538(n313 ,n7[1]);
    not g539(n312 ,n7[3]);
    not g540(n311 ,n7[9]);
    not g541(n310 ,n7[8]);
    not g542(n309 ,n7[6]);
    not g543(n308 ,n14[0]);
    not g544(n307 ,n7[5]);
    not g545(n306 ,n7[12]);
    not g546(n305 ,n714);
    not g547(n304 ,n778);
    not g548(n303 ,n755);
    not g549(n302 ,n772);
    not g550(n301 ,n749);
    not g551(n300 ,n770);
    not g552(n299 ,n716);
    not g553(n298 ,n776);
    not g554(n297 ,n752);
    not g555(n296 ,n795);
    not g556(n295 ,n780);
    not g557(n294 ,n794);
    not g558(n293 ,n712);
    not g559(n292 ,n748);
    not g560(n291 ,n747);
    not g561(n290 ,n12[1]);
    not g562(n289 ,n717);
    not g563(n288 ,n713);
    not g564(n287 ,n715);
    not g565(n286 ,n775);
    not g566(n285 ,n753);
    not g567(n284 ,n710);
    not g568(n283 ,n750);
    not g569(n282 ,n744);
    not g570(n281 ,n746);
    not g571(n280 ,n751);
    not g572(n279 ,n773);
    not g573(n278 ,n754);
    not g574(n277 ,n769);
    not g575(n276 ,n777);
    not g576(n275 ,n774);
    not g577(n274 ,n779);
    not g578(n273 ,n709);
    not g579(n272 ,n719);
    not g580(n271 ,n718);
    not g581(n270 ,n708);
    not g582(n269 ,n768);
    not g583(n268 ,n771);
    not g584(n267 ,n745);
    not g585(n266 ,n711);
    not g586(n265 ,n11[12]);
    not g587(n264 ,n11[5]);
    not g588(n263 ,n8[11]);
    not g589(n262 ,n11[1]);
    not g590(n261 ,n11[11]);
    not g591(n260 ,n11[8]);
    not g592(n259 ,n11[7]);
    not g593(n258 ,n11[9]);
    not g594(n257 ,n11[2]);
    not g595(n256 ,n707);
    not g596(n255 ,n11[4]);
    not g597(n254 ,n11[3]);
    not g598(n253 ,n11[10]);
    not g599(n252 ,n11[6]);
    not g600(n251 ,n3[0]);
    xnor g601(n780 ,n793 ,n81);
    nor g602(n81 ,n42 ,n80);
    xor g603(n779 ,n56 ,n79);
    nor g604(n80 ,n56 ,n79);
    nor g605(n79 ,n39 ,n78);
    xor g606(n778 ,n54 ,n77);
    nor g607(n78 ,n54 ,n77);
    nor g608(n77 ,n45 ,n76);
    xor g609(n777 ,n52 ,n75);
    nor g610(n76 ,n52 ,n75);
    nor g611(n75 ,n35 ,n74);
    xor g612(n776 ,n50 ,n73);
    nor g613(n74 ,n50 ,n73);
    nor g614(n73 ,n46 ,n72);
    xor g615(n775 ,n55 ,n71);
    nor g616(n72 ,n55 ,n71);
    nor g617(n71 ,n44 ,n70);
    xor g618(n774 ,n53 ,n69);
    nor g619(n70 ,n53 ,n69);
    nor g620(n69 ,n43 ,n68);
    xor g621(n773 ,n57 ,n67);
    nor g622(n68 ,n57 ,n67);
    nor g623(n67 ,n40 ,n66);
    xor g624(n772 ,n51 ,n65);
    nor g625(n66 ,n51 ,n65);
    nor g626(n65 ,n38 ,n64);
    xnor g627(n771 ,n58 ,n62);
    nor g628(n64 ,n58 ,n63);
    not g629(n63 ,n62);
    nor g630(n62 ,n37 ,n61);
    xnor g631(n770 ,n49 ,n60);
    nor g632(n61 ,n49 ,n60);
    nor g633(n60 ,n36 ,n59);
    xnor g634(n769 ,n48 ,n47);
    nor g635(n59 ,n47 ,n48);
    nor g636(n768 ,n47 ,n41);
    xnor g637(n58 ,n784 ,n12[3]);
    xnor g638(n57 ,n786 ,n12[5]);
    xnor g639(n56 ,n792 ,n12[11]);
    xnor g640(n55 ,n788 ,n12[7]);
    xnor g641(n54 ,n791 ,n12[10]);
    xnor g642(n53 ,n787 ,n12[6]);
    xnor g643(n52 ,n790 ,n12[9]);
    xnor g644(n51 ,n785 ,n12[4]);
    xnor g645(n50 ,n789 ,n12[8]);
    xnor g646(n49 ,n783 ,n12[2]);
    xnor g647(n48 ,n782 ,n12[1]);
    nor g648(n46 ,n16 ,n24);
    nor g649(n45 ,n32 ,n33);
    nor g650(n44 ,n29 ,n28);
    nor g651(n43 ,n30 ,n20);
    nor g652(n42 ,n27 ,n19);
    nor g653(n47 ,n17 ,n15);
    nor g654(n41 ,n781 ,n11[1]);
    nor g655(n40 ,n18 ,n25);
    nor g656(n39 ,n31 ,n34);
    nor g657(n38 ,n21 ,n22);
    nor g658(n37 ,n783 ,n12[2]);
    nor g659(n36 ,n782 ,n12[1]);
    nor g660(n35 ,n23 ,n26);
    not g661(n34 ,n12[10]);
    not g662(n33 ,n12[9]);
    not g663(n32 ,n790);
    not g664(n31 ,n791);
    not g665(n30 ,n786);
    not g666(n29 ,n787);
    not g667(n28 ,n12[6]);
    not g668(n27 ,n792);
    not g669(n26 ,n12[8]);
    not g670(n25 ,n12[4]);
    not g671(n24 ,n12[7]);
    not g672(n23 ,n789);
    not g673(n22 ,n12[3]);
    not g674(n21 ,n784);
    not g675(n20 ,n12[5]);
    not g676(n19 ,n12[11]);
    not g677(n18 ,n785);
    not g678(n17 ,n781);
    not g679(n16 ,n788);
    not g680(n15 ,n11[1]);
    xor g681(n755 ,n767 ,n129);
    nor g682(n129 ,n93 ,n128);
    xnor g683(n754 ,n105 ,n127);
    nor g684(n128 ,n105 ,n127);
    nor g685(n127 ,n87 ,n126);
    xor g686(n753 ,n107 ,n124);
    nor g687(n126 ,n107 ,n125);
    not g688(n125 ,n124);
    nor g689(n124 ,n94 ,n123);
    xnor g690(n752 ,n106 ,n121);
    nor g691(n123 ,n106 ,n122);
    not g692(n122 ,n121);
    nor g693(n121 ,n89 ,n120);
    xnor g694(n751 ,n98 ,n119);
    nor g695(n120 ,n98 ,n119);
    nor g696(n119 ,n91 ,n118);
    xnor g697(n750 ,n104 ,n117);
    nor g698(n118 ,n104 ,n117);
    nor g699(n117 ,n92 ,n116);
    xnor g700(n749 ,n101 ,n115);
    nor g701(n116 ,n101 ,n115);
    nor g702(n115 ,n90 ,n114);
    xnor g703(n748 ,n100 ,n113);
    nor g704(n114 ,n100 ,n113);
    nor g705(n113 ,n88 ,n112);
    xnor g706(n747 ,n99 ,n111);
    nor g707(n112 ,n99 ,n111);
    nor g708(n111 ,n86 ,n110);
    xnor g709(n746 ,n102 ,n109);
    nor g710(n110 ,n102 ,n109);
    nor g711(n109 ,n95 ,n108);
    xnor g712(n745 ,n103 ,n97);
    nor g713(n108 ,n97 ,n103);
    nor g714(n744 ,n97 ,n96);
    xnor g715(n107 ,n765 ,n12[11]);
    xnor g716(n106 ,n764 ,n12[10]);
    xnor g717(n105 ,n766 ,n11[11]);
    xnor g718(n104 ,n762 ,n12[8]);
    xnor g719(n103 ,n757 ,n12[3]);
    xnor g720(n102 ,n758 ,n12[4]);
    xnor g721(n101 ,n761 ,n12[7]);
    xnor g722(n100 ,n760 ,n12[6]);
    xnor g723(n99 ,n759 ,n12[5]);
    xnor g724(n98 ,n763 ,n12[9]);
    nor g725(n96 ,n756 ,n12[2]);
    nor g726(n95 ,n757 ,n12[3]);
    nor g727(n94 ,n83 ,n85);
    nor g728(n93 ,n766 ,n11[11]);
    nor g729(n92 ,n761 ,n12[7]);
    nor g730(n97 ,n82 ,n84);
    nor g731(n91 ,n762 ,n12[8]);
    nor g732(n90 ,n760 ,n12[6]);
    nor g733(n89 ,n763 ,n12[9]);
    nor g734(n88 ,n759 ,n12[5]);
    nor g735(n87 ,n765 ,n12[11]);
    nor g736(n86 ,n758 ,n12[4]);
    not g737(n85 ,n12[10]);
    not g738(n84 ,n12[2]);
    not g739(n83 ,n764);
    not g740(n82 ,n756);
    xnor g741(n743 ,n149 ,n184);
    nor g742(n184 ,n137 ,n183);
    xnor g743(n741 ,n155 ,n182);
    nor g744(n183 ,n155 ,n182);
    nor g745(n182 ,n143 ,n181);
    xnor g746(n739 ,n153 ,n180);
    nor g747(n181 ,n153 ,n180);
    nor g748(n180 ,n138 ,n179);
    xnor g749(n737 ,n152 ,n178);
    nor g750(n179 ,n152 ,n178);
    nor g751(n178 ,n140 ,n177);
    xor g752(n735 ,n158 ,n175);
    nor g753(n177 ,n158 ,n176);
    not g754(n176 ,n175);
    nor g755(n175 ,n147 ,n174);
    xor g756(n733 ,n159 ,n173);
    nor g757(n174 ,n159 ,n173);
    nor g758(n173 ,n145 ,n172);
    xnor g759(n731 ,n160 ,n170);
    nor g760(n172 ,n160 ,n171);
    not g761(n171 ,n170);
    nor g762(n170 ,n139 ,n169);
    xnor g763(n729 ,n154 ,n168);
    nor g764(n169 ,n154 ,n168);
    nor g765(n168 ,n141 ,n167);
    xnor g766(n727 ,n151 ,n166);
    nor g767(n167 ,n151 ,n166);
    nor g768(n166 ,n144 ,n165);
    xnor g769(n725 ,n157 ,n164);
    nor g770(n165 ,n157 ,n164);
    nor g771(n164 ,n136 ,n163);
    xnor g772(n723 ,n156 ,n162);
    nor g773(n163 ,n156 ,n162);
    nor g774(n162 ,n146 ,n161);
    xnor g775(n721 ,n150 ,n148);
    nor g776(n161 ,n148 ,n150);
    nor g777(n707 ,n148 ,n142);
    xnor g778(n160 ,n2[6] ,n3[6]);
    xnor g779(n159 ,n2[7] ,n3[7]);
    xnor g780(n158 ,n2[8] ,n3[8]);
    xnor g781(n157 ,n2[3] ,n3[3]);
    xnor g782(n156 ,n2[2] ,n3[2]);
    xnor g783(n149 ,n2[12] ,n3[12]);
    xnor g784(n155 ,n2[11] ,n3[11]);
    xnor g785(n154 ,n2[5] ,n3[5]);
    xnor g786(n153 ,n2[10] ,n3[10]);
    xnor g787(n152 ,n2[9] ,n3[9]);
    xnor g788(n151 ,n2[4] ,n3[4]);
    xnor g789(n150 ,n2[1] ,n3[1]);
    nor g790(n147 ,n134 ,n135);
    nor g791(n146 ,n2[1] ,n3[1]);
    nor g792(n145 ,n132 ,n131);
    nor g793(n144 ,n2[3] ,n3[3]);
    nor g794(n143 ,n2[10] ,n3[10]);
    nor g795(n148 ,n133 ,n130);
    nor g796(n142 ,n2[0] ,n3[0]);
    nor g797(n141 ,n2[4] ,n3[4]);
    nor g798(n140 ,n2[8] ,n3[8]);
    nor g799(n139 ,n2[5] ,n3[5]);
    nor g800(n138 ,n2[9] ,n3[9]);
    nor g801(n137 ,n2[11] ,n3[11]);
    nor g802(n136 ,n2[2] ,n3[2]);
    not g803(n135 ,n3[7]);
    not g804(n134 ,n2[7]);
    not g805(n133 ,n2[0]);
    not g806(n132 ,n2[6]);
    not g807(n131 ,n3[6]);
    not g808(n130 ,n3[0]);
    xor g809(n719 ,n215 ,n246);
    nor g810(n246 ,n210 ,n245);
    xor g811(n718 ,n221 ,n244);
    nor g812(n245 ,n221 ,n244);
    nor g813(n244 ,n213 ,n243);
    xor g814(n717 ,n223 ,n242);
    nor g815(n243 ,n223 ,n242);
    nor g816(n242 ,n209 ,n241);
    xor g817(n716 ,n220 ,n240);
    nor g818(n241 ,n220 ,n240);
    nor g819(n240 ,n206 ,n239);
    xor g820(n715 ,n222 ,n238);
    nor g821(n239 ,n222 ,n238);
    nor g822(n238 ,n212 ,n237);
    xor g823(n714 ,n225 ,n236);
    nor g824(n237 ,n225 ,n236);
    nor g825(n236 ,n203 ,n235);
    xor g826(n713 ,n224 ,n234);
    nor g827(n235 ,n224 ,n234);
    nor g828(n234 ,n211 ,n233);
    xor g829(n712 ,n219 ,n232);
    nor g830(n233 ,n219 ,n232);
    nor g831(n232 ,n207 ,n231);
    xnor g832(n711 ,n218 ,n229);
    nor g833(n231 ,n218 ,n230);
    not g834(n230 ,n229);
    nor g835(n229 ,n205 ,n228);
    xnor g836(n710 ,n217 ,n227);
    nor g837(n228 ,n217 ,n227);
    nor g838(n227 ,n204 ,n226);
    xnor g839(n709 ,n216 ,n214);
    nor g840(n226 ,n214 ,n216);
    nor g841(n708 ,n214 ,n208);
    xnor g842(n225 ,n732 ,n12[6]);
    xnor g843(n224 ,n730 ,n12[5]);
    xnor g844(n223 ,n738 ,n12[9]);
    xnor g845(n222 ,n734 ,n12[7]);
    xnor g846(n221 ,n740 ,n12[10]);
    xnor g847(n220 ,n736 ,n12[8]);
    xnor g848(n219 ,n728 ,n12[4]);
    xnor g849(n218 ,n726 ,n12[3]);
    xnor g850(n217 ,n724 ,n12[2]);
    xnor g851(n216 ,n722 ,n12[1]);
    xnor g852(n215 ,n12[11] ,n742);
    nor g853(n213 ,n201 ,n186);
    nor g854(n212 ,n198 ,n194);
    nor g855(n211 ,n187 ,n188);
    nor g856(n210 ,n199 ,n185);
    nor g857(n209 ,n200 ,n202);
    nor g858(n214 ,n191 ,n189);
    nor g859(n208 ,n720 ,n11[1]);
    nor g860(n207 ,n190 ,n197);
    nor g861(n206 ,n195 ,n193);
    nor g862(n205 ,n724 ,n12[2]);
    nor g863(n204 ,n722 ,n12[1]);
    nor g864(n203 ,n192 ,n196);
    not g865(n202 ,n12[8]);
    not g866(n201 ,n738);
    not g867(n200 ,n736);
    not g868(n199 ,n740);
    not g869(n198 ,n732);
    not g870(n197 ,n12[3]);
    not g871(n196 ,n12[5]);
    not g872(n195 ,n734);
    not g873(n194 ,n12[6]);
    not g874(n193 ,n12[7]);
    not g875(n192 ,n730);
    not g876(n191 ,n720);
    not g877(n190 ,n726);
    not g878(n189 ,n11[1]);
    not g879(n188 ,n12[4]);
    not g880(n187 ,n728);
    not g881(n186 ,n12[9]);
    not g882(n185 ,n12[10]);
    xor g883(n794 ,n13[2] ,n250);
    nor g884(n795 ,n250 ,n249);
    nor g885(n250 ,n248 ,n247);
    nor g886(n249 ,n13[1] ,n13[0]);
    not g887(n248 ,n13[1]);
    not g888(n247 ,n13[0]);
    not g889(n847 ,n1);
    nor g890(n848 ,n847 ,n846);
    or g891(n846 ,n843 ,n845);
    nor g892(n845 ,n844 ,n842);
    or g893(n844 ,n840 ,n841);
    nor g894(n843 ,n2[13] ,n2[12]);
    nor g895(n842 ,n2[11] ,n2[10]);
    not g896(n841 ,n2[12]);
    not g897(n840 ,n2[13]);
    xor g898(n11[12] ,n3[12] ,n839);
    nor g899(n11[11] ,n838 ,n839);
    nor g900(n839 ,n805 ,n837);
    nor g901(n838 ,n3[11] ,n836);
    nor g902(n11[10] ,n835 ,n836);
    not g903(n837 ,n836);
    nor g904(n836 ,n798 ,n834);
    nor g905(n835 ,n3[10] ,n833);
    nor g906(n11[9] ,n832 ,n833);
    not g907(n834 ,n833);
    nor g908(n833 ,n799 ,n831);
    nor g909(n832 ,n3[9] ,n830);
    nor g910(n11[8] ,n829 ,n830);
    not g911(n831 ,n830);
    nor g912(n830 ,n803 ,n828);
    nor g913(n829 ,n3[8] ,n827);
    nor g914(n11[7] ,n826 ,n827);
    not g915(n828 ,n827);
    nor g916(n827 ,n797 ,n825);
    nor g917(n826 ,n3[7] ,n824);
    nor g918(n11[6] ,n823 ,n824);
    not g919(n825 ,n824);
    nor g920(n824 ,n802 ,n822);
    nor g921(n823 ,n3[6] ,n821);
    nor g922(n11[5] ,n820 ,n821);
    not g923(n822 ,n821);
    nor g924(n821 ,n800 ,n819);
    nor g925(n820 ,n3[5] ,n818);
    nor g926(n11[4] ,n817 ,n818);
    not g927(n819 ,n818);
    nor g928(n818 ,n801 ,n816);
    nor g929(n817 ,n3[4] ,n815);
    nor g930(n11[3] ,n814 ,n815);
    not g931(n816 ,n815);
    nor g932(n815 ,n806 ,n813);
    nor g933(n814 ,n3[3] ,n812);
    nor g934(n11[2] ,n811 ,n812);
    not g935(n813 ,n812);
    nor g936(n812 ,n807 ,n810);
    nor g937(n811 ,n3[2] ,n809);
    nor g938(n11[1] ,n809 ,n808);
    not g939(n810 ,n809);
    nor g940(n809 ,n796 ,n804);
    nor g941(n808 ,n3[1] ,n848);
    not g942(n807 ,n3[2]);
    not g943(n806 ,n3[3]);
    not g944(n805 ,n3[11]);
    not g945(n804 ,n848);
    not g946(n803 ,n3[8]);
    not g947(n802 ,n3[6]);
    not g948(n801 ,n3[4]);
    not g949(n800 ,n3[5]);
    not g950(n799 ,n3[9]);
    not g951(n798 ,n3[10]);
    not g952(n797 ,n3[7]);
    not g953(n796 ,n3[1]);
endmodule
