module top(n0, n1, n2, n3, n4, n5, n6, n7, n8);
    input n0, n1, n2;
    input [11:0] n3, n4;
    input [2:0] n5;
    output n6, n7;
    output [11:0] n8;
    wire n0, n1, n2;
    wire [11:0] n3, n4;
    wire [2:0] n5;
    wire n6, n7;
    wire [11:0] n8;
    wire [11:0] n9;
    wire [11:0] n10;
    wire [2:0] n11;
    wire [11:0] n12;
    wire [18:0] n13;
    wire [19:0] n14;
    wire [12:0] n15;
    wire [12:0] n16;
    wire [12:0] n17;
    wire [12:0] n18;
    wire [3:0] n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
    wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
    wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627;
    wire n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635;
    wire n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643;
    wire n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
    wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
    wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
    wire n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675;
    wire n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683;
    wire n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
    wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
    wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707;
    wire n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715;
    wire n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723;
    wire n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
    wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
    wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
    wire n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755;
    wire n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763;
    wire n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
    wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
    wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787;
    wire n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795;
    wire n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803;
    wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
    wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
    wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
    wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
    wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
    wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
    wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
    wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
    wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
    wire n1876, n1877, n1878;
    not g0(n1693 ,n1877);
    or g1(n1704 ,n1692 ,n1670);
    or g2(n1703 ,n1683 ,n1662);
    or g3(n1698 ,n1689 ,n1665);
    or g4(n1724 ,n1690 ,n1669);
    or g5(n1723 ,n1688 ,n1666);
    or g6(n1722 ,n1687 ,n1663);
    or g7(n1701 ,n1685 ,n1659);
    or g8(n1697 ,n1686 ,n1661);
    or g9(n1721 ,n1684 ,n1668);
    or g10(n1696 ,n1681 ,n1664);
    or g11(n1720 ,n1682 ,n1660);
    or g12(n1719 ,n1680 ,n1658);
    or g13(n1702 ,n1691 ,n1667);
    or g14(n1700 ,n1677 ,n1654);
    or g15(n1695 ,n1678 ,n1656);
    or g16(n1718 ,n1679 ,n1657);
    or g17(n1717 ,n1676 ,n1655);
    or g18(n1699 ,n1653 ,n1672);
    or g19(n1726 ,n1675 ,n1673);
    or g20(n1725 ,n1674 ,n1671);
    nor g21(n1692 ,n1611 ,n1610);
    nor g22(n1691 ,n1638 ,n1610);
    nor g23(n1690 ,n1637 ,n1609);
    nor g24(n1689 ,n1634 ,n1610);
    nor g25(n1688 ,n1620 ,n1609);
    nor g26(n1687 ,n1642 ,n1609);
    nor g27(n1705 ,n1643 ,n1610);
    nor g28(n1686 ,n1648 ,n1610);
    nor g29(n1685 ,n1636 ,n1610);
    nor g30(n1684 ,n1623 ,n1609);
    nor g31(n1683 ,n1628 ,n1610);
    nor g32(n1682 ,n1630 ,n1609);
    nor g33(n1681 ,n1622 ,n1610);
    nor g34(n1680 ,n1615 ,n1609);
    nor g35(n1679 ,n1650 ,n1609);
    nor g36(n1678 ,n1649 ,n1610);
    nor g37(n1677 ,n1612 ,n1610);
    nor g38(n1676 ,n1621 ,n1609);
    nor g39(n1727 ,n1618 ,n1609);
    nor g40(n1675 ,n1627 ,n1609);
    nor g41(n1674 ,n1625 ,n1609);
    nor g42(n1673 ,n1616 ,n9[11]);
    nor g43(n1672 ,n1619 ,n10[11]);
    nor g44(n1671 ,n1624 ,n9[11]);
    nor g45(n1670 ,n1633 ,n10[11]);
    nor g46(n1669 ,n1632 ,n9[11]);
    nor g47(n1668 ,n1644 ,n9[11]);
    nor g48(n1667 ,n1641 ,n10[11]);
    nor g49(n1666 ,n1647 ,n9[11]);
    nor g50(n1665 ,n1629 ,n10[11]);
    nor g51(n1664 ,n1640 ,n10[11]);
    nor g52(n1663 ,n1646 ,n9[11]);
    nor g53(n1662 ,n1635 ,n10[11]);
    nor g54(n1661 ,n1652 ,n10[11]);
    nor g55(n1660 ,n1626 ,n9[11]);
    nor g56(n1659 ,n1613 ,n10[11]);
    nor g57(n1658 ,n1614 ,n9[11]);
    nor g58(n1657 ,n1639 ,n9[11]);
    nor g59(n1656 ,n1631 ,n10[11]);
    nor g60(n1655 ,n1651 ,n9[11]);
    nor g61(n1654 ,n1617 ,n10[11]);
    nor g62(n1653 ,n1645 ,n1610);
    not g63(n1652 ,n10[3]);
    not g64(n1651 ,n9[1]);
    not g65(n1783 ,n1);
    not g66(n1650 ,n1729);
    not g67(n1649 ,n1706);
    not g68(n1648 ,n1708);
    not g69(n1647 ,n9[7]);
    not g70(n1646 ,n9[6]);
    not g71(n1645 ,n1710);
    not g72(n1644 ,n9[5]);
    not g73(n1643 ,n1716);
    not g74(n1642 ,n1733);
    not g75(n1641 ,n10[8]);
    not g76(n1640 ,n10[2]);
    not g77(n1639 ,n9[2]);
    not g78(n1638 ,n1713);
    not g79(n1637 ,n1735);
    not g80(n1636 ,n1712);
    not g81(n1635 ,n10[9]);
    not g82(n1634 ,n1709);
    not g83(n1633 ,n10[10]);
    not g84(n1632 ,n9[8]);
    not g85(n1631 ,n10[1]);
    not g86(n1630 ,n1731);
    not g87(n1629 ,n10[4]);
    not g88(n1628 ,n1714);
    not g89(n1627 ,n1737);
    not g90(n1626 ,n9[4]);
    not g91(n1625 ,n1736);
    not g92(n1624 ,n9[9]);
    not g93(n1623 ,n1732);
    not g94(n1622 ,n1707);
    not g95(n1621 ,n1728);
    not g96(n1620 ,n1734);
    not g97(n1619 ,n10[5]);
    not g98(n1618 ,n1738);
    not g99(n1617 ,n10[6]);
    not g100(n1616 ,n9[10]);
    not g101(n1615 ,n1730);
    not g102(n1614 ,n9[3]);
    not g103(n1613 ,n10[7]);
    not g104(n1612 ,n1711);
    not g105(n1611 ,n1715);
    not g106(n1610 ,n10[11]);
    not g107(n1609 ,n9[11]);
    dff g108(.RN(n1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n8[0]));
    dff g109(.RN(n1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n8[1]));
    dff g110(.RN(n1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n8[2]));
    dff g111(.RN(n1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n8[3]));
    dff g112(.RN(n1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n8[4]));
    dff g113(.RN(n1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n8[5]));
    dff g114(.RN(n1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n8[6]));
    dff g115(.RN(n1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n8[7]));
    dff g116(.RN(n1), .SN(1'b1), .CK(n0), .D(n1606), .Q(n8[8]));
    dff g117(.RN(n1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n8[9]));
    dff g118(.RN(n1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n8[10]));
    dff g119(.RN(n1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n8[11]));
    dff g120(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[0]), .Q(n9[0]));
    dff g121(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[1]), .Q(n9[1]));
    dff g122(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[2]), .Q(n9[2]));
    dff g123(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[3]), .Q(n9[3]));
    dff g124(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[4]), .Q(n9[4]));
    dff g125(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[5]), .Q(n9[5]));
    dff g126(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[6]), .Q(n9[6]));
    dff g127(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[7]), .Q(n9[7]));
    dff g128(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[8]), .Q(n9[8]));
    dff g129(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[9]), .Q(n9[9]));
    dff g130(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[10]), .Q(n9[10]));
    dff g131(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[11]), .Q(n9[11]));
    dff g132(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[0]), .Q(n10[0]));
    dff g133(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[1]), .Q(n10[1]));
    dff g134(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[2]), .Q(n10[2]));
    dff g135(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[3]), .Q(n10[3]));
    dff g136(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[4]), .Q(n10[4]));
    dff g137(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[5]), .Q(n10[5]));
    dff g138(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[6]), .Q(n10[6]));
    dff g139(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[7]), .Q(n10[7]));
    dff g140(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[8]), .Q(n10[8]));
    dff g141(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[9]), .Q(n10[9]));
    dff g142(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[10]), .Q(n10[10]));
    dff g143(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[11]), .Q(n1608));
    dff g144(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[0]), .Q(n11[0]));
    dff g145(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[1]), .Q(n11[1]));
    dff g146(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[2]), .Q(n11[2]));
    dff g147(.RN(n1), .SN(1'b1), .CK(n0), .D(n1518), .Q(n12[0]));
    dff g148(.RN(n1), .SN(1'b1), .CK(n0), .D(n1517), .Q(n12[1]));
    dff g149(.RN(n1), .SN(1'b1), .CK(n0), .D(n1516), .Q(n12[2]));
    dff g150(.RN(n1), .SN(1'b1), .CK(n0), .D(n1515), .Q(n12[3]));
    dff g151(.RN(n1), .SN(1'b1), .CK(n0), .D(n1514), .Q(n12[4]));
    dff g152(.RN(n1), .SN(1'b1), .CK(n0), .D(n1512), .Q(n12[5]));
    dff g153(.RN(n1), .SN(1'b1), .CK(n0), .D(n1531), .Q(n12[6]));
    dff g154(.RN(n1), .SN(1'b1), .CK(n0), .D(n1535), .Q(n12[7]));
    dff g155(.RN(n1), .SN(1'b1), .CK(n0), .D(n1534), .Q(n12[8]));
    dff g156(.RN(n1), .SN(1'b1), .CK(n0), .D(n1533), .Q(n12[9]));
    dff g157(.RN(n1), .SN(1'b1), .CK(n0), .D(n1532), .Q(n12[10]));
    dff g158(.RN(n1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n12[11]));
    dff g159(.RN(n1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n1095));
    dff g160(.RN(n1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n7));
    dff g161(.RN(n1), .SN(1'b1), .CK(n0), .D(n2), .Q(n1878));
    dff g162(.RN(n1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n6));
    or g163(n1607 ,n1529 ,n1600);
    or g164(n1606 ,n1498 ,n1593);
    or g165(n1605 ,n1509 ,n1587);
    or g166(n1604 ,n1507 ,n1591);
    or g167(n1603 ,n1505 ,n1590);
    or g168(n1602 ,n1503 ,n1589);
    or g169(n1601 ,n1501 ,n1588);
    or g170(n1600 ,n1567 ,n1586);
    or g171(n1599 ,n1492 ,n1584);
    or g172(n1598 ,n1494 ,n1585);
    or g173(n1597 ,n1499 ,n1592);
    or g174(n1596 ,n1488 ,n1582);
    or g175(n1595 ,n1299 ,n1581);
    or g176(n1594 ,n1496 ,n1580);
    or g177(n1593 ,n1462 ,n1579);
    or g178(n1592 ,n1463 ,n1576);
    or g179(n1591 ,n1468 ,n1578);
    or g180(n1590 ,n1466 ,n1577);
    or g181(n1589 ,n1465 ,n1575);
    or g182(n1588 ,n1464 ,n1574);
    or g183(n1587 ,n1471 ,n1573);
    nor g184(n1586 ,n1319 ,n1572);
    or g185(n1585 ,n1460 ,n1571);
    or g186(n1584 ,n1459 ,n1570);
    or g187(n1583 ,n1342 ,n1569);
    or g188(n1582 ,n1458 ,n1568);
    nor g189(n1581 ,n1373 ,n1572);
    or g190(n1580 ,n1461 ,n1566);
    or g191(n1579 ,n1560 ,n1541);
    or g192(n1578 ,n1564 ,n1546);
    or g193(n1577 ,n1563 ,n1545);
    or g194(n1576 ,n1543 ,n1557);
    or g195(n1575 ,n1562 ,n1544);
    or g196(n1574 ,n1561 ,n1542);
    or g197(n1573 ,n1565 ,n1549);
    or g198(n1571 ,n1558 ,n1539);
    or g199(n1570 ,n1555 ,n1537);
    or g200(n1569 ,n1538 ,n1556);
    or g201(n1568 ,n1554 ,n1536);
    nor g202(n1567 ,n1320 ,n1552);
    or g203(n1566 ,n1559 ,n1540);
    nor g204(n1572 ,n1095 ,n1553);
    or g205(n1565 ,n1456 ,n1530);
    or g206(n1564 ,n1453 ,n1528);
    or g207(n1563 ,n1450 ,n1527);
    or g208(n1562 ,n1447 ,n1526);
    or g209(n1561 ,n1444 ,n1525);
    or g210(n1560 ,n1440 ,n1524);
    or g211(n1559 ,n1437 ,n1523);
    or g212(n1558 ,n1432 ,n1522);
    or g213(n1557 ,n1521 ,n1433);
    or g214(n1556 ,n1426 ,n1519);
    or g215(n1555 ,n1425 ,n1520);
    or g216(n1554 ,n1429 ,n1513);
    nor g217(n1553 ,n1551 ,n1550);
    or g218(n1552 ,n1548 ,n1547);
    nor g219(n1551 ,n1303 ,n1473);
    nor g220(n1550 ,n1266 ,n1472);
    or g221(n1549 ,n1455 ,n1454);
    nor g222(n1548 ,n1306 ,n1467);
    nor g223(n1547 ,n1265 ,n1510);
    or g224(n1546 ,n1452 ,n1451);
    or g225(n1545 ,n1449 ,n1448);
    or g226(n1544 ,n1446 ,n1445);
    or g227(n1543 ,n1441 ,n1436);
    or g228(n1542 ,n1443 ,n1442);
    or g229(n1541 ,n1439 ,n1438);
    or g230(n1540 ,n1435 ,n1434);
    or g231(n1539 ,n1431 ,n1430);
    or g232(n1538 ,n1428 ,n1427);
    or g233(n1537 ,n1423 ,n1424);
    or g234(n1536 ,n1422 ,n1457);
    or g235(n1535 ,n1292 ,n1486);
    or g236(n1534 ,n1312 ,n1485);
    or g237(n1533 ,n1315 ,n1484);
    or g238(n1532 ,n1295 ,n1483);
    or g239(n1531 ,n1277 ,n1475);
    or g240(n1530 ,n1407 ,n1508);
    or g241(n1529 ,n1470 ,n1469);
    or g242(n1528 ,n1406 ,n1506);
    or g243(n1527 ,n1405 ,n1504);
    or g244(n1526 ,n1404 ,n1502);
    or g245(n1525 ,n1403 ,n1500);
    or g246(n1524 ,n1401 ,n1497);
    or g247(n1523 ,n1400 ,n1495);
    or g248(n1522 ,n1399 ,n1493);
    or g249(n1521 ,n1374 ,n1474);
    or g250(n1520 ,n1420 ,n1489);
    or g251(n1519 ,n1491 ,n1490);
    or g252(n1518 ,n1278 ,n1481);
    or g253(n1517 ,n1275 ,n1480);
    or g254(n1516 ,n1281 ,n1479);
    or g255(n1515 ,n1274 ,n1478);
    or g256(n1514 ,n1296 ,n1477);
    or g257(n1513 ,n1396 ,n1487);
    or g258(n1512 ,n1313 ,n1476);
    or g259(n1511 ,n1304 ,n1482);
    or g260(n1510 ,n13[15] ,n1340);
    nor g261(n1509 ,n1252 ,n1375);
    nor g262(n1508 ,n1192 ,n1421);
    nor g263(n1507 ,n1181 ,n1375);
    nor g264(n1506 ,n1182 ,n1421);
    nor g265(n1505 ,n1177 ,n1375);
    nor g266(n1504 ,n1167 ,n1421);
    nor g267(n1503 ,n1186 ,n1375);
    nor g268(n1502 ,n1255 ,n1421);
    nor g269(n1501 ,n1258 ,n1375);
    nor g270(n1500 ,n1199 ,n1421);
    nor g271(n1499 ,n1210 ,n1375);
    nor g272(n1498 ,n1173 ,n1375);
    nor g273(n1497 ,n1253 ,n1421);
    nor g274(n1496 ,n1257 ,n1375);
    nor g275(n1495 ,n1189 ,n1421);
    nor g276(n1494 ,n1176 ,n1375);
    nor g277(n1493 ,n1196 ,n1421);
    nor g278(n1492 ,n1185 ,n1375);
    nor g279(n1491 ,n1254 ,n1421);
    nor g280(n1490 ,n1195 ,n1375);
    nor g281(n1489 ,n1174 ,n1421);
    nor g282(n1488 ,n1191 ,n1375);
    nor g283(n1487 ,n1194 ,n1421);
    nor g284(n1486 ,n1159 ,n1373);
    nor g285(n1485 ,n1154 ,n1373);
    nor g286(n1484 ,n1156 ,n1373);
    nor g287(n1483 ,n1164 ,n1373);
    nor g288(n1482 ,n1137 ,n1373);
    nor g289(n1481 ,n1162 ,n1373);
    nor g290(n1480 ,n1151 ,n1373);
    nor g291(n1479 ,n1230 ,n1373);
    nor g292(n1478 ,n1144 ,n1373);
    nor g293(n1477 ,n1147 ,n1373);
    nor g294(n1476 ,n1152 ,n1373);
    nor g295(n1475 ,n1238 ,n1373);
    nor g296(n1474 ,n1136 ,n1421);
    or g297(n1473 ,n1307 ,n1397);
    nor g298(n1471 ,n1309 ,n1338);
    nor g299(n1470 ,n1310 ,n1343);
    nor g300(n1469 ,n1308 ,n1353);
    nor g301(n1468 ,n1282 ,n1337);
    or g302(n1467 ,n1149 ,n1419);
    nor g303(n1466 ,n1298 ,n1336);
    nor g304(n1465 ,n1294 ,n1335);
    nor g305(n1464 ,n1291 ,n1334);
    nor g306(n1463 ,n1271 ,n1333);
    nor g307(n1462 ,n1288 ,n1332);
    nor g308(n1461 ,n1289 ,n1331);
    nor g309(n1460 ,n1284 ,n1330);
    nor g310(n1459 ,n1280 ,n1329);
    nor g311(n1458 ,n1300 ,n1339);
    or g312(n1457 ,n1371 ,n1417);
    or g313(n1456 ,n1362 ,n1395);
    or g314(n1455 ,n1369 ,n1374);
    or g315(n1454 ,n1394 ,n1411);
    or g316(n1453 ,n1367 ,n1393);
    or g317(n1452 ,n1366 ,n1374);
    or g318(n1451 ,n1392 ,n1416);
    or g319(n1450 ,n1364 ,n1391);
    or g320(n1449 ,n1363 ,n1374);
    or g321(n1448 ,n1390 ,n1415);
    or g322(n1447 ,n1361 ,n1389);
    or g323(n1446 ,n1360 ,n1374);
    or g324(n1445 ,n1388 ,n1414);
    or g325(n1444 ,n1359 ,n1387);
    or g326(n1443 ,n1358 ,n1374);
    or g327(n1442 ,n1386 ,n1413);
    or g328(n1441 ,n1357 ,n1402);
    or g329(n1440 ,n1347 ,n1385);
    or g330(n1439 ,n1356 ,n1374);
    or g331(n1438 ,n1384 ,n1412);
    or g332(n1437 ,n1354 ,n1382);
    or g333(n1436 ,n1381 ,n1355);
    or g334(n1435 ,n1365 ,n1374);
    or g335(n1434 ,n1380 ,n1409);
    or g336(n1433 ,n1379 ,n1344);
    or g337(n1432 ,n1368 ,n1378);
    or g338(n1431 ,n1352 ,n1374);
    or g339(n1430 ,n1377 ,n1410);
    or g340(n1429 ,n1345 ,n1370);
    or g341(n1428 ,n1376 ,n1351);
    or g342(n1427 ,n1383 ,n1374);
    or g343(n1426 ,n1372 ,n1398);
    or g344(n1425 ,n1350 ,n1418);
    or g345(n1424 ,n1349 ,n1408);
    or g346(n1423 ,n1348 ,n1374);
    or g347(n1422 ,n1346 ,n1374);
    nor g348(n1420 ,n1155 ,n1327);
    nor g349(n1418 ,n1184 ,n1320);
    nor g350(n1417 ,n1208 ,n1322);
    nor g351(n1416 ,n1213 ,n1322);
    nor g352(n1415 ,n1207 ,n1322);
    nor g353(n1414 ,n1215 ,n1322);
    nor g354(n1413 ,n1211 ,n1322);
    nor g355(n1412 ,n1206 ,n1322);
    nor g356(n1411 ,n1205 ,n1322);
    nor g357(n1410 ,n1209 ,n1322);
    nor g358(n1409 ,n1214 ,n1322);
    nor g359(n1408 ,n1212 ,n1322);
    nor g360(n1407 ,n1158 ,n1327);
    nor g361(n1406 ,n1236 ,n1327);
    nor g362(n1405 ,n1235 ,n1327);
    nor g363(n1404 ,n1227 ,n1327);
    nor g364(n1403 ,n1143 ,n1327);
    nor g365(n1402 ,n1160 ,n1327);
    nor g366(n1401 ,n1145 ,n1327);
    nor g367(n1400 ,n1231 ,n1327);
    nor g368(n1399 ,n1138 ,n1327);
    nor g369(n1398 ,n1140 ,n1327);
    or g370(n1397 ,n1157 ,n1323);
    nor g371(n1396 ,n1247 ,n1327);
    nor g372(n1395 ,n1180 ,n1320);
    nor g373(n1394 ,n1168 ,n1321);
    nor g374(n1393 ,n1169 ,n1320);
    nor g375(n1392 ,n1188 ,n1321);
    nor g376(n1391 ,n1198 ,n1320);
    nor g377(n1390 ,n1200 ,n1321);
    nor g378(n1389 ,n1166 ,n1320);
    nor g379(n1388 ,n1172 ,n1321);
    nor g380(n1387 ,n1251 ,n1320);
    nor g381(n1386 ,n1259 ,n1321);
    nor g382(n1385 ,n1175 ,n1320);
    nor g383(n1384 ,n1250 ,n1321);
    nor g384(n1383 ,n1141 ,n1321);
    nor g385(n1382 ,n1183 ,n1320);
    nor g386(n1381 ,n1171 ,n1320);
    nor g387(n1380 ,n1190 ,n1321);
    nor g388(n1379 ,n1170 ,n1321);
    nor g389(n1378 ,n1193 ,n1320);
    nor g390(n1377 ,n1178 ,n1321);
    nor g391(n1376 ,n1139 ,n1320);
    or g392(n1421 ,n1228 ,n1328);
    nor g393(n1372 ,n1137 ,n1319);
    nor g394(n1371 ,n1197 ,n1321);
    nor g395(n1370 ,n1179 ,n1320);
    nor g396(n1369 ,n1247 ,n1318);
    nor g397(n1368 ,n1164 ,n1319);
    nor g398(n1367 ,n1147 ,n1319);
    nor g399(n1366 ,n1158 ,n1318);
    nor g400(n1365 ,n1145 ,n1318);
    nor g401(n1364 ,n1152 ,n1319);
    nor g402(n1363 ,n1236 ,n1318);
    nor g403(n1362 ,n1144 ,n1319);
    nor g404(n1361 ,n1238 ,n1319);
    nor g405(n1360 ,n1235 ,n1318);
    nor g406(n1359 ,n1159 ,n1319);
    nor g407(n1358 ,n1227 ,n1318);
    nor g408(n1357 ,n1162 ,n1319);
    nor g409(n1356 ,n1143 ,n1318);
    nor g410(n1355 ,n1187 ,n1318);
    nor g411(n1354 ,n1156 ,n1319);
    or g412(n1353 ,n1262 ,n1318);
    nor g413(n1352 ,n1231 ,n1318);
    nor g414(n1351 ,n1138 ,n1318);
    nor g415(n1350 ,n1151 ,n1319);
    nor g416(n1349 ,n1256 ,n1321);
    nor g417(n1348 ,n1160 ,n1318);
    nor g418(n1347 ,n1154 ,n1319);
    nor g419(n1346 ,n1155 ,n1318);
    nor g420(n1345 ,n1230 ,n1319);
    nor g421(n1344 ,n1136 ,n1322);
    or g422(n1343 ,n1267 ,n1321);
    nor g423(n1342 ,n1326 ,n1317);
    or g424(n1341 ,n14[11] ,n1324);
    or g425(n1339 ,n1276 ,n1326);
    or g426(n1338 ,n1314 ,n1326);
    or g427(n1337 ,n1305 ,n1326);
    or g428(n1336 ,n1297 ,n1326);
    or g429(n1335 ,n1293 ,n1326);
    or g430(n1334 ,n1286 ,n1326);
    or g431(n1333 ,n1290 ,n1326);
    or g432(n1332 ,n1287 ,n1326);
    or g433(n1331 ,n1285 ,n1326);
    or g434(n1330 ,n1283 ,n1326);
    or g435(n1329 ,n1279 ,n1326);
    or g436(n1375 ,n1694 ,n1328);
    nor g437(n1374 ,n1693 ,n1318);
    or g438(n1373 ,n1201 ,n1319);
    or g439(n1325 ,n1264 ,n1261);
    or g440(n1324 ,n1263 ,n1260);
    or g441(n1328 ,n1203 ,n1273);
    or g442(n1327 ,n1202 ,n1134);
    or g443(n1326 ,n1202 ,n1135);
    xor g444(n1317 ,n9[11] ,n1608);
    or g445(n1316 ,n1302 ,n1311);
    or g446(n1322 ,n1268 ,n1269);
    or g447(n1321 ,n11[2] ,n1270);
    or g448(n1320 ,n11[2] ,n1134);
    or g449(n1319 ,n11[2] ,n1272);
    or g450(n1318 ,n11[2] ,n1135);
    nor g451(n1315 ,n1237 ,n1878);
    nor g452(n1314 ,n1220 ,n9[3]);
    nor g453(n1313 ,n1249 ,n1878);
    nor g454(n1312 ,n1242 ,n1878);
    or g455(n1311 ,n1150 ,n1139);
    nor g456(n1310 ,n1142 ,n1141);
    nor g457(n1309 ,n1205 ,n10[3]);
    nor g458(n1308 ,n1140 ,n1138);
    or g459(n1307 ,n1163 ,n1153);
    or g460(n1306 ,n1241 ,n1226);
    nor g461(n1305 ,n1224 ,n9[4]);
    nor g462(n1304 ,n1229 ,n1878);
    or g463(n1303 ,n1146 ,n1137);
    or g464(n1302 ,n1165 ,n1239);
    or g465(n1301 ,n1161 ,n1148);
    nor g466(n1300 ,n1208 ,n10[2]);
    nor g467(n1299 ,n1245 ,n1878);
    nor g468(n1298 ,n1207 ,n10[5]);
    nor g469(n1297 ,n1225 ,n9[5]);
    nor g470(n1296 ,n1246 ,n1878);
    nor g471(n1295 ,n1234 ,n1878);
    nor g472(n1294 ,n1215 ,n10[6]);
    nor g473(n1293 ,n1222 ,n9[6]);
    nor g474(n1292 ,n1248 ,n1878);
    nor g475(n1291 ,n1211 ,n10[7]);
    nor g476(n1290 ,n1210 ,n9[0]);
    nor g477(n1289 ,n1214 ,n10[9]);
    nor g478(n1288 ,n1206 ,n10[8]);
    nor g479(n1287 ,n1219 ,n9[8]);
    nor g480(n1286 ,n1223 ,n9[7]);
    nor g481(n1285 ,n1216 ,n9[9]);
    nor g482(n1284 ,n1209 ,n10[10]);
    nor g483(n1283 ,n1218 ,n9[10]);
    nor g484(n1282 ,n1213 ,n10[4]);
    nor g485(n1281 ,n1232 ,n1878);
    nor g486(n1280 ,n1212 ,n10[1]);
    nor g487(n1279 ,n1221 ,n9[1]);
    nor g488(n1278 ,n1243 ,n1878);
    nor g489(n1277 ,n1244 ,n1878);
    nor g490(n1276 ,n1217 ,n9[2]);
    nor g491(n1275 ,n1233 ,n1878);
    nor g492(n1274 ,n1240 ,n1878);
    or g493(n1273 ,n1204 ,n1202);
    or g494(n1272 ,n1204 ,n1203);
    nor g495(n1271 ,n1136 ,n10[0]);
    or g496(n1270 ,n1204 ,n11[1]);
    or g497(n1269 ,n1202 ,n11[1]);
    or g498(n1268 ,n1204 ,n9[11]);
    nor g499(n1267 ,n15[12] ,n16[11]);
    or g500(n1266 ,n14[17] ,n14[16]);
    or g501(n1265 ,n13[17] ,n13[16]);
    or g502(n1264 ,n13[14] ,n13[13]);
    or g503(n1263 ,n14[15] ,n14[14]);
    nor g504(n1262 ,n17[12] ,n18[11]);
    or g505(n1261 ,n13[12] ,n13[11]);
    or g506(n1260 ,n14[13] ,n14[12]);
    not g507(n1259 ,n1757);
    not g508(n1258 ,n1701);
    not g509(n1257 ,n1703);
    not g510(n1256 ,n1751);
    not g511(n1255 ,n1722);
    not g512(n1254 ,n1727);
    not g513(n1253 ,n1724);
    not g514(n1252 ,n1697);
    not g515(n1251 ,n1779);
    not g516(n1250 ,n1758);
    not g517(n1249 ,n12[5]);
    not g518(n1248 ,n12[7]);
    not g519(n1247 ,n1764);
    not g520(n1246 ,n12[4]);
    not g521(n1245 ,n1095);
    not g522(n1244 ,n12[6]);
    not g523(n1243 ,n12[0]);
    not g524(n1242 ,n12[8]);
    not g525(n1241 ,n13[17]);
    not g526(n1240 ,n12[3]);
    not g527(n1239 ,n13[13]);
    not g528(n1238 ,n1745);
    not g529(n1237 ,n12[9]);
    not g530(n1236 ,n1766);
    not g531(n1235 ,n1767);
    not g532(n1234 ,n12[10]);
    not g533(n1233 ,n12[1]);
    not g534(n1232 ,n12[2]);
    not g535(n1231 ,n1771);
    not g536(n1230 ,n1741);
    not g537(n1229 ,n12[11]);
    not g538(n1228 ,n1694);
    not g539(n1227 ,n1768);
    not g540(n1226 ,n13[16]);
    not g541(n1225 ,n10[5]);
    not g542(n1224 ,n10[4]);
    not g543(n1223 ,n10[7]);
    buf g544(n10[11] ,n1608);
    not g545(n1222 ,n10[6]);
    not g546(n1221 ,n10[1]);
    not g547(n1220 ,n10[3]);
    not g548(n1219 ,n10[8]);
    not g549(n1218 ,n10[10]);
    not g550(n1217 ,n10[2]);
    not g551(n1216 ,n10[9]);
    not g552(n1215 ,n9[6]);
    not g553(n1214 ,n9[9]);
    not g554(n1213 ,n9[4]);
    not g555(n1212 ,n9[1]);
    not g556(n1211 ,n9[7]);
    not g557(n1210 ,n10[0]);
    not g558(n1209 ,n9[10]);
    not g559(n1208 ,n9[2]);
    not g560(n1207 ,n9[5]);
    not g561(n1206 ,n9[8]);
    not g562(n1205 ,n9[3]);
    not g563(n1136 ,n9[0]);
    not g564(n1204 ,n11[0]);
    not g565(n1203 ,n11[1]);
    not g566(n1202 ,n11[2]);
    not g567(n1201 ,n1878);
    not g568(n1200 ,n1755);
    not g569(n1199 ,n1723);
    not g570(n1198 ,n1777);
    not g571(n1197 ,n1752);
    not g572(n1196 ,n1726);
    not g573(n1195 ,n1705);
    not g574(n1194 ,n1718);
    not g575(n1193 ,n1782);
    not g576(n1192 ,n1719);
    not g577(n1191 ,n1696);
    not g578(n1190 ,n1759);
    not g579(n1189 ,n1725);
    not g580(n1188 ,n1754);
    not g581(n1187 ,n1761);
    not g582(n1186 ,n1700);
    not g583(n1185 ,n1695);
    not g584(n1184 ,n1773);
    not g585(n1183 ,n1781);
    not g586(n1182 ,n1720);
    not g587(n1181 ,n1698);
    not g588(n1180 ,n1775);
    not g589(n1179 ,n1774);
    not g590(n1178 ,n1760);
    not g591(n1177 ,n1699);
    not g592(n1176 ,n1704);
    not g593(n1175 ,n1780);
    not g594(n1174 ,n1717);
    not g595(n1173 ,n1702);
    not g596(n1172 ,n1756);
    not g597(n1171 ,n1772);
    not g598(n1170 ,n1750);
    not g599(n1169 ,n1776);
    not g600(n1168 ,n1753);
    not g601(n1167 ,n1721);
    not g602(n1166 ,n1778);
    not g603(n1165 ,n13[14]);
    not g604(n1164 ,n1749);
    not g605(n1163 ,n14[14]);
    not g606(n1162 ,n1739);
    not g607(n1161 ,n14[17]);
    not g608(n1160 ,n1762);
    not g609(n1159 ,n1746);
    not g610(n1158 ,n1765);
    not g611(n1157 ,n14[15]);
    not g612(n1156 ,n1748);
    not g613(n1155 ,n1763);
    not g614(n1154 ,n1747);
    not g615(n1153 ,n14[13]);
    not g616(n1152 ,n1744);
    not g617(n1151 ,n1740);
    not g618(n1150 ,n13[12]);
    not g619(n1149 ,n13[15]);
    not g620(n1148 ,n14[16]);
    not g621(n1147 ,n1743);
    not g622(n1146 ,n14[12]);
    not g623(n1145 ,n1770);
    not g624(n1144 ,n1742);
    not g625(n1143 ,n1769);
    not g626(n1142 ,n15[12]);
    not g627(n1141 ,n16[11]);
    not g628(n1140 ,n17[12]);
    not g629(n1139 ,n13[11]);
    not g630(n1138 ,n18[11]);
    not g631(n1137 ,n14[11]);
    or g632(n1135 ,n11[0] ,n11[1]);
    or g633(n1134 ,n1203 ,n11[0]);
    xnor g634(n13[17] ,n516 ,n881);
    nor g635(n881 ,n605 ,n880);
    xnor g636(n13[16] ,n626 ,n879);
    nor g637(n880 ,n609 ,n879);
    nor g638(n879 ,n704 ,n878);
    xnor g639(n13[15] ,n714 ,n877);
    nor g640(n878 ,n706 ,n877);
    nor g641(n877 ,n760 ,n876);
    xnor g642(n13[14] ,n772 ,n875);
    nor g643(n876 ,n767 ,n875);
    nor g644(n875 ,n786 ,n874);
    xnor g645(n13[13] ,n800 ,n873);
    nor g646(n874 ,n787 ,n873);
    nor g647(n873 ,n807 ,n872);
    xnor g648(n13[12] ,n813 ,n871);
    nor g649(n872 ,n806 ,n871);
    nor g650(n871 ,n823 ,n870);
    xnor g651(n13[11] ,n832 ,n869);
    nor g652(n870 ,n824 ,n869);
    nor g653(n869 ,n834 ,n868);
    xnor g654(n1782 ,n847 ,n867);
    nor g655(n868 ,n836 ,n867);
    nor g656(n867 ,n849 ,n866);
    xnor g657(n1781 ,n851 ,n865);
    nor g658(n866 ,n865 ,n850);
    nor g659(n865 ,n864 ,n835);
    xnor g660(n1780 ,n845 ,n863);
    nor g661(n864 ,n841 ,n863);
    nor g662(n863 ,n842 ,n862);
    xnor g663(n1779 ,n844 ,n861);
    nor g664(n862 ,n843 ,n861);
    nor g665(n861 ,n840 ,n860);
    xnor g666(n1778 ,n846 ,n859);
    nor g667(n860 ,n839 ,n859);
    nor g668(n859 ,n801 ,n858);
    xor g669(n1777 ,n814 ,n857);
    nor g670(n858 ,n804 ,n857);
    nor g671(n857 ,n791 ,n856);
    xnor g672(n1776 ,n798 ,n855);
    nor g673(n856 ,n790 ,n855);
    nor g674(n855 ,n774 ,n854);
    xor g675(n1775 ,n797 ,n853);
    nor g676(n854 ,n788 ,n853);
    nor g677(n853 ,n763 ,n852);
    xnor g678(n1774 ,n773 ,n848);
    nor g679(n852 ,n762 ,n848);
    xnor g680(n851 ,n837 ,n825);
    nor g681(n850 ,n826 ,n837);
    nor g682(n849 ,n825 ,n838);
    nor g683(n848 ,n728 ,n833);
    xnor g684(n847 ,n815 ,n829);
    xnor g685(n846 ,n817 ,n779);
    xnor g686(n845 ,n821 ,n827);
    xnor g687(n844 ,n819 ,n809);
    xnor g688(n1773 ,n740 ,n831);
    nor g689(n843 ,n810 ,n819);
    nor g690(n842 ,n809 ,n820);
    nor g691(n841 ,n828 ,n821);
    nor g692(n840 ,n779 ,n818);
    nor g693(n839 ,n780 ,n817);
    not g694(n838 ,n837);
    nor g695(n836 ,n830 ,n815);
    nor g696(n835 ,n827 ,n822);
    nor g697(n834 ,n829 ,n816);
    nor g698(n833 ,n729 ,n831);
    xnor g699(n832 ,n777 ,n811);
    xnor g700(n837 ,n799 ,n725);
    not g701(n830 ,n829);
    not g702(n828 ,n827);
    not g703(n826 ,n825);
    nor g704(n824 ,n812 ,n777);
    nor g705(n823 ,n811 ,n778);
    nor g706(n831 ,n687 ,n802);
    nor g707(n829 ,n785 ,n803);
    nor g708(n827 ,n793 ,n805);
    nor g709(n825 ,n784 ,n808);
    not g710(n822 ,n821);
    not g711(n820 ,n819);
    not g712(n818 ,n817);
    not g713(n816 ,n815);
    xnor g714(n1772 ,n713 ,n783);
    xnor g715(n814 ,n781 ,n754);
    xnor g716(n813 ,n744 ,n795);
    xnor g717(n821 ,n771 ,n742);
    xnor g718(n819 ,n770 ,n756);
    xnor g719(n817 ,n769 ,n735);
    xnor g720(n815 ,n768 ,n736);
    not g721(n812 ,n811);
    not g722(n810 ,n809);
    nor g723(n808 ,n738 ,n789);
    nor g724(n807 ,n745 ,n795);
    nor g725(n806 ,n744 ,n796);
    nor g726(n805 ,n737 ,n792);
    nor g727(n804 ,n755 ,n782);
    nor g728(n811 ,n761 ,n776);
    nor g729(n809 ,n766 ,n775);
    nor g730(n803 ,n725 ,n794);
    nor g731(n802 ,n709 ,n783);
    nor g732(n801 ,n754 ,n781);
    xnor g733(n800 ,n746 ,n731);
    xnor g734(n799 ,n752 ,n641);
    xnor g735(n798 ,n750 ,n733);
    xnor g736(n797 ,n748 ,n715);
    not g737(n796 ,n795);
    nor g738(n794 ,n642 ,n752);
    nor g739(n793 ,n649 ,n757);
    nor g740(n792 ,n650 ,n756);
    nor g741(n791 ,n733 ,n751);
    nor g742(n790 ,n734 ,n750);
    nor g743(n789 ,n648 ,n742);
    nor g744(n788 ,n716 ,n749);
    nor g745(n787 ,n732 ,n746);
    nor g746(n786 ,n731 ,n747);
    nor g747(n785 ,n641 ,n753);
    nor g748(n784 ,n647 ,n743);
    nor g749(n795 ,n707 ,n758);
    not g750(n782 ,n781);
    not g751(n780 ,n779);
    not g752(n778 ,n777);
    nor g753(n776 ,n736 ,n764);
    nor g754(n775 ,n735 ,n765);
    nor g755(n774 ,n715 ,n748);
    xnor g756(n773 ,n717 ,n691);
    xnor g757(n772 ,n639 ,n723);
    xnor g758(n771 ,n738 ,n647);
    xnor g759(n770 ,n737 ,n649);
    xnor g760(n769 ,n599 ,n719);
    xnor g761(n768 ,n721 ,n566);
    nor g762(n783 ,n663 ,n759);
    xnor g763(n781 ,n712 ,n726);
    nor g764(n779 ,n686 ,n741);
    xnor g765(n777 ,n711 ,n739);
    nor g766(n767 ,n639 ,n724);
    nor g767(n766 ,n600 ,n719);
    nor g768(n765 ,n599 ,n720);
    nor g769(n764 ,n567 ,n721);
    nor g770(n763 ,n691 ,n718);
    nor g771(n762 ,n692 ,n717);
    nor g772(n761 ,n566 ,n722);
    nor g773(n760 ,n640 ,n723);
    nor g774(n759 ,n661 ,n730);
    nor g775(n758 ,n739 ,n705);
    not g776(n757 ,n756);
    not g777(n755 ,n754);
    not g778(n753 ,n752);
    not g779(n751 ,n750);
    not g780(n749 ,n748);
    not g781(n747 ,n746);
    not g782(n745 ,n744);
    not g783(n743 ,n742);
    nor g784(n741 ,n697 ,n726);
    xnor g785(n740 ,n693 ,n645);
    xnor g786(n756 ,n682 ,n621);
    nor g787(n754 ,n634 ,n727);
    xnor g788(n752 ,n680 ,n619);
    xnor g789(n750 ,n681 ,n695);
    xnor g790(n748 ,n679 ,n583);
    xnor g791(n746 ,n685 ,n571);
    xnor g792(n744 ,n683 ,n655);
    xnor g793(n742 ,n684 ,n656);
    not g794(n734 ,n733);
    not g795(n732 ,n731);
    nor g796(n730 ,n633 ,n708);
    nor g797(n729 ,n646 ,n693);
    nor g798(n728 ,n645 ,n694);
    nor g799(n727 ,n675 ,n696);
    nor g800(n739 ,n678 ,n700);
    nor g801(n738 ,n672 ,n701);
    nor g802(n737 ,n636 ,n699);
    nor g803(n736 ,n669 ,n710);
    nor g804(n735 ,n676 ,n698);
    nor g805(n733 ,n674 ,n689);
    nor g806(n731 ,n662 ,n688);
    not g807(n724 ,n723);
    not g808(n722 ,n721);
    not g809(n720 ,n719);
    not g810(n718 ,n717);
    not g811(n716 ,n715);
    xnor g812(n714 ,n617 ,n643);
    xnor g813(n713 ,n616 ,n637);
    xnor g814(n712 ,n593 ,n653);
    xnor g815(n711 ,n613 ,n651);
    xnor g816(n726 ,n630 ,n597);
    nor g817(n725 ,n631 ,n703);
    nor g818(n723 ,n664 ,n702);
    xnor g819(n721 ,n628 ,n587);
    xnor g820(n719 ,n629 ,n577);
    xnor g821(n717 ,n627 ,n581);
    nor g822(n715 ,n668 ,n690);
    nor g823(n710 ,n551 ,n660);
    nor g824(n709 ,n616 ,n638);
    nor g825(n708 ,n520 ,n658);
    nor g826(n707 ,n614 ,n651);
    nor g827(n706 ,n644 ,n617);
    nor g828(n705 ,n613 ,n652);
    nor g829(n704 ,n643 ,n618);
    nor g830(n703 ,n673 ,n657);
    nor g831(n702 ,n571 ,n659);
    nor g832(n701 ,n621 ,n671);
    nor g833(n700 ,n570 ,n670);
    nor g834(n699 ,n569 ,n677);
    nor g835(n698 ,n553 ,n635);
    nor g836(n697 ,n594 ,n654);
    not g837(n696 ,n695);
    not g838(n694 ,n693);
    not g839(n692 ,n691);
    nor g840(n690 ,n554 ,n667);
    nor g841(n689 ,n556 ,n632);
    nor g842(n688 ,n655 ,n666);
    nor g843(n687 ,n615 ,n637);
    nor g844(n686 ,n593 ,n653);
    xnor g845(n685 ,n373 ,n575);
    xnor g846(n684 ,n481 ,n579);
    xnor g847(n683 ,n612 ,n545);
    xnor g848(n682 ,n539 ,n591);
    xnor g849(n681 ,n589 ,n549);
    xnor g850(n680 ,n595 ,n551);
    xnor g851(n679 ,n585 ,n556);
    xnor g852(n695 ,n573 ,n558);
    xnor g853(n693 ,n574 ,n601);
    nor g854(n691 ,n544 ,n665);
    nor g855(n678 ,n305 ,n587);
    nor g856(n677 ,n565 ,n578);
    nor g857(n676 ,n483 ,n598);
    nor g858(n675 ,n550 ,n590);
    nor g859(n674 ,n586 ,n584);
    nor g860(n673 ,n480 ,n580);
    nor g861(n672 ,n540 ,n591);
    nor g862(n671 ,n539 ,n592);
    nor g863(n670 ,n306 ,n588);
    nor g864(n669 ,n619 ,n596);
    nor g865(n668 ,n510 ,n581);
    nor g866(n667 ,n509 ,n582);
    nor g867(n666 ,n546 ,n612);
    nor g868(n665 ,n559 ,n602);
    nor g869(n664 ,n373 ,n576);
    nor g870(n663 ,n485 ,n624);
    nor g871(n662 ,n545 ,n611);
    nor g872(n661 ,n484 ,n625);
    nor g873(n660 ,n620 ,n595);
    nor g874(n659 ,n372 ,n575);
    nor g875(n658 ,n422 ,n623);
    not g876(n657 ,n656);
    not g877(n654 ,n653);
    not g878(n652 ,n651);
    not g879(n650 ,n649);
    not g880(n648 ,n647);
    not g881(n646 ,n645);
    not g882(n644 ,n643);
    not g883(n642 ,n641);
    not g884(n640 ,n639);
    not g885(n638 ,n637);
    nor g886(n636 ,n564 ,n577);
    nor g887(n635 ,n482 ,n597);
    nor g888(n634 ,n549 ,n589);
    nor g889(n633 ,n421 ,n622);
    nor g890(n632 ,n585 ,n583);
    nor g891(n631 ,n481 ,n579);
    xor g892(n630 ,n483 ,n553);
    xor g893(n629 ,n565 ,n569);
    xnor g894(n628 ,n306 ,n570);
    xnor g895(n627 ,n509 ,n554);
    xnor g896(n626 ,n371 ,n547);
    xnor g897(n656 ,n507 ,n557);
    nor g898(n655 ,n429 ,n604);
    nor g899(n653 ,n563 ,n606);
    xnor g900(n651 ,n515 ,n555);
    xnor g901(n649 ,n543 ,n572);
    nor g902(n647 ,n525 ,n603);
    nor g903(n645 ,n435 ,n608);
    nor g904(n643 ,n441 ,n607);
    nor g905(n641 ,n439 ,n610);
    xnor g906(n639 ,n506 ,n568);
    xnor g907(n637 ,n501 ,n552);
    not g908(n625 ,n624);
    not g909(n623 ,n622);
    not g910(n620 ,n619);
    not g911(n618 ,n617);
    not g912(n616 ,n615);
    not g913(n614 ,n613);
    not g914(n612 ,n611);
    nor g915(n610 ,n448 ,n557);
    nor g916(n609 ,n371 ,n548);
    nor g917(n608 ,n469 ,n552);
    nor g918(n607 ,n462 ,n568);
    nor g919(n606 ,n558 ,n560);
    nor g920(n605 ,n370 ,n547);
    nor g921(n604 ,n467 ,n555);
    nor g922(n603 ,n517 ,n572);
    xnor g923(n624 ,n495 ,n356);
    nor g924(n622 ,n465 ,n561);
    nor g925(n621 ,n436 ,n562);
    xnor g926(n619 ,n369 ,n508);
    xnor g927(n617 ,n367 ,n488);
    xnor g928(n615 ,n212 ,n498);
    xnor g929(n613 ,n505 ,n350);
    xnor g930(n611 ,n372 ,n491);
    not g931(n602 ,n601);
    not g932(n600 ,n599);
    not g933(n598 ,n597);
    not g934(n596 ,n595);
    not g935(n594 ,n593);
    not g936(n592 ,n591);
    not g937(n590 ,n589);
    not g938(n588 ,n587);
    not g939(n586 ,n585);
    not g940(n584 ,n583);
    not g941(n582 ,n581);
    not g942(n580 ,n579);
    not g943(n578 ,n577);
    not g944(n576 ,n575);
    xnor g945(n574 ,n541 ,n317);
    xnor g946(n573 ,n511 ,n325);
    xnor g947(n601 ,n492 ,n355);
    xnor g948(n599 ,n497 ,n513);
    xnor g949(n597 ,n496 ,n412);
    xnor g950(n595 ,n494 ,n413);
    xnor g951(n593 ,n493 ,n416);
    xnor g952(n591 ,n502 ,n415);
    xnor g953(n589 ,n490 ,n414);
    xnor g954(n587 ,n487 ,n352);
    xnor g955(n585 ,n489 ,n353);
    xnor g956(n583 ,n504 ,n453);
    xnor g957(n581 ,n486 ,n357);
    xnor g958(n579 ,n499 ,n351);
    xnor g959(n577 ,n500 ,n358);
    xnor g960(n575 ,n503 ,n360);
    not g961(n567 ,n566);
    not g962(n565 ,n564);
    nor g963(n563 ,n325 ,n512);
    nor g964(n562 ,n478 ,n514);
    nor g965(n561 ,n537 ,n463);
    nor g966(n560 ,n326 ,n511);
    nor g967(n559 ,n318 ,n542);
    nor g968(n572 ,n449 ,n534);
    nor g969(n571 ,n450 ,n535);
    nor g970(n570 ,n464 ,n532);
    nor g971(n569 ,n434 ,n531);
    nor g972(n568 ,n460 ,n523);
    nor g973(n566 ,n433 ,n530);
    nor g974(n564 ,n461 ,n533);
    not g975(n550 ,n549);
    not g976(n548 ,n547);
    not g977(n546 ,n545);
    nor g978(n544 ,n317 ,n541);
    xnor g979(n543 ,n451 ,n311);
    nor g980(n558 ,n455 ,n526);
    nor g981(n557 ,n428 ,n538);
    nor g982(n556 ,n427 ,n524);
    nor g983(n555 ,n426 ,n521);
    nor g984(n554 ,n446 ,n522);
    nor g985(n553 ,n432 ,n529);
    nor g986(n552 ,n443 ,n518);
    nor g987(n551 ,n431 ,n527);
    nor g988(n549 ,n430 ,n536);
    nor g989(n547 ,n444 ,n519);
    nor g990(n545 ,n457 ,n528);
    not g991(n542 ,n541);
    not g992(n540 ,n539);
    nor g993(n538 ,n415 ,n472);
    or g994(n537 ,n38 ,n442);
    nor g995(n536 ,n454 ,n473);
    nor g996(n535 ,n372 ,n477);
    nor g997(n534 ,n358 ,n466);
    nor g998(n533 ,n412 ,n459);
    nor g999(n532 ,n413 ,n458);
    nor g1000(n531 ,n416 ,n476);
    nor g1001(n530 ,n417 ,n468);
    nor g1002(n529 ,n414 ,n475);
    nor g1003(n528 ,n350 ,n437);
    nor g1004(n527 ,n351 ,n474);
    nor g1005(n526 ,n456 ,n353);
    nor g1006(n525 ,n312 ,n452);
    nor g1007(n524 ,n357 ,n471);
    nor g1008(n523 ,n360 ,n447);
    nor g1009(n522 ,n445 ,n355);
    nor g1010(n521 ,n352 ,n470);
    xor g1011(n520 ,n423 ,n302);
    nor g1012(n519 ,n420 ,n440);
    nor g1013(n518 ,n356 ,n479);
    nor g1014(n517 ,n311 ,n451);
    xnor g1015(n516 ,n371 ,n339);
    xnor g1016(n515 ,n306 ,n346);
    or g1017(n539 ,n438 ,n481);
    not g1018(n514 ,n513);
    not g1019(n512 ,n511);
    not g1020(n510 ,n509);
    xnor g1021(n508 ,n417 ,n396);
    xnor g1022(n507 ,n369 ,n307);
    xnor g1023(n506 ,n367 ,n404);
    xnor g1024(n505 ,n376 ,n384);
    xnor g1025(n504 ,n321 ,n323);
    xnor g1026(n503 ,n378 ,n402);
    xnor g1027(n502 ,n342 ,n344);
    xnor g1028(n501 ,n309 ,n406);
    xnor g1029(n500 ,n348 ,n410);
    xnor g1030(n499 ,n315 ,n333);
    xnor g1031(n498 ,n419 ,n295);
    xnor g1032(n497 ,n394 ,n382);
    xnor g1033(n496 ,n215 ,n408);
    xnor g1034(n495 ,n212 ,n319);
    xnor g1035(n494 ,n374 ,n392);
    xnor g1036(n493 ,n400 ,n331);
    xnor g1037(n492 ,n213 ,n327);
    xnor g1038(n491 ,n398 ,n380);
    xnor g1039(n490 ,n388 ,n386);
    xnor g1040(n489 ,n217 ,n313);
    xnor g1041(n488 ,n390 ,n420);
    xnor g1042(n487 ,n340 ,n329);
    xnor g1043(n486 ,n335 ,n337);
    xnor g1044(n513 ,n354 ,n298);
    xnor g1045(n511 ,n418 ,n296);
    xnor g1046(n509 ,n359 ,n300);
    not g1047(n485 ,n484);
    not g1048(n483 ,n482);
    not g1049(n480 ,n481);
    nor g1050(n479 ,n211 ,n320);
    nor g1051(n478 ,n383 ,n395);
    nor g1052(n477 ,n381 ,n399);
    nor g1053(n476 ,n332 ,n401);
    nor g1054(n475 ,n387 ,n389);
    nor g1055(n474 ,n334 ,n316);
    nor g1056(n473 ,n324 ,n322);
    nor g1057(n472 ,n345 ,n343);
    nor g1058(n471 ,n338 ,n336);
    nor g1059(n470 ,n330 ,n341);
    nor g1060(n469 ,n407 ,n310);
    nor g1061(n468 ,n397 ,n368);
    nor g1062(n467 ,n347 ,n305);
    nor g1063(n466 ,n411 ,n349);
    nor g1064(n465 ,n220 ,n424);
    nor g1065(n464 ,n392 ,n375);
    nor g1066(n462 ,n367 ,n405);
    nor g1067(n461 ,n216 ,n408);
    nor g1068(n460 ,n402 ,n379);
    nor g1069(n459 ,n215 ,n409);
    nor g1070(n458 ,n374 ,n393);
    nor g1071(n457 ,n384 ,n377);
    nor g1072(n456 ,n217 ,n314);
    nor g1073(n455 ,n218 ,n313);
    nor g1074(n484 ,n303 ,n423);
    nor g1075(n482 ,n297 ,n418);
    nor g1076(n481 ,n362 ,n364);
    not g1077(n454 ,n453);
    not g1078(n452 ,n451);
    nor g1079(n450 ,n380 ,n398);
    nor g1080(n449 ,n410 ,n348);
    nor g1081(n448 ,n369 ,n308);
    nor g1082(n447 ,n378 ,n403);
    nor g1083(n446 ,n214 ,n327);
    nor g1084(n445 ,n213 ,n328);
    nor g1085(n444 ,n367 ,n391);
    nor g1086(n443 ,n212 ,n319);
    or g1087(n442 ,n21 ,n365);
    nor g1088(n441 ,n404 ,n366);
    nor g1089(n440 ,n390 ,n366);
    nor g1090(n439 ,n307 ,n368);
    nor g1091(n438 ,n361 ,n363);
    nor g1092(n437 ,n376 ,n385);
    nor g1093(n436 ,n382 ,n394);
    nor g1094(n435 ,n406 ,n309);
    nor g1095(n434 ,n331 ,n400);
    nor g1096(n433 ,n396 ,n369);
    nor g1097(n432 ,n386 ,n388);
    nor g1098(n431 ,n333 ,n315);
    nor g1099(n430 ,n323 ,n321);
    nor g1100(n429 ,n346 ,n306);
    nor g1101(n428 ,n344 ,n342);
    nor g1102(n427 ,n337 ,n335);
    nor g1103(n426 ,n329 ,n340);
    nor g1104(n425 ,n304 ,n419);
    nor g1105(n453 ,n301 ,n359);
    nor g1106(n451 ,n299 ,n354);
    not g1107(n422 ,n421);
    not g1108(n411 ,n410);
    not g1109(n409 ,n408);
    not g1110(n407 ,n406);
    not g1111(n405 ,n404);
    not g1112(n403 ,n402);
    not g1113(n401 ,n400);
    not g1114(n399 ,n398);
    not g1115(n397 ,n396);
    not g1116(n395 ,n394);
    not g1117(n393 ,n392);
    not g1118(n391 ,n390);
    not g1119(n389 ,n388);
    not g1120(n387 ,n386);
    not g1121(n385 ,n384);
    not g1122(n383 ,n382);
    not g1123(n381 ,n380);
    not g1124(n379 ,n378);
    not g1125(n377 ,n376);
    not g1126(n375 ,n374);
    not g1127(n372 ,n373);
    not g1128(n370 ,n371);
    not g1129(n368 ,n369);
    not g1130(n366 ,n367);
    nor g1131(n365 ,n196 ,n229);
    nor g1132(n424 ,n194 ,n289);
    nor g1133(n423 ,n201 ,n291);
    nor g1134(n421 ,n150 ,n290);
    nor g1135(n420 ,n142 ,n227);
    nor g1136(n419 ,n198 ,n230);
    nor g1137(n418 ,n163 ,n264);
    nor g1138(n417 ,n165 ,n265);
    nor g1139(n416 ,n171 ,n271);
    nor g1140(n415 ,n139 ,n240);
    nor g1141(n414 ,n197 ,n259);
    nor g1142(n413 ,n190 ,n275);
    nor g1143(n412 ,n189 ,n276);
    nor g1144(n410 ,n169 ,n292);
    nor g1145(n408 ,n188 ,n277);
    nor g1146(n406 ,n186 ,n248);
    nor g1147(n404 ,n175 ,n284);
    nor g1148(n402 ,n203 ,n270);
    nor g1149(n400 ,n160 ,n273);
    nor g1150(n398 ,n176 ,n294);
    nor g1151(n396 ,n170 ,n269);
    nor g1152(n394 ,n185 ,n281);
    nor g1153(n392 ,n182 ,n283);
    nor g1154(n390 ,n175 ,n238);
    nor g1155(n388 ,n161 ,n260);
    nor g1156(n386 ,n162 ,n278);
    nor g1157(n384 ,n183 ,n244);
    nor g1158(n382 ,n145 ,n224);
    nor g1159(n380 ,n141 ,n282);
    nor g1160(n378 ,n176 ,n254);
    nor g1161(n376 ,n173 ,n263);
    nor g1162(n374 ,n174 ,n279);
    nor g1163(n373 ,n159 ,n293);
    nor g1164(n371 ,n221 ,n262);
    nor g1165(n369 ,n167 ,n267);
    nor g1166(n367 ,n192 ,n280);
    not g1167(n364 ,n363);
    not g1168(n362 ,n361);
    not g1169(n349 ,n348);
    not g1170(n347 ,n346);
    not g1171(n345 ,n344);
    not g1172(n343 ,n342);
    not g1173(n341 ,n340);
    not g1174(n338 ,n337);
    not g1175(n336 ,n335);
    not g1176(n334 ,n333);
    not g1177(n332 ,n331);
    not g1178(n330 ,n329);
    not g1179(n328 ,n327);
    not g1180(n326 ,n325);
    not g1181(n324 ,n323);
    not g1182(n322 ,n321);
    not g1183(n320 ,n319);
    not g1184(n318 ,n317);
    not g1185(n316 ,n315);
    not g1186(n314 ,n313);
    not g1187(n312 ,n311);
    not g1188(n310 ,n309);
    not g1189(n308 ,n307);
    not g1190(n305 ,n306);
    nor g1191(n304 ,n212 ,n295);
    nor g1192(n363 ,n184 ,n286);
    nor g1193(n361 ,n156 ,n268);
    nor g1194(n360 ,n191 ,n228);
    nor g1195(n359 ,n204 ,n245);
    nor g1196(n358 ,n222 ,n257);
    nor g1197(n357 ,n158 ,n236);
    nor g1198(n356 ,n199 ,n233);
    nor g1199(n355 ,n137 ,n232);
    nor g1200(n354 ,n178 ,n258);
    nor g1201(n353 ,n146 ,n250);
    nor g1202(n352 ,n168 ,n235);
    nor g1203(n351 ,n153 ,n249);
    nor g1204(n350 ,n157 ,n251);
    nor g1205(n348 ,n152 ,n285);
    nor g1206(n346 ,n154 ,n231);
    nor g1207(n344 ,n143 ,n243);
    nor g1208(n342 ,n166 ,n287);
    nor g1209(n340 ,n173 ,n242);
    nor g1210(n339 ,n221 ,n247);
    nor g1211(n337 ,n136 ,n239);
    nor g1212(n335 ,n193 ,n237);
    nor g1213(n333 ,n138 ,n255);
    nor g1214(n331 ,n200 ,n274);
    nor g1215(n329 ,n187 ,n241);
    nor g1216(n327 ,n195 ,n234);
    nor g1217(n325 ,n140 ,n256);
    nor g1218(n323 ,n149 ,n246);
    nor g1219(n321 ,n144 ,n272);
    nor g1220(n319 ,n151 ,n225);
    nor g1221(n317 ,n147 ,n266);
    nor g1222(n315 ,n177 ,n253);
    nor g1223(n313 ,n202 ,n252);
    nor g1224(n311 ,n222 ,n223);
    nor g1225(n309 ,n181 ,n226);
    nor g1226(n307 ,n174 ,n288);
    nor g1227(n306 ,n179 ,n261);
    not g1228(n303 ,n302);
    not g1229(n301 ,n300);
    not g1230(n299 ,n298);
    not g1231(n297 ,n296);
    nor g1232(n294 ,n126 ,n208);
    nor g1233(n293 ,n119 ,n209);
    nor g1234(n292 ,n134 ,n209);
    nor g1235(n291 ,n59 ,n210);
    nor g1236(n290 ,n99 ,n206);
    nor g1237(n289 ,n133 ,n210);
    nor g1238(n288 ,n104 ,n206);
    nor g1239(n287 ,n123 ,n207);
    nor g1240(n286 ,n91 ,n206);
    nor g1241(n285 ,n122 ,n208);
    nor g1242(n284 ,n124 ,n209);
    nor g1243(n283 ,n125 ,n207);
    nor g1244(n282 ,n92 ,n205);
    nor g1245(n281 ,n120 ,n207);
    nor g1246(n280 ,n72 ,n205);
    nor g1247(n279 ,n112 ,n206);
    nor g1248(n278 ,n103 ,n209);
    nor g1249(n277 ,n117 ,n206);
    nor g1250(n276 ,n135 ,n208);
    nor g1251(n275 ,n116 ,n209);
    nor g1252(n274 ,n114 ,n210);
    nor g1253(n273 ,n113 ,n209);
    nor g1254(n272 ,n86 ,n206);
    nor g1255(n271 ,n85 ,n207);
    nor g1256(n270 ,n63 ,n209);
    nor g1257(n269 ,n71 ,n205);
    nor g1258(n268 ,n108 ,n208);
    nor g1259(n267 ,n109 ,n207);
    nor g1260(n266 ,n83 ,n207);
    nor g1261(n265 ,n82 ,n208);
    nor g1262(n264 ,n131 ,n206);
    nor g1263(n263 ,n106 ,n207);
    nor g1264(n262 ,n69 ,n205);
    nor g1265(n302 ,n25 ,n172);
    nor g1266(n300 ,n20 ,n148);
    nor g1267(n298 ,n23 ,n180);
    nor g1268(n296 ,n26 ,n164);
    nor g1269(n295 ,n22 ,n155);
    nor g1270(n261 ,n121 ,n208);
    nor g1271(n260 ,n105 ,n208);
    nor g1272(n259 ,n89 ,n210);
    nor g1273(n258 ,n129 ,n206);
    nor g1274(n257 ,n132 ,n210);
    nor g1275(n256 ,n111 ,n207);
    nor g1276(n255 ,n70 ,n205);
    nor g1277(n254 ,n81 ,n208);
    nor g1278(n253 ,n80 ,n209);
    nor g1279(n252 ,n127 ,n210);
    nor g1280(n251 ,n65 ,n205);
    nor g1281(n250 ,n79 ,n208);
    nor g1282(n249 ,n73 ,n208);
    nor g1283(n248 ,n96 ,n207);
    nor g1284(n247 ,n66 ,n205);
    nor g1285(n246 ,n88 ,n207);
    nor g1286(n245 ,n107 ,n210);
    nor g1287(n244 ,n60 ,n208);
    nor g1288(n243 ,n76 ,n209);
    nor g1289(n242 ,n115 ,n207);
    nor g1290(n241 ,n67 ,n205);
    nor g1291(n240 ,n68 ,n205);
    nor g1292(n239 ,n97 ,n208);
    nor g1293(n238 ,n62 ,n209);
    nor g1294(n237 ,n64 ,n206);
    nor g1295(n236 ,n78 ,n207);
    nor g1296(n235 ,n77 ,n209);
    nor g1297(n234 ,n130 ,n210);
    nor g1298(n233 ,n87 ,n210);
    nor g1299(n232 ,n84 ,n206);
    nor g1300(n231 ,n110 ,n209);
    nor g1301(n230 ,n128 ,n210);
    nor g1302(n228 ,n75 ,n205);
    nor g1303(n227 ,n74 ,n205);
    nor g1304(n226 ,n118 ,n206);
    nor g1305(n225 ,n90 ,n206);
    nor g1306(n224 ,n95 ,n205);
    nor g1307(n223 ,n61 ,n210);
    not g1308(n220 ,n219);
    not g1309(n218 ,n217);
    not g1310(n216 ,n215);
    not g1311(n214 ,n213);
    not g1312(n211 ,n212);
    nor g1313(n204 ,n28 ,n127);
    nor g1314(n203 ,n124 ,n50);
    nor g1315(n202 ,n28 ,n89);
    nor g1316(n201 ,n28 ,n87);
    nor g1317(n200 ,n28 ,n132);
    nor g1318(n199 ,n28 ,n128);
    nor g1319(n198 ,n28 ,n130);
    nor g1320(n197 ,n28 ,n114);
    nor g1321(n195 ,n28 ,n107);
    nor g1322(n194 ,n28 ,n59);
    nor g1323(n193 ,n86 ,n52);
    nor g1324(n192 ,n74 ,n54);
    nor g1325(n191 ,n72 ,n54);
    nor g1326(n190 ,n77 ,n50);
    nor g1327(n189 ,n122 ,n58);
    nor g1328(n188 ,n129 ,n52);
    nor g1329(n187 ,n65 ,n54);
    nor g1330(n186 ,n83 ,n56);
    nor g1331(n185 ,n123 ,n56);
    nor g1332(n184 ,n104 ,n52);
    nor g1333(n183 ,n126 ,n58);
    nor g1334(n182 ,n115 ,n56);
    nor g1335(n181 ,n84 ,n52);
    nor g1336(n180 ,n36 ,n101);
    nor g1337(n179 ,n60 ,n58);
    nor g1338(n178 ,n91 ,n52);
    nor g1339(n177 ,n116 ,n50);
    nor g1340(n222 ,n28 ,n61);
    nor g1341(n221 ,n66 ,n54);
    nor g1342(n219 ,n27 ,n52);
    nor g1343(n217 ,n27 ,n50);
    nor g1344(n215 ,n27 ,n54);
    nor g1345(n213 ,n27 ,n58);
    nor g1346(n212 ,n27 ,n56);
    or g1347(n210 ,n10[0] ,n94);
    or g1348(n209 ,n47 ,n49);
    or g1349(n208 ,n45 ,n57);
    or g1350(n207 ,n46 ,n55);
    or g1351(n206 ,n44 ,n51);
    or g1352(n205 ,n48 ,n53);
    nor g1353(n172 ,n37 ,n93);
    nor g1354(n171 ,n120 ,n56);
    nor g1355(n170 ,n67 ,n54);
    nor g1356(n169 ,n76 ,n50);
    nor g1357(n168 ,n110 ,n50);
    nor g1358(n167 ,n125 ,n56);
    nor g1359(n166 ,n109 ,n56);
    nor g1360(n165 ,n121 ,n58);
    nor g1361(n164 ,n35 ,n98);
    nor g1362(n163 ,n117 ,n52);
    nor g1363(n162 ,n113 ,n50);
    nor g1364(n161 ,n135 ,n58);
    nor g1365(n160 ,n134 ,n50);
    nor g1366(n159 ,n63 ,n50);
    nor g1367(n158 ,n88 ,n56);
    nor g1368(n157 ,n92 ,n54);
    nor g1369(n156 ,n73 ,n58);
    nor g1370(n155 ,n34 ,n100);
    nor g1371(n154 ,n119 ,n50);
    nor g1372(n153 ,n82 ,n58);
    nor g1373(n152 ,n108 ,n58);
    nor g1374(n151 ,n118 ,n52);
    nor g1375(n150 ,n90 ,n52);
    nor g1376(n149 ,n111 ,n56);
    nor g1377(n148 ,n33 ,n102);
    nor g1378(n147 ,n78 ,n56);
    nor g1379(n146 ,n105 ,n58);
    nor g1380(n145 ,n68 ,n54);
    nor g1381(n144 ,n131 ,n52);
    nor g1382(n143 ,n80 ,n50);
    nor g1383(n142 ,n69 ,n54);
    nor g1384(n141 ,n75 ,n54);
    nor g1385(n140 ,n85 ,n56);
    nor g1386(n139 ,n70 ,n54);
    nor g1387(n138 ,n71 ,n54);
    nor g1388(n137 ,n64 ,n52);
    nor g1389(n136 ,n79 ,n58);
    nor g1390(n176 ,n81 ,n58);
    nor g1391(n175 ,n62 ,n50);
    nor g1392(n174 ,n112 ,n52);
    nor g1393(n173 ,n106 ,n56);
    xnor g1394(n103 ,n9[0] ,n10[9]);
    nor g1395(n102 ,n10[5] ,n42);
    nor g1396(n101 ,n10[9] ,n41);
    nor g1397(n100 ,n10[3] ,n40);
    xnor g1398(n99 ,n9[0] ,n10[3]);
    nor g1399(n98 ,n10[7] ,n43);
    xnor g1400(n97 ,n9[0] ,n10[7]);
    xnor g1401(n96 ,n9[0] ,n10[5]);
    xnor g1402(n95 ,n9[0] ,n10[11]);
    nor g1403(n93 ,n10[1] ,n39);
    xnor g1404(n135 ,n10[7] ,n9[3]);
    xnor g1405(n134 ,n10[9] ,n9[2]);
    xnor g1406(n132 ,n10[1] ,n9[10]);
    xnor g1407(n131 ,n10[3] ,n9[6]);
    xnor g1408(n130 ,n10[1] ,n9[5]);
    xnor g1409(n129 ,n10[3] ,n9[8]);
    xnor g1410(n128 ,n10[1] ,n9[4]);
    xnor g1411(n127 ,n10[1] ,n9[7]);
    xnor g1412(n126 ,n10[7] ,n9[10]);
    xnor g1413(n125 ,n10[5] ,n9[9]);
    xnor g1414(n124 ,n10[9] ,n9[10]);
    xnor g1415(n123 ,n10[5] ,n9[7]);
    xnor g1416(n122 ,n10[7] ,n9[4]);
    xnor g1417(n121 ,n10[7] ,n9[8]);
    xnor g1418(n120 ,n10[5] ,n9[6]);
    xnor g1419(n119 ,n10[9] ,n9[8]);
    xnor g1420(n118 ,n10[3] ,n9[2]);
    xnor g1421(n117 ,n10[3] ,n9[7]);
    xnor g1422(n116 ,n10[9] ,n9[5]);
    xnor g1423(n115 ,n10[5] ,n9[10]);
    xnor g1424(n114 ,n10[1] ,n9[9]);
    xnor g1425(n113 ,n10[9] ,n9[1]);
    xnor g1426(n112 ,n10[3] ,n9[11]);
    xnor g1427(n111 ,n10[5] ,n9[4]);
    xnor g1428(n110 ,n10[9] ,n9[7]);
    xnor g1429(n109 ,n10[5] ,n9[8]);
    xnor g1430(n108 ,n10[7] ,n9[5]);
    xnor g1431(n107 ,n10[1] ,n9[6]);
    xnor g1432(n106 ,n10[5] ,n9[11]);
    xnor g1433(n105 ,n10[7] ,n9[2]);
    xnor g1434(n104 ,n10[3] ,n9[10]);
    not g1435(n58 ,n57);
    not g1436(n56 ,n55);
    not g1437(n54 ,n53);
    not g1438(n52 ,n51);
    not g1439(n50 ,n49);
    xnor g1440(n48 ,n10[10] ,n10[11]);
    xnor g1441(n47 ,n10[8] ,n10[9]);
    xnor g1442(n46 ,n10[4] ,n10[5]);
    xnor g1443(n45 ,n10[6] ,n10[7]);
    xnor g1444(n44 ,n10[2] ,n10[3]);
    xnor g1445(n92 ,n10[11] ,n9[6]);
    xnor g1446(n91 ,n10[3] ,n9[9]);
    xnor g1447(n90 ,n10[3] ,n9[1]);
    xnor g1448(n89 ,n10[1] ,n9[8]);
    xnor g1449(n88 ,n10[5] ,n9[3]);
    xnor g1450(n87 ,n10[1] ,n9[3]);
    xnor g1451(n86 ,n10[3] ,n9[5]);
    xnor g1452(n85 ,n10[5] ,n9[5]);
    xnor g1453(n84 ,n10[3] ,n9[3]);
    xnor g1454(n83 ,n10[5] ,n9[1]);
    xnor g1455(n82 ,n10[7] ,n9[7]);
    xnor g1456(n81 ,n10[7] ,n9[11]);
    xnor g1457(n80 ,n10[9] ,n9[4]);
    xnor g1458(n79 ,n10[7] ,n9[1]);
    xnor g1459(n78 ,n10[5] ,n9[2]);
    xnor g1460(n77 ,n10[9] ,n9[6]);
    xnor g1461(n76 ,n10[9] ,n9[3]);
    xnor g1462(n75 ,n10[11] ,n9[7]);
    xnor g1463(n74 ,n10[11] ,n9[9]);
    xnor g1464(n73 ,n10[7] ,n9[6]);
    xnor g1465(n72 ,n10[11] ,n9[8]);
    xnor g1466(n71 ,n10[11] ,n9[3]);
    xnor g1467(n70 ,n10[11] ,n9[2]);
    xnor g1468(n69 ,n10[11] ,n9[10]);
    xnor g1469(n68 ,n10[11] ,n9[1]);
    xnor g1470(n67 ,n10[11] ,n9[4]);
    xnor g1471(n66 ,n10[11] ,n9[11]);
    xnor g1472(n65 ,n10[11] ,n9[5]);
    xnor g1473(n64 ,n10[3] ,n9[4]);
    xnor g1474(n63 ,n10[9] ,n9[9]);
    xnor g1475(n62 ,n10[9] ,n9[11]);
    xnor g1476(n61 ,n10[1] ,n9[11]);
    xnor g1477(n60 ,n10[7] ,n9[9]);
    xnor g1478(n59 ,n10[1] ,n9[2]);
    xnor g1479(n57 ,n10[6] ,n22);
    xnor g1480(n55 ,n10[4] ,n25);
    xnor g1481(n53 ,n10[10] ,n26);
    xnor g1482(n51 ,n10[2] ,n21);
    xnor g1483(n49 ,n10[8] ,n20);
    nor g1484(n43 ,n27 ,n31);
    nor g1485(n42 ,n27 ,n30);
    nor g1486(n41 ,n27 ,n32);
    nor g1487(n40 ,n27 ,n29);
    nor g1488(n39 ,n27 ,n24);
    nor g1489(n37 ,n9[0] ,n10[2]);
    nor g1490(n36 ,n9[0] ,n10[10]);
    nor g1491(n35 ,n9[0] ,n10[8]);
    nor g1492(n34 ,n9[0] ,n10[4]);
    nor g1493(n33 ,n9[0] ,n10[6]);
    not g1494(n32 ,n10[10]);
    not g1495(n31 ,n10[8]);
    not g1496(n30 ,n10[6]);
    not g1497(n29 ,n10[4]);
    not g1498(n28 ,n10[0]);
    not g1499(n27 ,n9[0]);
    not g1500(n26 ,n10[9]);
    not g1501(n25 ,n10[3]);
    not g1502(n24 ,n10[2]);
    not g1503(n23 ,n10[11]);
    not g1504(n22 ,n10[5]);
    not g1505(n21 ,n10[1]);
    not g1506(n20 ,n10[7]);
    or g1507(n17[12] ,n903 ,n944);
    xnor g1508(n18[11] ,n916 ,n943);
    nor g1509(n944 ,n916 ,n943);
    nor g1510(n943 ,n900 ,n942);
    xor g1511(n1771 ,n910 ,n940);
    nor g1512(n942 ,n910 ,n941);
    not g1513(n941 ,n940);
    nor g1514(n940 ,n907 ,n939);
    xor g1515(n1770 ,n917 ,n938);
    nor g1516(n939 ,n917 ,n938);
    nor g1517(n938 ,n897 ,n937);
    xor g1518(n1769 ,n915 ,n936);
    nor g1519(n937 ,n915 ,n936);
    nor g1520(n936 ,n904 ,n935);
    xor g1521(n1768 ,n919 ,n934);
    nor g1522(n935 ,n919 ,n934);
    nor g1523(n934 ,n905 ,n933);
    xnor g1524(n1767 ,n918 ,n931);
    nor g1525(n933 ,n918 ,n932);
    not g1526(n932 ,n931);
    nor g1527(n931 ,n899 ,n930);
    xor g1528(n1766 ,n911 ,n928);
    nor g1529(n930 ,n911 ,n929);
    not g1530(n929 ,n928);
    nor g1531(n928 ,n906 ,n927);
    xnor g1532(n1765 ,n914 ,n925);
    nor g1533(n927 ,n914 ,n926);
    not g1534(n926 ,n925);
    nor g1535(n925 ,n898 ,n924);
    xnor g1536(n1764 ,n909 ,n923);
    nor g1537(n924 ,n909 ,n923);
    nor g1538(n923 ,n896 ,n922);
    xnor g1539(n1763 ,n913 ,n921);
    nor g1540(n922 ,n913 ,n921);
    nor g1541(n921 ,n901 ,n920);
    xnor g1542(n1762 ,n912 ,n908);
    nor g1543(n920 ,n908 ,n912);
    nor g1544(n1761 ,n908 ,n902);
    xnor g1545(n919 ,n9[7] ,n10[7]);
    xnor g1546(n918 ,n9[6] ,n10[6]);
    xnor g1547(n917 ,n9[9] ,n10[9]);
    xnor g1548(n916 ,n9[11] ,n10[11]);
    xnor g1549(n915 ,n9[8] ,n10[8]);
    xnor g1550(n914 ,n9[4] ,n10[4]);
    xnor g1551(n913 ,n9[2] ,n10[2]);
    xnor g1552(n912 ,n9[1] ,n10[1]);
    xnor g1553(n911 ,n9[5] ,n10[5]);
    xnor g1554(n910 ,n9[10] ,n10[10]);
    xnor g1555(n909 ,n9[3] ,n10[3]);
    nor g1556(n907 ,n894 ,n888);
    nor g1557(n906 ,n889 ,n890);
    nor g1558(n905 ,n891 ,n885);
    nor g1559(n904 ,n882 ,n883);
    nor g1560(n903 ,n886 ,n884);
    nor g1561(n908 ,n895 ,n892);
    nor g1562(n902 ,n9[0] ,n10[0]);
    nor g1563(n901 ,n9[1] ,n10[1]);
    nor g1564(n900 ,n9[10] ,n10[10]);
    nor g1565(n899 ,n9[5] ,n10[5]);
    nor g1566(n898 ,n9[3] ,n10[3]);
    nor g1567(n897 ,n887 ,n893);
    nor g1568(n896 ,n9[2] ,n10[2]);
    not g1569(n895 ,n9[0]);
    not g1570(n894 ,n9[9]);
    not g1571(n893 ,n10[8]);
    not g1572(n892 ,n10[0]);
    not g1573(n891 ,n9[6]);
    not g1574(n890 ,n10[4]);
    not g1575(n889 ,n9[4]);
    not g1576(n888 ,n10[9]);
    not g1577(n887 ,n9[8]);
    not g1578(n886 ,n9[11]);
    not g1579(n885 ,n10[6]);
    not g1580(n884 ,n10[11]);
    not g1581(n883 ,n10[7]);
    not g1582(n882 ,n9[7]);
    xnor g1583(n14[17] ,n13[17] ,n1027);
    xnor g1584(n14[16] ,n13[16] ,n1024);
    nor g1585(n1027 ,n1026 ,n1025);
    xnor g1586(n14[15] ,n13[15] ,n1020);
    nor g1587(n1026 ,n946 ,n1023);
    nor g1588(n1024 ,n1022 ,n1021);
    xnor g1589(n14[14] ,n13[14] ,n1016);
    not g1590(n1023 ,n1022);
    nor g1591(n1022 ,n945 ,n1019);
    nor g1592(n1020 ,n1018 ,n1017);
    xnor g1593(n14[13] ,n13[13] ,n1012);
    not g1594(n1019 ,n1018);
    nor g1595(n1018 ,n951 ,n1015);
    nor g1596(n1016 ,n1014 ,n1013);
    xnor g1597(n14[12] ,n13[12] ,n1008);
    not g1598(n1015 ,n1014);
    nor g1599(n1014 ,n950 ,n1011);
    nor g1600(n1012 ,n1010 ,n1009);
    not g1601(n1011 ,n1010);
    nor g1602(n1010 ,n949 ,n1006);
    nor g1603(n1008 ,n1005 ,n1007);
    xor g1604(n14[11] ,n978 ,n1003);
    nor g1605(n1007 ,n967 ,n1004);
    not g1606(n1006 ,n1005);
    nor g1607(n1005 ,n966 ,n1003);
    not g1608(n1004 ,n1003);
    nor g1609(n1003 ,n969 ,n1002);
    xor g1610(n1749 ,n982 ,n1001);
    nor g1611(n1002 ,n982 ,n1001);
    nor g1612(n1001 ,n968 ,n1000);
    xnor g1613(n1748 ,n981 ,n998);
    nor g1614(n1000 ,n981 ,n999);
    not g1615(n999 ,n998);
    nor g1616(n998 ,n959 ,n997);
    xnor g1617(n1747 ,n974 ,n996);
    nor g1618(n997 ,n974 ,n996);
    nor g1619(n996 ,n958 ,n995);
    xnor g1620(n1746 ,n976 ,n994);
    nor g1621(n995 ,n976 ,n994);
    nor g1622(n994 ,n962 ,n993);
    xnor g1623(n1745 ,n975 ,n992);
    nor g1624(n993 ,n975 ,n992);
    nor g1625(n992 ,n965 ,n991);
    xnor g1626(n1744 ,n973 ,n990);
    nor g1627(n991 ,n973 ,n990);
    nor g1628(n990 ,n963 ,n989);
    xnor g1629(n1743 ,n972 ,n988);
    nor g1630(n989 ,n972 ,n988);
    nor g1631(n988 ,n961 ,n987);
    xnor g1632(n1742 ,n980 ,n986);
    nor g1633(n987 ,n980 ,n986);
    nor g1634(n986 ,n960 ,n985);
    xnor g1635(n1741 ,n979 ,n984);
    nor g1636(n985 ,n979 ,n984);
    nor g1637(n984 ,n970 ,n983);
    xnor g1638(n1740 ,n977 ,n971);
    nor g1639(n983 ,n971 ,n977);
    nor g1640(n1739 ,n971 ,n964);
    xnor g1641(n978 ,n13[11] ,n12[11]);
    xnor g1642(n982 ,n1782 ,n12[10]);
    xnor g1643(n981 ,n1781 ,n12[9]);
    xnor g1644(n980 ,n1775 ,n12[3]);
    xnor g1645(n979 ,n1774 ,n12[2]);
    xnor g1646(n977 ,n1773 ,n12[1]);
    xnor g1647(n976 ,n1779 ,n12[7]);
    xnor g1648(n975 ,n1778 ,n12[6]);
    xnor g1649(n974 ,n1780 ,n12[8]);
    xnor g1650(n973 ,n1777 ,n12[5]);
    xnor g1651(n972 ,n1776 ,n12[4]);
    nor g1652(n970 ,n1773 ,n12[1]);
    nor g1653(n969 ,n957 ,n956);
    nor g1654(n968 ,n952 ,n948);
    or g1655(n967 ,n953 ,n13[11]);
    or g1656(n966 ,n955 ,n12[11]);
    nor g1657(n965 ,n1777 ,n12[5]);
    nor g1658(n971 ,n954 ,n947);
    nor g1659(n964 ,n1772 ,n12[0]);
    nor g1660(n963 ,n1776 ,n12[4]);
    nor g1661(n962 ,n1778 ,n12[6]);
    nor g1662(n961 ,n1775 ,n12[3]);
    nor g1663(n960 ,n1774 ,n12[2]);
    nor g1664(n959 ,n1780 ,n12[8]);
    nor g1665(n958 ,n1779 ,n12[7]);
    not g1666(n957 ,n1782);
    not g1667(n956 ,n12[10]);
    not g1668(n955 ,n13[11]);
    not g1669(n954 ,n1772);
    not g1670(n953 ,n12[11]);
    not g1671(n952 ,n1781);
    not g1672(n951 ,n13[14]);
    not g1673(n950 ,n13[13]);
    not g1674(n949 ,n13[12]);
    not g1675(n948 ,n12[9]);
    not g1676(n947 ,n12[0]);
    not g1677(n946 ,n13[16]);
    not g1678(n945 ,n13[15]);
    nor g1679(n1694 ,n1061 ,n1094);
    nor g1680(n1094 ,n1076 ,n1093);
    nor g1681(n1093 ,n1078 ,n1092);
    nor g1682(n1092 ,n1083 ,n1091);
    nor g1683(n1091 ,n1080 ,n1090);
    nor g1684(n1090 ,n1075 ,n1089);
    nor g1685(n1089 ,n1084 ,n1088);
    nor g1686(n1088 ,n1081 ,n1087);
    nor g1687(n1087 ,n1079 ,n1086);
    nor g1688(n1086 ,n1077 ,n1085);
    nor g1689(n1085 ,n1074 ,n1082);
    or g1690(n1084 ,n1067 ,n1065);
    or g1691(n1083 ,n1066 ,n1064);
    or g1692(n1082 ,n1073 ,n1072);
    or g1693(n1081 ,n1063 ,n1056);
    or g1694(n1080 ,n1057 ,n1055);
    or g1695(n1079 ,n1058 ,n1060);
    or g1696(n1078 ,n1062 ,n1068);
    or g1697(n1077 ,n1054 ,n1053);
    or g1698(n1076 ,n1052 ,n1069);
    or g1699(n1075 ,n1051 ,n1070);
    nor g1700(n1074 ,n1059 ,n1071);
    nor g1701(n1073 ,n1046 ,n1718);
    nor g1702(n1072 ,n1028 ,n1717);
    nor g1703(n1071 ,n1050 ,n10[0]);
    nor g1704(n1070 ,n1033 ,n1700);
    nor g1705(n1069 ,n1042 ,n1704);
    nor g1706(n1068 ,n1043 ,n1725);
    nor g1707(n1067 ,n1035 ,n1722);
    nor g1708(n1066 ,n1047 ,n1703);
    nor g1709(n1065 ,n1037 ,n1721);
    nor g1710(n1064 ,n1030 ,n1702);
    nor g1711(n1063 ,n1048 ,n1699);
    nor g1712(n1062 ,n1036 ,n1726);
    nor g1713(n1061 ,n1045 ,n1727);
    nor g1714(n1060 ,n1041 ,n1719);
    nor g1715(n1059 ,n1039 ,n1695);
    nor g1716(n1058 ,n1034 ,n1720);
    nor g1717(n1057 ,n1044 ,n1724);
    nor g1718(n1056 ,n1031 ,n1698);
    nor g1719(n1055 ,n1049 ,n1723);
    nor g1720(n1054 ,n1032 ,n1697);
    nor g1721(n1053 ,n1029 ,n1696);
    nor g1722(n1052 ,n1038 ,n1705);
    nor g1723(n1051 ,n1040 ,n1701);
    not g1724(n1050 ,n9[0]);
    not g1725(n1049 ,n1701);
    not g1726(n1048 ,n1721);
    not g1727(n1047 ,n1725);
    not g1728(n1046 ,n1696);
    not g1729(n1045 ,n1705);
    not g1730(n1044 ,n1702);
    not g1731(n1043 ,n1703);
    not g1732(n1042 ,n1726);
    not g1733(n1041 ,n1697);
    not g1734(n1040 ,n1723);
    not g1735(n1039 ,n1717);
    not g1736(n1038 ,n1727);
    not g1737(n1037 ,n1699);
    not g1738(n1036 ,n1704);
    not g1739(n1035 ,n1700);
    not g1740(n1034 ,n1698);
    not g1741(n1033 ,n1722);
    not g1742(n1032 ,n1719);
    not g1743(n1031 ,n1720);
    not g1744(n1030 ,n1724);
    not g1745(n1029 ,n1718);
    not g1746(n1028 ,n1695);
    xnor g1747(n1737 ,n9[10] ,n1112);
    nor g1748(n1114 ,n9[10] ,n1113);
    xnor g1749(n1736 ,n9[9] ,n1110);
    not g1750(n1113 ,n1112);
    nor g1751(n1112 ,n9[9] ,n1111);
    xnor g1752(n1735 ,n9[8] ,n1108);
    not g1753(n1111 ,n1110);
    nor g1754(n1110 ,n9[8] ,n1109);
    xnor g1755(n1734 ,n9[7] ,n1106);
    not g1756(n1109 ,n1108);
    nor g1757(n1108 ,n9[7] ,n1107);
    xnor g1758(n1733 ,n9[6] ,n1104);
    not g1759(n1107 ,n1106);
    nor g1760(n1106 ,n9[6] ,n1105);
    xnor g1761(n1732 ,n9[5] ,n1102);
    not g1762(n1105 ,n1104);
    nor g1763(n1104 ,n9[5] ,n1103);
    xnor g1764(n1731 ,n9[4] ,n1100);
    not g1765(n1103 ,n1102);
    nor g1766(n1102 ,n9[4] ,n1101);
    xnor g1767(n1730 ,n9[3] ,n1098);
    not g1768(n1101 ,n1100);
    nor g1769(n1100 ,n9[3] ,n1099);
    xnor g1770(n1729 ,n9[2] ,n1096);
    not g1771(n1099 ,n1098);
    nor g1772(n1098 ,n9[2] ,n1097);
    xor g1773(n1728 ,n9[1] ,n9[0]);
    not g1774(n1097 ,n1096);
    nor g1775(n1096 ,n9[1] ,n9[0]);
    xnor g1776(n1715 ,n10[10] ,n1131);
    nor g1777(n1133 ,n10[10] ,n1132);
    xnor g1778(n1714 ,n10[9] ,n1129);
    not g1779(n1132 ,n1131);
    nor g1780(n1131 ,n10[9] ,n1130);
    xnor g1781(n1713 ,n10[8] ,n1127);
    not g1782(n1130 ,n1129);
    nor g1783(n1129 ,n10[8] ,n1128);
    xnor g1784(n1712 ,n10[7] ,n1125);
    not g1785(n1128 ,n1127);
    nor g1786(n1127 ,n10[7] ,n1126);
    xnor g1787(n1711 ,n10[6] ,n1123);
    not g1788(n1126 ,n1125);
    nor g1789(n1125 ,n10[6] ,n1124);
    xnor g1790(n1710 ,n10[5] ,n1121);
    not g1791(n1124 ,n1123);
    nor g1792(n1123 ,n10[5] ,n1122);
    xnor g1793(n1709 ,n10[4] ,n1119);
    not g1794(n1122 ,n1121);
    nor g1795(n1121 ,n10[4] ,n1120);
    xnor g1796(n1708 ,n10[3] ,n1117);
    not g1797(n1120 ,n1119);
    nor g1798(n1119 ,n10[3] ,n1118);
    xnor g1799(n1707 ,n10[2] ,n1115);
    not g1800(n1118 ,n1117);
    nor g1801(n1117 ,n10[2] ,n1116);
    xor g1802(n1706 ,n10[1] ,n10[0]);
    not g1803(n1116 ,n1115);
    nor g1804(n1115 ,n10[1] ,n10[0]);
    or g1805(n15[12] ,n1799 ,n1851);
    xor g1806(n16[11] ,n1850 ,n1815);
    nor g1807(n1851 ,n1816 ,n1850);
    nor g1808(n1850 ,n1798 ,n1849);
    xor g1809(n1760 ,n1848 ,n1817);
    nor g1810(n1849 ,n1818 ,n1848);
    nor g1811(n1848 ,n1808 ,n1847);
    xor g1812(n1759 ,n1846 ,n1819);
    nor g1813(n1847 ,n1820 ,n1846);
    nor g1814(n1846 ,n1796 ,n1845);
    xor g1815(n1758 ,n1844 ,n1813);
    nor g1816(n1845 ,n1814 ,n1844);
    nor g1817(n1844 ,n1805 ,n1843);
    xor g1818(n1757 ,n1842 ,n1827);
    nor g1819(n1843 ,n1828 ,n1842);
    nor g1820(n1842 ,n1803 ,n1841);
    xor g1821(n1756 ,n1840 ,n1823);
    nor g1822(n1841 ,n1824 ,n1840);
    nor g1823(n1840 ,n1797 ,n1839);
    xor g1824(n1755 ,n1838 ,n1821);
    nor g1825(n1839 ,n1822 ,n1838);
    nor g1826(n1838 ,n1806 ,n1837);
    xor g1827(n1754 ,n1836 ,n1811);
    nor g1828(n1837 ,n1812 ,n1836);
    nor g1829(n1836 ,n1800 ,n1835);
    xor g1830(n1753 ,n1834 ,n1809);
    nor g1831(n1835 ,n1810 ,n1834);
    nor g1832(n1834 ,n1807 ,n1833);
    xor g1833(n1752 ,n1832 ,n1829);
    nor g1834(n1833 ,n1830 ,n1832);
    nor g1835(n1832 ,n1804 ,n1831);
    xnor g1836(n1751 ,n1825 ,n1801);
    nor g1837(n1831 ,n1802 ,n1826);
    not g1838(n1830 ,n1829);
    not g1839(n1828 ,n1827);
    not g1840(n1826 ,n1825);
    not g1841(n1824 ,n1823);
    not g1842(n1822 ,n1821);
    xor g1843(n1750 ,n9[0] ,n10[0]);
    xnor g1844(n1829 ,n9[2] ,n10[2]);
    xnor g1845(n1827 ,n9[7] ,n10[7]);
    xnor g1846(n1825 ,n9[1] ,n10[1]);
    xnor g1847(n1823 ,n9[6] ,n10[6]);
    xnor g1848(n1821 ,n9[5] ,n10[5]);
    not g1849(n1820 ,n1819);
    not g1850(n1818 ,n1817);
    not g1851(n1816 ,n1815);
    not g1852(n1814 ,n1813);
    not g1853(n1812 ,n1811);
    not g1854(n1810 ,n1809);
    xnor g1855(n1819 ,n9[9] ,n10[9]);
    xnor g1856(n1817 ,n9[10] ,n10[10]);
    xnor g1857(n1815 ,n9[11] ,n10[11]);
    xnor g1858(n1813 ,n9[8] ,n10[8]);
    xnor g1859(n1811 ,n9[4] ,n10[4]);
    xnor g1860(n1809 ,n9[3] ,n10[3]);
    nor g1861(n1808 ,n1784 ,n9[9]);
    nor g1862(n1807 ,n1785 ,n9[2]);
    nor g1863(n1806 ,n1790 ,n9[4]);
    nor g1864(n1805 ,n1793 ,n9[7]);
    nor g1865(n1804 ,n1786 ,n9[1]);
    nor g1866(n1803 ,n1789 ,n9[6]);
    not g1867(n1802 ,n1801);
    nor g1868(n1800 ,n1795 ,n9[3]);
    nor g1869(n1799 ,n1791 ,n10[11]);
    nor g1870(n1798 ,n1792 ,n9[10]);
    nor g1871(n1797 ,n1787 ,n9[5]);
    nor g1872(n1796 ,n1788 ,n9[8]);
    nor g1873(n1801 ,n1794 ,n9[0]);
    not g1874(n1795 ,n10[3]);
    not g1875(n1794 ,n10[0]);
    not g1876(n1793 ,n10[7]);
    not g1877(n1792 ,n10[10]);
    not g1878(n1791 ,n9[11]);
    not g1879(n1790 ,n10[4]);
    not g1880(n1789 ,n10[6]);
    not g1881(n1788 ,n10[8]);
    not g1882(n1787 ,n10[5]);
    not g1883(n1786 ,n10[1]);
    not g1884(n1785 ,n10[2]);
    not g1885(n1784 ,n10[9]);
    buf g1886(n133 ,n9[1]);
    not g1887(n94 ,n10[1]);
    buf g1888(n38 ,n9[0]);
    not g1889(n196 ,n133);
    not g1890(n229 ,n210);
    buf g1891(n463 ,n424);
    not g1892(n541 ,n425);
    buf g1893(n1716 ,n1133);
    buf g1894(n1738 ,n1114);
    buf g1895(n1009 ,n1007);
    buf g1896(n1013 ,n1009);
    buf g1897(n1340 ,n1325);
    buf g1898(n1017 ,n1013);
    buf g1899(n1021 ,n1017);
    buf g1900(n1025 ,n1021);
    buf g1901(n1419 ,n1316);
    buf g1902(n1472 ,n1341);
    buf g1903(n1323 ,n1301);
    not g1904(n1868 ,n19[0]);
    not g1905(n1867 ,n19[2]);
    not g1906(n1866 ,n19[1]);
    nor g1907(n1872 ,n1864 ,n1865);
    nor g1908(n1871 ,n1864 ,n1867);
    nor g1909(n1869 ,n1864 ,n1868);
    nor g1910(n1870 ,n1864 ,n1866);
    not g1911(n1865 ,n1877);
    not g1912(n1864 ,n1783);
    dff g1913(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n19[0]));
    dff g1914(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n19[1]));
    dff g1915(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n19[2]));
    dff g1916(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n1877));
    xor g1917(n1873 ,n1872 ,n1863);
    nor g1918(n1874 ,n1862 ,n1863);
    nor g1919(n1863 ,n1853 ,n1861);
    nor g1920(n1862 ,n1871 ,n1860);
    nor g1921(n1875 ,n1859 ,n1860);
    not g1922(n1861 ,n1860);
    nor g1923(n1860 ,n1855 ,n1858);
    nor g1924(n1859 ,n1870 ,n1857);
    nor g1925(n1876 ,n1857 ,n1856);
    not g1926(n1858 ,n1857);
    nor g1927(n1857 ,n1852 ,n1854);
    nor g1928(n1856 ,n1869 ,n9[0]);
    not g1929(n1855 ,n1870);
    not g1930(n1854 ,n9[0]);
    not g1931(n1853 ,n1871);
    not g1932(n1852 ,n1869);
endmodule
