module top (n0, n1, n2, n3, n4);
    input n0, n1;
    input [63:0] n2;
    input [7:0] n3;
    output [31:0] n4;
    wire n0, n1;
    wire [63:0] n2;
    wire [7:0] n3;
    wire [31:0] n4;
    wire [7:0] n5;
    wire [31:0] n6;
    wire [15:0] n7;
    wire [7:0] n8;
    wire [15:0] n9;
    wire [15:0] n10;
    wire [7:0] n11;
    wire [3:0] n12;
    wire [15:0] n13;
    wire [7:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581;
    nor g0(n294 ,n126 ,n285);
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n354), .Q(n6[14]));
    not g2(n471 ,n14[6]);
    nor g3(n352 ,n13[0] ,n322);
    xor g4(n7[9] ,n2[25] ,n2[9]);
    nor g5(n251 ,n156 ,n209);
    or g6(n513 ,n558 ,n7[14]);
    not g7(n152 ,n2[0]);
    not g8(n476 ,n14[5]);
    or g9(n539 ,n558 ,n499);
    not g10(n385 ,n5[3]);
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n242), .Q(n10[12]));
    not g12(n390 ,n406);
    not g13(n101 ,n100);
    buf g14(n4[18], n4[31]);
    nor g15(n325 ,n137 ,n307);
    or g16(n199 ,n197 ,n9[6]);
    nor g17(n247 ,n164 ,n209);
    nor g18(n573 ,n434 ,n435);
    not g19(n170 ,n391);
    nor g20(n269 ,n143 ,n257);
    nor g21(n266 ,n174 ,n260);
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n245), .Q(n10[7]));
    nor g23(n225 ,n189 ,n126);
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n303), .Q(n8[0]));
    not g25(n155 ,n408);
    or g26(n38 ,n8[4] ,n37);
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n296), .Q(n8[5]));
    not g28(n51 ,n50);
    nor g29(n114 ,n10[13] ,n112);
    or g30(n364 ,n329 ,n348);
    dff g31(.RN(n520), .SN(n537), .CK(n0), .D(n569), .Q(n13[6]));
    nor g32(n81 ,n10[2] ,n79);
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n295), .Q(n8[6]));
    not g34(n73 ,n10[11]);
    nor g35(n435 ,n416 ,n433);
    not g36(n473 ,n14[4]);
    dff g37(.RN(n558), .SN(1'b1), .CK(n0), .D(n577), .Q(n14[5]));
    nor g38(n370 ,n126 ,n334);
    nor g39(n440 ,n417 ,n438);
    not g40(n544 ,n14[2]);
    not g41(n427 ,n7[10]);
    not g42(n426 ,n7[8]);
    xnor g43(n378 ,n9[0] ,n10[0]);
    nor g44(n220 ,n126 ,n152);
    xnor g45(n124 ,n2[5] ,n3[5]);
    not g46(n86 ,n85);
    or g47(n535 ,n558 ,n506);
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n225), .Q(n5[3]));
    nor g49(n411 ,n52 ,n53);
    nor g50(n434 ,n7[2] ,n432);
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n250), .Q(n10[1]));
    or g52(n304 ,n126 ,n301);
    xor g53(n7[11] ,n2[27] ,n2[11]);
    xnor g54(n120 ,n2[1] ,n3[1]);
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n203), .Q(n11[3]));
    nor g56(n398 ,n99 ,n100);
    nor g57(n289 ,n269 ,n270);
    or g58(n371 ,n333 ,n347);
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n254), .Q(n10[15]));
    nor g60(n491 ,n476 ,n489);
    nor g61(n410 ,n55 ,n56);
    not g62(n68 ,n10[5]);
    nor g63(n91 ,n68 ,n89);
    nor g64(n253 ,n161 ,n209);
    not g65(n418 ,n7[6]);
    not g66(n113 ,n112);
    nor g67(n52 ,n8[3] ,n50);
    not g68(n416 ,n7[2]);
    nor g69(n432 ,n430 ,n425);
    nor g70(n291 ,n273 ,n280);
    xnor g71(n7[6] ,n2[22] ,n125);
    nor g72(n302 ,n215 ,n284);
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n232), .Q(n9[3]));
    not g74(n145 ,n415);
    not g75(n30 ,n8[1]);
    nor g76(n334 ,n313 ,n310);
    not g77(n104 ,n103);
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n205), .Q(n9[6]));
    xnor g79(n123 ,n2[7] ,n3[7]);
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n249), .Q(n10[2]));
    or g81(n519 ,n558 ,n7[15]);
    nor g82(n323 ,n140 ,n307);
    nor g83(n562 ,n466 ,n467);
    not g84(n307 ,n306);
    or g85(n37 ,n8[7] ,n36);
    not g86(n176 ,n9[0]);
    dff g87(.RN(n514), .SN(n530), .CK(n0), .D(n562), .Q(n13[13]));
    nor g88(n412 ,n49 ,n50);
    xnor g89(n4[13] ,n384 ,n6[13]);
    not g90(n502 ,n7[9]);
    nor g91(n281 ,n167 ,n256);
    or g92(n198 ,n190 ,n9[2]);
    nor g93(n559 ,n554 ,n557);
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n241), .Q(n10[13]));
    not g95(n140 ,n13[11]);
    not g96(n501 ,n7[13]);
    not g97(n74 ,n10[14]);
    dff g98(.RN(n558), .SN(1'b1), .CK(n0), .D(n580), .Q(n14[2]));
    nor g99(n223 ,n176 ,n126);
    or g100(n264 ,n214 ,n237);
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n8[1]));
    dff g102(.RN(n517), .SN(n534), .CK(n0), .D(n566), .Q(n13[9]));
    xnor g103(n376 ,n2[0] ,n3[0]);
    or g104(n382 ,n388 ,n380);
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n229), .Q(n5[4]));
    or g106(n543 ,n558 ,n510);
    not g107(n161 ,n401);
    not g108(n506 ,n7[8]);
    or g109(n365 ,n330 ,n349);
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n5[0]));
    nor g111(n111 ,n10[12] ,n109);
    nor g112(n445 ,n7[6] ,n443);
    xor g113(n7[8] ,n2[24] ,n2[8]);
    xnor g114(n4[10] ,n384 ,n6[10]);
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n321), .Q(n6[16]));
    nor g116(n82 ,n67 ,n80);
    nor g117(n564 ,n460 ,n461);
    not g118(n496 ,n7[11]);
    not g119(n456 ,n455);
    not g120(n558 ,n1);
    or g121(n293 ,n266 ,n290);
    nor g122(n395 ,n90 ,n91);
    or g123(n18 ,n10[7] ,n10[6]);
    nor g124(n55 ,n8[4] ,n53);
    nor g125(n87 ,n10[4] ,n85);
    not g126(n67 ,n10[2]);
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n204), .Q(n9[7]));
    not g128(n48 ,n47);
    xor g129(n7[15] ,n2[31] ,n2[15]);
    nor g130(n466 ,n7[13] ,n464);
    not g131(n95 ,n94);
    not g132(n188 ,n9[2]);
    nor g133(n315 ,n173 ,n308);
    nor g134(n284 ,n216 ,n265);
    or g135(n522 ,n558 ,n7[5]);
    not g136(n187 ,n5[4]);
    not g137(n489 ,n488);
    xnor g138(n4[5] ,n384 ,n6[5]);
    nor g139(n292 ,n272 ,n281);
    not g140(n441 ,n440);
    xnor g141(n4[11] ,n384 ,n6[11]);
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n206), .Q(n11[0]));
    nor g143(n262 ,n231 ,n239);
    nor g144(n100 ,n69 ,n98);
    nor g145(n341 ,n13[11] ,n322);
    or g146(n217 ,n175 ,n169);
    nor g147(n338 ,n13[14] ,n322);
    buf g148(n4[28], n4[31]);
    or g149(n24 ,n22 ,n19);
    or g150(n362 ,n327 ,n346);
    not g151(n507 ,n7[5]);
    not g152(n138 ,n13[7]);
    nor g153(n479 ,n475 ,n472);
    xnor g154(n122 ,n2[4] ,n3[4]);
    nor g155(n340 ,n13[12] ,n322);
    not g156(n308 ,n309);
    nor g157(n310 ,n263 ,n309);
    nor g158(n296 ,n126 ,n287);
    nor g159(n577 ,n490 ,n491);
    nor g160(n470 ,n423 ,n468);
    nor g161(n574 ,n432 ,n431);
    nor g162(n53 ,n42 ,n51);
    not g163(n131 ,n13[12]);
    nor g164(n59 ,n44 ,n57);
    or g165(n527 ,n558 ,n7[0]);
    nor g166(n36 ,n32 ,n35);
    not g167(n486 ,n485);
    nor g168(n201 ,n185 ,n126);
    nor g169(n350 ,n13[2] ,n322);
    not g170(n40 ,n8[0]);
    not g171(n545 ,n14[0]);
    xnor g172(n7[1] ,n2[17] ,n120);
    nor g173(n347 ,n13[5] ,n322);
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n219), .Q(n9[2]));
    not g175(n150 ,n392);
    xor g176(n7[13] ,n2[29] ,n2[13]);
    dff g177(.RN(n525), .SN(n543), .CK(n0), .D(n573), .Q(n13[2]));
    not g178(n211 ,n210);
    nor g179(n115 ,n64 ,n113);
    not g180(n172 ,n12[1]);
    nor g181(n286 ,n268 ,n276);
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n297), .Q(n8[4]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n11[1]));
    nor g184(n34 ,n30 ,n31);
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n222), .Q(n5[2]));
    nor g186(n327 ,n147 ,n307);
    buf g187(n4[24], n4[31]);
    nor g188(n260 ,n145 ,n213);
    nor g189(n324 ,n141 ,n307);
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n246), .Q(n10[6]));
    not g191(n428 ,n7[7]);
    or g192(n305 ,n258 ,n293);
    nor g193(n216 ,n128 ,n12[1]);
    or g194(n283 ,n12[2] ,n262);
    dff g195(.RN(n558), .SN(1'b1), .CK(n0), .D(n576), .Q(n14[6]));
    dff g196(.RN(n522), .SN(n538), .CK(n0), .D(n570), .Q(n13[5]));
    or g197(n541 ,n558 ,n504);
    nor g198(n485 ,n474 ,n483);
    or g199(n360 ,n325 ,n344);
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n357), .Q(n6[11]));
    nor g201(n330 ,n130 ,n307);
    not g202(n171 ,n398);
    nor g203(n278 ,n154 ,n256);
    or g204(n239 ,n12[0] ,n216);
    xor g205(n383 ,n415 ,n381);
    nor g206(n255 ,n145 ,n214);
    or g207(n361 ,n326 ,n345);
    not g208(n549 ,n14[1]);
    xnor g209(n4[8] ,n384 ,n6[8]);
    nor g210(n481 ,n14[2] ,n479);
    not g211(n422 ,n7[9]);
    nor g212(n118 ,n74 ,n116);
    nor g213(n50 ,n45 ,n48);
    nor g214(n403 ,n114 ,n115);
    not g215(n425 ,n559);
    xnor g216(n7[0] ,n2[16] ,n376);
    not g217(n387 ,n5[7]);
    nor g218(n446 ,n418 ,n444);
    nor g219(n487 ,n14[4] ,n485);
    buf g220(n4[23], n4[31]);
    nor g221(n280 ,n153 ,n256);
    nor g222(n221 ,n175 ,n126);
    not g223(n70 ,n10[7]);
    xnor g224(n4[15] ,n384 ,n6[15]);
    nor g225(n272 ,n191 ,n257);
    buf g226(n4[19], n4[31]);
    nor g227(n265 ,n217 ,n259);
    nor g228(n460 ,n7[11] ,n458);
    not g229(n60 ,n59);
    xnor g230(n4[2] ,n384 ,n6[2]);
    or g231(n557 ,n546 ,n556);
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n362), .Q(n6[6]));
    dff g233(.RN(n519), .SN(n528), .CK(n0), .D(n560), .Q(n13[15]));
    not g234(n420 ,n7[11]);
    nor g235(n35 ,n8[2] ,n34);
    nor g236(n463 ,n7[12] ,n461);
    not g237(n511 ,n7[15]);
    nor g238(n580 ,n481 ,n482);
    not g239(n178 ,n5[3]);
    xor g240(n560 ,n7[15] ,n470);
    nor g241(n342 ,n13[10] ,n322);
    not g242(n141 ,n13[9]);
    not g243(n510 ,n7[2]);
    xnor g244(n384 ,n377 ,n383);
    not g245(n179 ,n9[1]);
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n356), .Q(n6[12]));
    not g247(n181 ,n9[6]);
    nor g248(n457 ,n7[10] ,n455);
    xnor g249(n381 ,n378 ,n8[0]);
    nor g250(n243 ,n158 ,n209);
    not g251(n127 ,n13[0]);
    nor g252(n299 ,n126 ,n292);
    nor g253(n207 ,n144 ,n126);
    not g254(n500 ,n7[7]);
    nor g255(n316 ,n127 ,n307);
    not g256(n130 ,n13[3]);
    or g257(n529 ,n558 ,n497);
    or g258(n21 ,n10[15] ,n10[14]);
    nor g259(n254 ,n159 ,n209);
    dff g260(.RN(n521), .SN(n536), .CK(n0), .D(n568), .Q(n13[7]));
    or g261(n553 ,n547 ,n544);
    not g262(n136 ,n13[5]);
    not g263(n143 ,n8[3]);
    buf g264(n4[25], n4[31]);
    not g265(n509 ,n14[0]);
    or g266(n29 ,n10[13] ,n28);
    nor g267(n402 ,n111 ,n112);
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n253), .Q(n10[11]));
    nor g269(n565 ,n457 ,n458);
    not g270(n92 ,n91);
    nor g271(n312 ,n236 ,n309);
    not g272(n57 ,n56);
    xnor g273(n4[9] ,n384 ,n6[9]);
    nor g274(n571 ,n439 ,n440);
    nor g275(n240 ,n151 ,n209);
    xnor g276(n377 ,n11[0] ,n12[0]);
    nor g277(n106 ,n75 ,n104);
    or g278(n537 ,n558 ,n503);
    not g279(n472 ,n14[0]);
    dff g280(.RN(n516), .SN(n533), .CK(n0), .D(n565), .Q(n13[10]));
    not g281(n195 ,n11[2]);
    nor g282(n46 ,n8[1] ,n8[0]);
    nor g283(n581 ,n479 ,n478);
    nor g284(n568 ,n448 ,n449);
    not g285(n429 ,n7[12]);
    dff g286(.RN(n558), .SN(1'b1), .CK(n0), .D(n509), .Q(n14[0]));
    nor g287(n242 ,n163 ,n209);
    nor g288(n570 ,n442 ,n443);
    nor g289(n320 ,n174 ,n308);
    not g290(n388 ,n5[1]);
    nor g291(n569 ,n445 ,n446);
    nor g292(n494 ,n471 ,n492);
    nor g293(n464 ,n429 ,n462);
    not g294(n196 ,n5[5]);
    nor g295(n303 ,n126 ,n282);
    nor g296(n443 ,n421 ,n441);
    nor g297(n337 ,n13[15] ,n322);
    dff g298(.RN(n558), .SN(1'b1), .CK(n0), .D(n575), .Q(n14[7]));
    xnor g299(n4[14] ,n384 ,n6[14]);
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n369), .Q(n12[2]));
    nor g301(n493 ,n14[6] ,n491);
    xnor g302(n4[3] ,n384 ,n6[3]);
    nor g303(n306 ,n274 ,n304);
    not g304(n459 ,n458);
    not g305(n66 ,n10[4]);
    nor g306(n454 ,n7[9] ,n452);
    not g307(n132 ,n5[6]);
    not g308(n417 ,n7[4]);
    nor g309(n442 ,n7[5] ,n440);
    nor g310(n62 ,n39 ,n60);
    not g311(n492 ,n491);
    not g312(n495 ,n7[0]);
    nor g313(n394 ,n87 ,n88);
    or g314(n359 ,n324 ,n343);
    or g315(n355 ,n319 ,n339);
    not g316(n256 ,n257);
    not g317(n149 ,n396);
    not g318(n64 ,n10[13]);
    nor g319(n409 ,n58 ,n59);
    nor g320(n399 ,n102 ,n103);
    nor g321(n326 ,n138 ,n307);
    nor g322(n274 ,n175 ,n256);
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n358), .Q(n6[10]));
    not g324(n89 ,n88);
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n251), .Q(n10[10]));
    nor g326(n219 ,n179 ,n126);
    nor g327(n245 ,n166 ,n209);
    buf g328(n4[29], n4[31]);
    nor g329(n47 ,n43 ,n40);
    not g330(n197 ,n9[7]);
    not g331(n110 ,n109);
    not g332(n167 ,n412);
    or g333(n556 ,n551 ,n555);
    or g334(n555 ,n553 ,n552);
    not g335(n546 ,n14[4]);
    or g336(n33 ,n8[6] ,n8[5]);
    not g337(n107 ,n106);
    nor g338(n567 ,n451 ,n452);
    or g339(n526 ,n558 ,n7[1]);
    nor g340(n258 ,n389 ,n211);
    not g341(n389 ,n414);
    not g342(n192 ,n8[5]);
    or g343(n552 ,n549 ,n545);
    nor g344(n84 ,n10[3] ,n82);
    nor g345(n298 ,n126 ,n289);
    xor g346(n407 ,n8[7] ,n62);
    or g347(n25 ,n24 ,n23);
    nor g348(n234 ,n10[0] ,n209);
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n247), .Q(n10[5]));
    nor g350(n490 ,n14[5] ,n488);
    or g351(n534 ,n558 ,n502);
    nor g352(n329 ,n135 ,n307);
    not g353(n504 ,n7[1]);
    nor g354(n208 ,n190 ,n126);
    nor g355(n408 ,n61 ,n62);
    not g356(n184 ,n8[1]);
    not g357(n174 ,n12[2]);
    dff g358(.RN(n527), .SN(n542), .CK(n0), .D(n7[0]), .Q(n13[0]));
    not g359(n498 ,n7[12]);
    or g360(n415 ,n372 ,n382);
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n355), .Q(n6[13]));
    not g362(n182 ,n8[6]);
    not g363(n503 ,n7[6]);
    dff g364(.RN(n526), .SN(n541), .CK(n0), .D(n574), .Q(n13[1]));
    not g365(n168 ,n411);
    not g366(n75 ,n10[10]);
    not g367(n550 ,n14[5]);
    nor g368(n321 ,n126 ,n306);
    not g369(n162 ,n409);
    nor g370(n439 ,n7[4] ,n437);
    dff g371(.RN(n558), .SN(1'b1), .CK(n0), .D(n581), .Q(n14[1]));
    not g372(n116 ,n115);
    not g373(n83 ,n82);
    nor g374(n109 ,n73 ,n107);
    or g375(n19 ,n10[9] ,n10[8]);
    not g376(n444 ,n443);
    not g377(n183 ,n5[1]);
    dff g378(.RN(n524), .SN(n540), .CK(n0), .D(n572), .Q(n13[3]));
    nor g379(n563 ,n463 ,n464);
    or g380(n512 ,n558 ,n7[12]);
    nor g381(n467 ,n419 ,n465);
    buf g382(n4[16], n4[31]);
    nor g383(n351 ,n13[1] ,n322);
    not g384(n193 ,n9[5]);
    nor g385(n449 ,n428 ,n447);
    nor g386(n235 ,n9[0] ,n211);
    nor g387(n397 ,n96 ,n97);
    or g388(n375 ,n387 ,n5[6]);
    nor g389(n99 ,n10[8] ,n97);
    nor g390(n301 ,n261 ,n283);
    not g391(n45 ,n8[2]);
    nor g392(n319 ,n129 ,n307);
    nor g393(n413 ,n47 ,n46);
    xnor g394(n7[2] ,n2[2] ,n121);
    nor g395(n401 ,n108 ,n109);
    nor g396(n27 ,n20 ,n26);
    nor g397(n249 ,n150 ,n209);
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n294), .Q(n8[7]));
    not g399(n453 ,n452);
    buf g400(n4[22], n4[31]);
    or g401(n517 ,n558 ,n7[9]);
    not g402(n41 ,n8[4]);
    dff g403(.RN(n558), .SN(1'b1), .CK(n0), .D(n578), .Q(n14[4]));
    nor g404(n102 ,n10[9] ,n100);
    or g405(n367 ,n331 ,n350);
    not g406(n31 ,n8[0]);
    not g407(n191 ,n8[2]);
    nor g408(n204 ,n181 ,n126);
    nor g409(n224 ,n187 ,n126);
    not g410(n160 ,n407);
    nor g411(n277 ,n162 ,n256);
    or g412(n540 ,n558 ,n505);
    or g413(n200 ,n179 ,n9[0]);
    nor g414(n271 ,n186 ,n257);
    or g415(n17 ,n10[1] ,n10[0]);
    nor g416(n97 ,n70 ,n95);
    dff g417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n243), .Q(n10[3]));
    nor g418(n285 ,n279 ,n275);
    not g419(n128 ,n3[0]);
    dff g420(.RN(n518), .SN(n535), .CK(n0), .D(n567), .Q(n13[8]));
    nor g421(n314 ,n131 ,n307);
    nor g422(n431 ,n7[1] ,n559);
    or g423(n368 ,n316 ,n352);
    nor g424(n257 ,n174 ,n213);
    or g425(n214 ,n173 ,n12[1]);
    xnor g426(n4[12] ,n384 ,n6[12]);
    not g427(n465 ,n464);
    nor g428(n339 ,n13[13] ,n322);
    or g429(n514 ,n558 ,n7[13]);
    nor g430(n90 ,n10[5] ,n88);
    not g431(n165 ,n403);
    nor g432(n458 ,n427 ,n456);
    or g433(n236 ,n12[2] ,n211);
    nor g434(n331 ,n134 ,n307);
    xnor g435(n121 ,n2[18] ,n3[2]);
    nor g436(n343 ,n13[9] ,n322);
    not g437(n175 ,n11[0]);
    or g438(n202 ,n193 ,n9[4]);
    not g439(n438 ,n437);
    xor g440(n7[14] ,n2[30] ,n2[14]);
    nor g441(n346 ,n13[6] ,n322);
    not g442(n166 ,n397);
    nor g443(n579 ,n484 ,n485);
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n371), .Q(n6[5]));
    or g445(n414 ,n21 ,n29);
    nor g446(n345 ,n13[7] ,n322);
    not g447(n39 ,n8[6]);
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n363), .Q(n12[0]));
    nor g449(n290 ,n238 ,n264);
    or g450(n238 ,n202 ,n199);
    nor g451(n311 ,n215 ,n309);
    nor g452(n212 ,n12[0] ,n12[1]);
    dff g453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n298), .Q(n8[3]));
    not g454(n480 ,n479);
    nor g455(n275 ,n160 ,n256);
    not g456(n134 ,n13[2]);
    xnor g457(n7[5] ,n2[21] ,n124);
    not g458(n433 ,n432);
    or g459(n542 ,n558 ,n495);
    or g460(n516 ,n558 ,n7[10]);
    nor g461(n93 ,n10[6] ,n91);
    not g462(n65 ,n10[3]);
    buf g463(n4[17], n4[31]);
    xor g464(n405 ,n10[15] ,n118);
    not g465(n185 ,n5[0]);
    xnor g466(n125 ,n2[6] ,n3[6]);
    nor g467(n369 ,n126 ,n335);
    nor g468(n363 ,n126 ,n336);
    nor g469(n226 ,n126 ,n127);
    nor g470(n488 ,n473 ,n486);
    nor g471(n210 ,n173 ,n172);
    not g472(n54 ,n53);
    nor g473(n392 ,n81 ,n82);
    not g474(n173 ,n12[0]);
    nor g475(n227 ,n132 ,n126);
    nor g476(n229 ,n178 ,n126);
    nor g477(n451 ,n7[8] ,n449);
    nor g478(n248 ,n157 ,n209);
    buf g479(n4[21], n4[31]);
    or g480(n521 ,n558 ,n7[7]);
    or g481(n373 ,n390 ,n5[0]);
    or g482(n554 ,n548 ,n550);
    nor g483(n349 ,n13[3] ,n322);
    nor g484(n268 ,n182 ,n257);
    not g485(n322 ,n321);
    xnor g486(n7[4] ,n2[20] ,n122);
    not g487(n156 ,n400);
    nor g488(n393 ,n84 ,n85);
    nor g489(n96 ,n10[7] ,n94);
    xnor g490(n4[0] ,n384 ,n6[0]);
    not g491(n151 ,n404);
    or g492(n380 ,n375 ,n379);
    nor g493(n250 ,n170 ,n209);
    nor g494(n576 ,n493 ,n494);
    not g495(n213 ,n212);
    not g496(n43 ,n8[1]);
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n223), .Q(n9[1]));
    not g498(n462 ,n461);
    nor g499(n56 ,n41 ,n54);
    not g500(n164 ,n395);
    not g501(n139 ,n13[1]);
    xnor g502(n4[4] ,n384 ,n6[4]);
    nor g503(n295 ,n126 ,n286);
    or g504(n209 ,n126 ,n128);
    not g505(n126 ,n1);
    buf g506(n4[20], n4[31]);
    not g507(n69 ,n10[8]);
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n234), .Q(n10[0]));
    not g509(n547 ,n14[3]);
    nor g510(n117 ,n10[14] ,n115);
    nor g511(n252 ,n148 ,n209);
    not g512(n450 ,n449);
    not g513(n159 ,n405);
    nor g514(n79 ,n71 ,n76);
    or g515(n230 ,n195 ,n172);
    nor g516(n452 ,n426 ,n450);
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n248), .Q(n10[4]));
    not g518(n386 ,n5[5]);
    or g519(n528 ,n558 ,n511);
    or g520(n379 ,n373 ,n374);
    or g521(n16 ,n10[5] ,n10[4]);
    or g522(n20 ,n10[3] ,n10[2]);
    not g523(n474 ,n14[3]);
    not g524(n189 ,n5[2]);
    xnor g525(n119 ,n2[3] ,n3[3]);
    buf g526(n4[26], n4[31]);
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n208), .Q(n9[4]));
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n353), .Q(n6[15]));
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n240), .Q(n10[14]));
    not g530(n436 ,n435);
    nor g531(n267 ,n192 ,n257);
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n252), .Q(n10[9]));
    not g533(n72 ,n10[9]);
    nor g534(n279 ,n194 ,n257);
    dff g535(.RN(n513), .SN(n529), .CK(n0), .D(n561), .Q(n13[14]));
    not g536(n468 ,n467);
    nor g537(n78 ,n10[1] ,n10[0]);
    or g538(n518 ,n558 ,n7[8]);
    or g539(n358 ,n332 ,n342);
    not g540(n180 ,n11[1]);
    nor g541(n469 ,n7[14] ,n467);
    dff g542(.RN(n558), .SN(1'b1), .CK(n0), .D(n579), .Q(n14[3]));
    nor g543(n566 ,n454 ,n455);
    nor g544(n309 ,n302 ,n305);
    xnor g545(n4[6] ,n384 ,n6[6]);
    not g546(n477 ,n14[2]);
    nor g547(n396 ,n93 ,n94);
    not g548(n158 ,n393);
    nor g549(n205 ,n193 ,n126);
    buf g550(n4[30], n4[31]);
    not g551(n153 ,n413);
    nor g552(n578 ,n487 ,n488);
    or g553(n515 ,n558 ,n7[11]);
    not g554(n129 ,n13[13]);
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n227), .Q(n5[7]));
    nor g556(n344 ,n13[8] ,n322);
    dff g557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n364), .Q(n6[4]));
    nor g558(n335 ,n320 ,n312);
    not g559(n135 ,n13[4]);
    nor g560(n336 ,n315 ,n311);
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n228), .Q(n5[6]));
    nor g562(n28 ,n15 ,n27);
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n361), .Q(n6[7]));
    nor g564(n287 ,n267 ,n277);
    not g565(n497 ,n7[14]);
    or g566(n525 ,n558 ,n7[2]);
    or g567(n536 ,n558 ,n500);
    not g568(n548 ,n14[6]);
    or g569(n532 ,n558 ,n496);
    not g570(n80 ,n79);
    nor g571(n478 ,n14[1] ,n14[0]);
    buf g572(n4[27], n4[31]);
    not g573(n32 ,n8[3]);
    not g574(n424 ,n7[3]);
    or g575(n520 ,n558 ,n7[6]);
    dff g576(.RN(n515), .SN(n532), .CK(n0), .D(n564), .Q(n13[11]));
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n365), .Q(n6[3]));
    not g578(n508 ,n7[10]);
    or g579(n23 ,n18 ,n16);
    or g580(n215 ,n12[0] ,n12[2]);
    xnor g581(n7[3] ,n119 ,n2[19]);
    nor g582(n112 ,n77 ,n110);
    or g583(n263 ,n210 ,n233);
    nor g584(n241 ,n165 ,n209);
    nor g585(n206 ,n126 ,n128);
    or g586(n366 ,n328 ,n351);
    xor g587(n7[10] ,n2[26] ,n2[10]);
    nor g588(n88 ,n66 ,n86);
    or g589(n261 ,n235 ,n255);
    not g590(n483 ,n482);
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n201), .Q(n5[1]));
    or g592(n531 ,n558 ,n498);
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n207), .Q(n9[5]));
    nor g594(n58 ,n8[5] ,n56);
    xnor g595(n4[7] ,n384 ,n6[7]);
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n368), .Q(n6[0]));
    nor g597(n61 ,n8[6] ,n59);
    not g598(n63 ,n10[6]);
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n366), .Q(n6[1]));
    or g600(n233 ,n12[2] ,n212);
    not g601(n146 ,n13[10]);
    xnor g602(n282 ,n257 ,n8[0]);
    or g603(n354 ,n318 ,n338);
    or g604(n26 ,n17 ,n25);
    dff g605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n218), .Q(n11[2]));
    not g606(n144 ,n9[4]);
    not g607(n505 ,n7[3]);
    or g608(n22 ,n10[11] ,n10[10]);
    dff g609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n370), .Q(n12[1]));
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n367), .Q(n6[2]));
    xor g611(n7[12] ,n2[28] ,n2[12]);
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n244), .Q(n10[8]));
    nor g613(n246 ,n149 ,n209);
    xor g614(n575 ,n14[7] ,n494);
    not g615(n430 ,n7[1]);
    not g616(n475 ,n14[1]);
    dff g617(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n360), .Q(n6[8]));
    dff g618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n299), .Q(n8[2]));
    nor g619(n105 ,n10[10] ,n103);
    nor g620(n218 ,n180 ,n126);
    nor g621(n49 ,n8[2] ,n47);
    nor g622(n482 ,n477 ,n480);
    not g623(n98 ,n97);
    not g624(n44 ,n8[5]);
    not g625(n147 ,n13[6]);
    not g626(n551 ,n14[7]);
    or g627(n523 ,n558 ,n7[4]);
    not g628(n421 ,n7[5]);
    dff g629(.RN(n512), .SN(n531), .CK(n0), .D(n563), .Q(n13[12]));
    not g630(n419 ,n7[13]);
    or g631(n357 ,n323 ,n341);
    not g632(n148 ,n399);
    xnor g633(n7[7] ,n2[23] ,n123);
    not g634(n142 ,n13[14]);
    nor g635(n313 ,n172 ,n308);
    nor g636(n404 ,n117 ,n118);
    not g637(n71 ,n10[1]);
    not g638(n499 ,n7[4]);
    or g639(n533 ,n558 ,n508);
    nor g640(n448 ,n7[7] ,n446);
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n359), .Q(n6[9]));
    nor g642(n244 ,n171 ,n209);
    not g643(n163 ,n402);
    or g644(n356 ,n314 ,n340);
    nor g645(n328 ,n139 ,n307);
    nor g646(n94 ,n63 ,n92);
    nor g647(n232 ,n188 ,n126);
    or g648(n538 ,n558 ,n507);
    not g649(n157 ,n394);
    not g650(n137 ,n13[8]);
    not g651(n177 ,n10[0]);
    nor g652(n288 ,n271 ,n278);
    nor g653(n317 ,n133 ,n307);
    nor g654(n85 ,n65 ,n83);
    nor g655(n461 ,n420 ,n459);
    nor g656(n297 ,n126 ,n288);
    not g657(n423 ,n7[14]);
    not g658(n194 ,n8[7]);
    not g659(n447 ,n446);
    not g660(n190 ,n9[3]);
    nor g661(n400 ,n105 ,n106);
    nor g662(n332 ,n146 ,n307);
    nor g663(n455 ,n422 ,n453);
    or g664(n530 ,n558 ,n501);
    nor g665(n276 ,n155 ,n256);
    not g666(n42 ,n8[3]);
    dff g667(.RN(n523), .SN(n539), .CK(n0), .D(n571), .Q(n13[4]));
    or g668(n372 ,n385 ,n5[2]);
    nor g669(n561 ,n469 ,n470);
    not g670(n133 ,n13[15]);
    not g671(n15 ,n10[12]);
    or g672(n374 ,n386 ,n5[4]);
    or g673(n524 ,n558 ,n7[3]);
    not g674(n76 ,n10[0]);
    nor g675(n348 ,n13[4] ,n322);
    nor g676(n103 ,n72 ,n101);
    nor g677(n391 ,n79 ,n78);
    nor g678(n318 ,n142 ,n307);
    not g679(n77 ,n10[12]);
    not g680(n169 ,n11[3]);
    not g681(n186 ,n8[4]);
    nor g682(n270 ,n168 ,n256);
    xnor g683(n4[1] ,n384 ,n6[1]);
    nor g684(n300 ,n126 ,n291);
    nor g685(n231 ,n177 ,n172);
    nor g686(n222 ,n183 ,n126);
    nor g687(n333 ,n136 ,n307);
    dff g688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n224), .Q(n5[5]));
    nor g689(n273 ,n184 ,n257);
    xnor g690(n4[31] ,n6[16] ,n384);
    not g691(n154 ,n410);
    xor g692(n572 ,n7[3] ,n435);
    nor g693(n437 ,n424 ,n436);
    or g694(n237 ,n200 ,n198);
    nor g695(n203 ,n195 ,n126);
    or g696(n259 ,n180 ,n230);
    or g697(n353 ,n317 ,n337);
    or g698(n406 ,n33 ,n38);
    nor g699(n108 ,n10[11] ,n106);
    nor g700(n484 ,n14[3] ,n482);
    nor g701(n228 ,n196 ,n126);
    dff g702(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n9[0]));
endmodule
