module top(n0, n1, n3, n5, n6, n7, n4, n2, n8, n9, n10, n11, n12, n14, n13);
    input n0, n1, n2;
    input [1:0] n3, n4;
    input [15:0] n5;
    input [31:0] n6;
    input [3:0] n7;
    output [31:0] n8;
    output n9, n10;
    output [3:0] n11;
    output [7:0] n12, n13;
    output [15:0] n14;
    wire n0, n1, n2;
    wire [1:0] n3, n4;
    wire [15:0] n5;
    wire [31:0] n6;
    wire [3:0] n7;
    wire [31:0] n8;
    wire n9, n10;
    wire [3:0] n11;
    wire [7:0] n12, n13;
    wire [15:0] n14;
    wire [3:0] n15;
    wire [2:0] n16;
    wire [15:0] n17;
    wire [3:0] n18;
    wire [1:0] n19;
    wire [31:0] n20;
    wire n21, n22, n23, n24, n25, n26, n27, n28;
    wire n29, n30, n31, n32, n33, n34, n35, n36;
    wire n37, n38, n39, n40, n41, n42, n43, n44;
    wire n45, n46, n47, n48, n49, n50, n51, n52;
    wire n53, n54, n55, n56, n57, n58, n59, n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591;
    buf g0(n13[0], 1'b0);
    buf g1(n13[1], 1'b0);
    buf g2(n12[0], 1'b0);
    buf g3(n12[1], 1'b0);
    buf g4(n12[2], 1'b0);
    buf g5(n12[3], 1'b0);
    buf g6(n12[4], 1'b0);
    buf g7(n12[5], 1'b0);
    buf g8(n12[6], 1'b0);
    buf g9(n12[7], 1'b0);
    buf g10(n8[20], 1'b0);
    buf g11(n8[21], 1'b0);
    buf g12(n8[22], 1'b0);
    buf g13(n8[23], 1'b0);
    buf g14(n8[24], 1'b0);
    buf g15(n8[25], 1'b0);
    buf g16(n8[26], 1'b0);
    buf g17(n8[27], 1'b0);
    buf g18(n8[28], 1'b0);
    buf g19(n8[29], 1'b0);
    buf g20(n8[30], 1'b0);
    buf g21(n8[31], 1'b0);
    not g22(n563 ,n591);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n562), .Q(n15[2]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n561), .Q(n15[0]));
    or g25(n562 ,n546 ,n559);
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n560), .Q(n15[1]));
    or g27(n561 ,n548 ,n556);
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n555), .Q(n16[1]));
    or g29(n560 ,n547 ,n557);
    or g30(n559 ,n425 ,n558);
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n552), .Q(n11[3]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n551), .Q(n11[2]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n553), .Q(n11[0]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n550), .Q(n11[1]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n544), .Q(n16[0]));
    nor g36(n558 ,n173 ,n554);
    nor g37(n557 ,n158 ,n554);
    nor g38(n556 ,n15[0] ,n554);
    or g39(n555 ,n511 ,n545);
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n549), .Q(n16[2]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n517), .Q(n8[14]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n531), .Q(n8[0]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n530), .Q(n8[1]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n529), .Q(n8[2]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n542), .Q(n8[3]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n527), .Q(n8[4]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n526), .Q(n8[5]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n525), .Q(n8[6]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n524), .Q(n8[7]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n523), .Q(n8[8]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n522), .Q(n8[9]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n521), .Q(n8[10]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n520), .Q(n8[11]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n519), .Q(n8[12]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n518), .Q(n8[13]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n535), .Q(n8[19]));
    or g57(n553 ,n421 ,n541);
    or g58(n552 ,n418 ,n539);
    or g59(n551 ,n419 ,n540);
    or g60(n550 ,n420 ,n528);
    or g61(n549 ,n465 ,n532);
    nor g62(n548 ,n193 ,n543);
    nor g63(n547 ,n201 ,n543);
    nor g64(n546 ,n199 ,n543);
    or g65(n545 ,n415 ,n533);
    or g66(n544 ,n411 ,n534);
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n514), .Q(n8[17]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n536), .Q(n8[18]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n537), .Q(n9));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n516), .Q(n8[15]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n515), .Q(n8[16]));
    or g72(n554 ,n121 ,n538);
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n458), .Q(n17[9]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n464), .Q(n17[10]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n463), .Q(n17[11]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n462), .Q(n17[12]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n461), .Q(n17[13]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n460), .Q(n17[14]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n457), .Q(n17[15]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n431), .Q(n17[3]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n430), .Q(n17[4]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n17[1]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n432), .Q(n14[15]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n435), .Q(n17[2]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n451), .Q(n14[1]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n450), .Q(n14[2]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n449), .Q(n14[3]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n448), .Q(n14[4]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n439), .Q(n17[0]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n446), .Q(n14[5]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n445), .Q(n14[6]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n444), .Q(n14[7]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n443), .Q(n14[8]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n14[9]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n440), .Q(n14[10]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n438), .Q(n14[11]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n436), .Q(n14[12]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n434), .Q(n14[13]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n433), .Q(n14[14]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n452), .Q(n14[0]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n454), .Q(n18[2]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n442), .Q(n19[1]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n453), .Q(n18[3]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n456), .Q(n18[0]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n455), .Q(n18[1]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n447), .Q(n19[0]));
    or g107(n542 ,n483 ,n504);
    nor g108(n541 ,n256 ,n469);
    nor g109(n540 ,n256 ,n512);
    nor g110(n539 ,n265 ,n512);
    nor g111(n537 ,n126 ,n468);
    or g112(n536 ,n510 ,n500);
    or g113(n535 ,n488 ,n508);
    or g114(n534 ,n417 ,n467);
    or g115(n533 ,n287 ,n513);
    or g116(n532 ,n513 ,n466);
    or g117(n531 ,n486 ,n507);
    or g118(n530 ,n485 ,n506);
    or g119(n529 ,n484 ,n505);
    nor g120(n528 ,n265 ,n469);
    or g121(n527 ,n482 ,n503);
    or g122(n526 ,n481 ,n502);
    or g123(n525 ,n480 ,n501);
    or g124(n524 ,n487 ,n499);
    or g125(n523 ,n479 ,n498);
    or g126(n522 ,n478 ,n497);
    or g127(n521 ,n477 ,n496);
    or g128(n520 ,n476 ,n495);
    or g129(n519 ,n475 ,n493);
    or g130(n518 ,n474 ,n492);
    or g131(n517 ,n473 ,n491);
    or g132(n516 ,n472 ,n490);
    or g133(n515 ,n471 ,n489);
    or g134(n514 ,n509 ,n494);
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n428), .Q(n17[6]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n459), .Q(n17[7]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n427), .Q(n17[8]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n429), .Q(n17[5]));
    or g139(n543 ,n121 ,n470);
    nor g140(n511 ,n191 ,n424);
    nor g141(n510 ,n207 ,n423);
    nor g142(n509 ,n131 ,n423);
    nor g143(n508 ,n237 ,n422);
    nor g144(n507 ,n194 ,n422);
    nor g145(n506 ,n197 ,n422);
    nor g146(n505 ,n198 ,n422);
    nor g147(n504 ,n196 ,n422);
    nor g148(n503 ,n234 ,n422);
    nor g149(n502 ,n238 ,n422);
    nor g150(n501 ,n223 ,n422);
    nor g151(n500 ,n205 ,n422);
    nor g152(n499 ,n217 ,n422);
    nor g153(n498 ,n224 ,n422);
    nor g154(n497 ,n139 ,n422);
    nor g155(n496 ,n226 ,n422);
    nor g156(n495 ,n218 ,n422);
    nor g157(n494 ,n216 ,n422);
    nor g158(n493 ,n245 ,n422);
    nor g159(n492 ,n243 ,n422);
    nor g160(n491 ,n134 ,n422);
    nor g161(n490 ,n222 ,n422);
    nor g162(n489 ,n233 ,n422);
    nor g163(n488 ,n219 ,n423);
    nor g164(n487 ,n231 ,n423);
    nor g165(n486 ,n212 ,n423);
    nor g166(n485 ,n232 ,n423);
    nor g167(n484 ,n242 ,n423);
    nor g168(n483 ,n211 ,n423);
    nor g169(n482 ,n140 ,n423);
    nor g170(n481 ,n138 ,n423);
    nor g171(n480 ,n225 ,n423);
    nor g172(n479 ,n236 ,n423);
    nor g173(n478 ,n213 ,n423);
    nor g174(n477 ,n229 ,n423);
    nor g175(n476 ,n214 ,n423);
    nor g176(n475 ,n209 ,n423);
    nor g177(n474 ,n137 ,n423);
    nor g178(n473 ,n133 ,n423);
    nor g179(n472 ,n208 ,n423);
    nor g180(n471 ,n240 ,n423);
    nor g181(n513 ,n136 ,n409);
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n396), .Q(n10));
    or g183(n512 ,n197 ,n426);
    nor g184(n468 ,n416 ,n407);
    nor g185(n467 ,n190 ,n424);
    nor g186(n466 ,n127 ,n424);
    nor g187(n465 ,n254 ,n408);
    nor g188(n464 ,n125 ,n405);
    nor g189(n463 ,n125 ,n404);
    nor g190(n462 ,n125 ,n403);
    nor g191(n461 ,n122 ,n402);
    nor g192(n460 ,n123 ,n401);
    nor g193(n459 ,n125 ,n372);
    nor g194(n458 ,n123 ,n406);
    nor g195(n457 ,n122 ,n400);
    nor g196(n456 ,n126 ,n399);
    nor g197(n455 ,n122 ,n410);
    nor g198(n454 ,n125 ,n412);
    nor g199(n453 ,n126 ,n413);
    nor g200(n452 ,n122 ,n398);
    nor g201(n451 ,n124 ,n397);
    nor g202(n450 ,n124 ,n395);
    nor g203(n449 ,n126 ,n394);
    nor g204(n448 ,n124 ,n392);
    nor g205(n447 ,n122 ,n391);
    nor g206(n446 ,n126 ,n390);
    nor g207(n445 ,n123 ,n388);
    nor g208(n444 ,n123 ,n387);
    nor g209(n443 ,n124 ,n386);
    nor g210(n442 ,n122 ,n389);
    nor g211(n441 ,n124 ,n385);
    nor g212(n440 ,n124 ,n383);
    nor g213(n439 ,n126 ,n384);
    nor g214(n438 ,n125 ,n382);
    nor g215(n437 ,n124 ,n379);
    nor g216(n436 ,n122 ,n381);
    nor g217(n435 ,n126 ,n377);
    nor g218(n434 ,n125 ,n380);
    nor g219(n433 ,n123 ,n378);
    nor g220(n432 ,n123 ,n376);
    nor g221(n431 ,n124 ,n375);
    nor g222(n430 ,n126 ,n374);
    nor g223(n429 ,n123 ,n371);
    nor g224(n428 ,n123 ,n393);
    nor g225(n427 ,n122 ,n373);
    nor g226(n470 ,n251 ,n414);
    or g227(n469 ,n18[1] ,n426);
    not g228(n422 ,n423);
    nor g229(n421 ,n200 ,n329);
    nor g230(n420 ,n128 ,n329);
    nor g231(n419 ,n239 ,n329);
    nor g232(n418 ,n220 ,n329);
    nor g233(n417 ,n132 ,n333);
    nor g234(n416 ,n129 ,n331);
    nor g235(n415 ,n255 ,n330);
    nor g236(n413 ,n313 ,n341);
    nor g237(n412 ,n314 ,n342);
    nor g238(n411 ,n19[0] ,n330);
    nor g239(n410 ,n315 ,n343);
    or g240(n409 ,n2 ,n333);
    or g241(n408 ,n259 ,n330);
    nor g242(n407 ,n251 ,n332);
    nor g243(n406 ,n327 ,n353);
    nor g244(n405 ,n311 ,n350);
    nor g245(n404 ,n324 ,n349);
    nor g246(n403 ,n323 ,n348);
    nor g247(n402 ,n322 ,n347);
    nor g248(n401 ,n320 ,n346);
    nor g249(n400 ,n318 ,n345);
    nor g250(n399 ,n317 ,n344);
    or g251(n426 ,n18[2] ,n330);
    nor g252(n425 ,n277 ,n288);
    or g253(n424 ,n276 ,n286);
    nor g254(n423 ,n264 ,n332);
    xnor g255(n398 ,n14[0] ,n275);
    nor g256(n397 ,n309 ,n368);
    or g257(n396 ,n369 ,n290);
    nor g258(n395 ,n316 ,n367);
    nor g259(n394 ,n308 ,n366);
    nor g260(n393 ,n319 ,n352);
    nor g261(n392 ,n307 ,n354);
    nor g262(n391 ,n289 ,n338);
    nor g263(n390 ,n293 ,n365);
    nor g264(n389 ,n306 ,n337);
    nor g265(n388 ,n298 ,n364);
    nor g266(n387 ,n328 ,n363);
    nor g267(n386 ,n302 ,n362);
    nor g268(n385 ,n294 ,n361);
    nor g269(n384 ,n300 ,n339);
    nor g270(n383 ,n296 ,n360);
    nor g271(n382 ,n297 ,n359);
    nor g272(n381 ,n304 ,n358);
    nor g273(n380 ,n292 ,n357);
    nor g274(n379 ,n326 ,n336);
    nor g275(n378 ,n295 ,n355);
    nor g276(n377 ,n299 ,n335);
    nor g277(n376 ,n303 ,n370);
    nor g278(n375 ,n312 ,n351);
    nor g279(n374 ,n291 ,n356);
    nor g280(n373 ,n321 ,n334);
    nor g281(n372 ,n325 ,n340);
    nor g282(n371 ,n301 ,n305);
    nor g283(n370 ,n188 ,n274);
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n284), .Q(n20[1]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n281), .Q(n20[2]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n20[3]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n270), .Q(n20[4]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n266), .Q(n20[5]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n285), .Q(n20[6]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n283), .Q(n20[7]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n271), .Q(n20[8]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n282), .Q(n20[9]));
    nor g293(n369 ,n221 ,n277);
    nor g294(n368 ,n182 ,n274);
    nor g295(n367 ,n180 ,n274);
    nor g296(n366 ,n174 ,n274);
    nor g297(n365 ,n171 ,n274);
    nor g298(n364 ,n142 ,n274);
    nor g299(n363 ,n156 ,n274);
    nor g300(n362 ,n185 ,n274);
    nor g301(n361 ,n159 ,n274);
    nor g302(n360 ,n165 ,n274);
    nor g303(n359 ,n179 ,n274);
    nor g304(n358 ,n170 ,n274);
    nor g305(n357 ,n175 ,n274);
    nor g306(n356 ,n160 ,n272);
    nor g307(n355 ,n164 ,n274);
    nor g308(n354 ,n176 ,n274);
    nor g309(n353 ,n146 ,n272);
    nor g310(n352 ,n166 ,n272);
    nor g311(n351 ,n162 ,n272);
    nor g312(n350 ,n172 ,n272);
    nor g313(n349 ,n151 ,n272);
    nor g314(n348 ,n145 ,n272);
    nor g315(n347 ,n144 ,n272);
    nor g316(n346 ,n189 ,n272);
    nor g317(n345 ,n154 ,n272);
    nor g318(n344 ,n186 ,n272);
    nor g319(n343 ,n177 ,n272);
    nor g320(n342 ,n163 ,n272);
    nor g321(n341 ,n181 ,n272);
    nor g322(n340 ,n155 ,n272);
    nor g323(n339 ,n152 ,n272);
    nor g324(n338 ,n184 ,n272);
    nor g325(n337 ,n187 ,n272);
    nor g326(n336 ,n153 ,n272);
    nor g327(n335 ,n157 ,n272);
    nor g328(n334 ,n161 ,n272);
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n267), .Q(n20[0]));
    not g330(n332 ,n331);
    nor g331(n328 ,n135 ,n275);
    nor g332(n327 ,n243 ,n273);
    nor g333(n326 ,n238 ,n273);
    nor g334(n325 ,n218 ,n273);
    nor g335(n324 ,n222 ,n273);
    nor g336(n323 ,n233 ,n273);
    nor g337(n322 ,n216 ,n273);
    nor g338(n321 ,n245 ,n273);
    nor g339(n320 ,n205 ,n273);
    nor g340(n319 ,n226 ,n273);
    nor g341(n318 ,n237 ,n273);
    nor g342(n317 ,n194 ,n273);
    nor g343(n316 ,n203 ,n275);
    nor g344(n315 ,n197 ,n273);
    nor g345(n314 ,n198 ,n273);
    nor g346(n313 ,n196 ,n273);
    nor g347(n312 ,n217 ,n273);
    nor g348(n311 ,n134 ,n273);
    nor g349(n310 ,n563 ,n276);
    nor g350(n309 ,n228 ,n275);
    nor g351(n308 ,n206 ,n275);
    nor g352(n307 ,n227 ,n275);
    nor g353(n306 ,n195 ,n273);
    nor g354(n305 ,n143 ,n272);
    nor g355(n304 ,n215 ,n275);
    nor g356(n303 ,n230 ,n275);
    nor g357(n302 ,n244 ,n275);
    nor g358(n301 ,n139 ,n273);
    nor g359(n300 ,n234 ,n273);
    nor g360(n299 ,n223 ,n273);
    nor g361(n298 ,n241 ,n275);
    nor g362(n297 ,n202 ,n275);
    nor g363(n296 ,n141 ,n275);
    nor g364(n295 ,n235 ,n275);
    nor g365(n294 ,n210 ,n275);
    nor g366(n293 ,n204 ,n275);
    nor g367(n292 ,n130 ,n275);
    nor g368(n291 ,n224 ,n273);
    nor g369(n290 ,n190 ,n280);
    nor g370(n289 ,n192 ,n273);
    or g371(n288 ,n250 ,n279);
    nor g372(n287 ,n125 ,n272);
    or g373(n286 ,n277 ,n278);
    or g374(n333 ,n16[0] ,n280);
    nor g375(n331 ,n249 ,n276);
    or g376(n330 ,n121 ,n274);
    or g377(n329 ,n121 ,n268);
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n257), .Q(n13[7]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n262), .Q(n13[3]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n258), .Q(n13[4]));
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n261), .Q(n13[5]));
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n263), .Q(n13[6]));
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n260), .Q(n13[2]));
    nor g384(n285 ,n149 ,n248);
    nor g385(n284 ,n169 ,n248);
    nor g386(n283 ,n183 ,n248);
    nor g387(n282 ,n167 ,n248);
    nor g388(n281 ,n150 ,n248);
    not g389(n279 ,n278);
    not g390(n274 ,n275);
    not g391(n272 ,n273);
    nor g392(n271 ,n147 ,n248);
    nor g393(n270 ,n168 ,n248);
    nor g394(n269 ,n148 ,n248);
    nor g395(n268 ,n127 ,n253);
    nor g396(n267 ,n20[0] ,n248);
    nor g397(n266 ,n178 ,n248);
    or g398(n280 ,n121 ,n252);
    nor g399(n278 ,n15[1] ,n246);
    or g400(n277 ,n121 ,n251);
    nor g401(n276 ,n191 ,n247);
    nor g402(n275 ,n16[2] ,n253);
    nor g403(n273 ,n16[2] ,n250);
    not g404(n264 ,n263);
    nor g405(n262 ,n128 ,n121);
    nor g406(n261 ,n195 ,n121);
    nor g407(n260 ,n200 ,n121);
    nor g408(n259 ,n192 ,n195);
    nor g409(n258 ,n192 ,n121);
    nor g410(n257 ,n191 ,n121);
    or g411(n265 ,n194 ,n18[3]);
    nor g412(n263 ,n190 ,n121);
    not g413(n255 ,n254);
    not g414(n252 ,n251);
    not g415(n250 ,n249);
    nor g416(n247 ,n190 ,n16[2]);
    or g417(n246 ,n15[0] ,n15[2]);
    or g418(n256 ,n18[0] ,n18[3]);
    nor g419(n254 ,n19[0] ,n19[1]);
    or g420(n253 ,n191 ,n16[0]);
    nor g421(n251 ,n16[1] ,n16[2]);
    nor g422(n249 ,n190 ,n16[1]);
    or g423(n248 ,n121 ,n575);
    not g424(n245 ,n17[8]);
    not g425(n244 ,n14[8]);
    not g426(n243 ,n17[9]);
    not g427(n242 ,n8[2]);
    not g428(n241 ,n14[6]);
    not g429(n240 ,n8[16]);
    not g430(n239 ,n11[2]);
    not g431(n238 ,n17[1]);
    not g432(n237 ,n17[15]);
    not g433(n236 ,n8[8]);
    not g434(n235 ,n14[14]);
    not g435(n234 ,n17[0]);
    not g436(n233 ,n17[12]);
    not g437(n232 ,n8[1]);
    not g438(n231 ,n8[7]);
    not g439(n230 ,n14[15]);
    not g440(n229 ,n8[10]);
    not g441(n228 ,n14[1]);
    not g442(n227 ,n14[4]);
    not g443(n226 ,n17[6]);
    not g444(n225 ,n8[6]);
    not g445(n224 ,n17[4]);
    not g446(n223 ,n17[2]);
    not g447(n222 ,n17[11]);
    not g448(n221 ,n10);
    not g449(n220 ,n11[3]);
    not g450(n219 ,n8[19]);
    not g451(n218 ,n17[7]);
    not g452(n217 ,n17[3]);
    not g453(n216 ,n17[13]);
    not g454(n215 ,n14[12]);
    not g455(n214 ,n8[11]);
    not g456(n213 ,n8[9]);
    not g457(n212 ,n8[0]);
    not g458(n211 ,n8[3]);
    not g459(n210 ,n14[9]);
    not g460(n209 ,n8[12]);
    not g461(n208 ,n8[15]);
    not g462(n207 ,n8[18]);
    not g463(n206 ,n14[3]);
    not g464(n205 ,n17[14]);
    not g465(n204 ,n14[5]);
    not g466(n203 ,n14[2]);
    not g467(n202 ,n14[11]);
    not g468(n201 ,n15[1]);
    not g469(n200 ,n11[0]);
    not g470(n199 ,n15[2]);
    not g471(n198 ,n18[2]);
    not g472(n197 ,n18[1]);
    not g473(n196 ,n18[3]);
    not g474(n195 ,n19[1]);
    not g475(n194 ,n18[0]);
    not g476(n193 ,n15[0]);
    not g477(n192 ,n19[0]);
    not g478(n191 ,n16[1]);
    not g479(n190 ,n16[0]);
    not g480(n189 ,n5[14]);
    not g481(n188 ,n576);
    not g482(n187 ,n3[1]);
    not g483(n186 ,n7[0]);
    not g484(n185 ,n583);
    not g485(n184 ,n3[0]);
    not g486(n183 ,n572);
    not g487(n182 ,n590);
    not g488(n181 ,n7[3]);
    not g489(n180 ,n589);
    not g490(n179 ,n580);
    not g491(n178 ,n570);
    not g492(n177 ,n7[1]);
    not g493(n176 ,n587);
    not g494(n175 ,n578);
    not g495(n174 ,n588);
    not g496(n173 ,n565);
    not g497(n172 ,n5[10]);
    not g498(n171 ,n586);
    not g499(n170 ,n579);
    not g500(n169 ,n566);
    not g501(n168 ,n569);
    not g502(n167 ,n574);
    not g503(n166 ,n5[6]);
    not g504(n165 ,n581);
    not g505(n164 ,n577);
    not g506(n163 ,n7[2]);
    not g507(n162 ,n5[3]);
    not g508(n161 ,n5[8]);
    not g509(n160 ,n5[4]);
    not g510(n159 ,n582);
    not g511(n158 ,n564);
    not g512(n157 ,n5[2]);
    not g513(n156 ,n584);
    not g514(n155 ,n5[7]);
    not g515(n154 ,n5[15]);
    not g516(n153 ,n5[1]);
    not g517(n152 ,n5[0]);
    not g518(n151 ,n5[11]);
    not g519(n150 ,n567);
    not g520(n149 ,n571);
    not g521(n148 ,n568);
    not g522(n147 ,n573);
    not g523(n146 ,n5[9]);
    not g524(n145 ,n5[12]);
    not g525(n144 ,n5[13]);
    not g526(n143 ,n5[5]);
    not g527(n142 ,n585);
    not g528(n141 ,n14[10]);
    not g529(n140 ,n8[4]);
    not g530(n139 ,n17[5]);
    not g531(n138 ,n8[5]);
    not g532(n137 ,n8[13]);
    not g533(n136 ,n575);
    not g534(n135 ,n14[7]);
    not g535(n134 ,n17[10]);
    not g536(n133 ,n8[14]);
    not g537(n132 ,n2);
    not g538(n131 ,n8[17]);
    not g539(n130 ,n14[13]);
    not g540(n129 ,n9);
    not g541(n128 ,n11[1]);
    not g542(n127 ,n16[2]);
    not g543(n126 ,n1);
    not g544(n125 ,n1);
    not g545(n124 ,n1);
    not g546(n123 ,n1);
    not g547(n122 ,n1);
    not g548(n121 ,n1);
    xor g549(n565 ,n15[2] ,n21);
    xnor g550(n564 ,n15[1] ,n15[0]);
    nor g551(n21 ,n15[1] ,n15[0]);
    or g552(n591 ,n15[0] ,n22);
    or g553(n22 ,n15[2] ,n15[1]);
    nor g554(n575 ,n29 ,n32);
    or g555(n32 ,n24 ,n31);
    or g556(n31 ,n30 ,n28);
    or g557(n30 ,n27 ,n23);
    or g558(n29 ,n25 ,n26);
    nor g559(n28 ,n20[4] ,n20[3]);
    not g560(n27 ,n20[9]);
    not g561(n26 ,n20[5]);
    not g562(n25 ,n20[6]);
    not g563(n24 ,n20[7]);
    not g564(n23 ,n20[8]);
    xor g565(n574 ,n20[9] ,n64);
    nor g566(n573 ,n63 ,n64);
    nor g567(n64 ,n39 ,n62);
    nor g568(n63 ,n20[8] ,n61);
    nor g569(n572 ,n60 ,n61);
    not g570(n62 ,n61);
    nor g571(n61 ,n35 ,n59);
    nor g572(n60 ,n20[7] ,n58);
    nor g573(n571 ,n57 ,n58);
    not g574(n59 ,n58);
    nor g575(n58 ,n36 ,n56);
    nor g576(n57 ,n20[6] ,n55);
    nor g577(n570 ,n54 ,n55);
    not g578(n56 ,n55);
    nor g579(n55 ,n33 ,n53);
    nor g580(n54 ,n20[5] ,n52);
    nor g581(n569 ,n51 ,n52);
    not g582(n53 ,n52);
    nor g583(n52 ,n40 ,n50);
    nor g584(n51 ,n20[4] ,n49);
    nor g585(n568 ,n48 ,n49);
    not g586(n50 ,n49);
    nor g587(n49 ,n41 ,n47);
    nor g588(n48 ,n20[3] ,n46);
    nor g589(n567 ,n45 ,n46);
    not g590(n47 ,n46);
    nor g591(n46 ,n34 ,n44);
    nor g592(n45 ,n20[2] ,n43);
    nor g593(n566 ,n43 ,n42);
    not g594(n44 ,n43);
    nor g595(n43 ,n37 ,n38);
    nor g596(n42 ,n20[1] ,n20[0]);
    not g597(n41 ,n20[3]);
    not g598(n40 ,n20[4]);
    not g599(n39 ,n20[8]);
    not g600(n38 ,n20[0]);
    not g601(n37 ,n20[1]);
    not g602(n36 ,n20[6]);
    not g603(n35 ,n20[7]);
    not g604(n34 ,n20[2]);
    not g605(n33 ,n20[5]);
    xor g606(n576 ,n14[15] ,n120);
    nor g607(n577 ,n119 ,n120);
    nor g608(n120 ,n76 ,n118);
    nor g609(n119 ,n14[14] ,n117);
    nor g610(n578 ,n116 ,n117);
    not g611(n118 ,n117);
    nor g612(n117 ,n66 ,n115);
    nor g613(n116 ,n14[13] ,n114);
    nor g614(n579 ,n113 ,n114);
    not g615(n115 ,n114);
    nor g616(n114 ,n79 ,n112);
    nor g617(n113 ,n14[12] ,n111);
    nor g618(n580 ,n110 ,n111);
    not g619(n112 ,n111);
    nor g620(n111 ,n75 ,n109);
    nor g621(n110 ,n14[11] ,n108);
    nor g622(n581 ,n107 ,n108);
    not g623(n109 ,n108);
    nor g624(n108 ,n77 ,n106);
    nor g625(n107 ,n14[10] ,n105);
    nor g626(n582 ,n104 ,n105);
    not g627(n106 ,n105);
    nor g628(n105 ,n74 ,n103);
    nor g629(n104 ,n14[9] ,n102);
    nor g630(n583 ,n101 ,n102);
    not g631(n103 ,n102);
    nor g632(n102 ,n71 ,n100);
    nor g633(n101 ,n14[8] ,n99);
    nor g634(n584 ,n98 ,n99);
    not g635(n100 ,n99);
    nor g636(n99 ,n72 ,n97);
    nor g637(n98 ,n14[7] ,n96);
    nor g638(n585 ,n95 ,n96);
    not g639(n97 ,n96);
    nor g640(n96 ,n65 ,n94);
    nor g641(n95 ,n14[6] ,n93);
    nor g642(n586 ,n92 ,n93);
    not g643(n94 ,n93);
    nor g644(n93 ,n70 ,n91);
    nor g645(n92 ,n14[5] ,n90);
    nor g646(n587 ,n89 ,n90);
    not g647(n91 ,n90);
    nor g648(n90 ,n68 ,n88);
    nor g649(n89 ,n14[4] ,n87);
    nor g650(n588 ,n86 ,n87);
    not g651(n88 ,n87);
    nor g652(n87 ,n67 ,n85);
    nor g653(n86 ,n14[3] ,n84);
    nor g654(n589 ,n83 ,n84);
    not g655(n85 ,n84);
    nor g656(n84 ,n69 ,n82);
    nor g657(n83 ,n14[2] ,n81);
    nor g658(n590 ,n81 ,n80);
    not g659(n82 ,n81);
    nor g660(n81 ,n73 ,n78);
    nor g661(n80 ,n14[1] ,n14[0]);
    not g662(n79 ,n14[12]);
    not g663(n78 ,n14[0]);
    not g664(n77 ,n14[10]);
    not g665(n76 ,n14[14]);
    not g666(n75 ,n14[11]);
    not g667(n74 ,n14[9]);
    not g668(n73 ,n14[1]);
    not g669(n72 ,n14[7]);
    not g670(n71 ,n14[8]);
    not g671(n70 ,n14[5]);
    not g672(n69 ,n14[2]);
    not g673(n68 ,n14[4]);
    not g674(n67 ,n14[3]);
    not g675(n66 ,n14[13]);
    not g676(n65 ,n14[6]);
    not g677(n414 ,n310);
    not g678(n538 ,n470);
endmodule
