module top(n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [63:0] n6;
    wire [63:0] n7;
    wire [63:0] n8;
    wire [63:0] n9;
    wire [63:0] n10;
    wire [63:0] n11;
    wire [2:0] n12;
    wire [3:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574;
    wire n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582;
    wire n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590;
    wire n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598;
    wire n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606;
    wire n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614;
    wire n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622;
    wire n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630;
    wire n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;
    wire n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646;
    wire n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
    wire n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662;
    wire n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670;
    wire n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678;
    wire n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686;
    wire n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694;
    wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
    wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
    wire n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718;
    wire n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726;
    wire n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734;
    wire n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742;
    wire n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
    wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
    wire n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766;
    wire n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774;
    wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
    wire n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790;
    wire n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
    wire n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806;
    wire n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814;
    wire n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822;
    wire n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830;
    wire n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838;
    wire n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846;
    wire n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854;
    wire n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862;
    wire n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870;
    wire n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878;
    wire n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886;
    wire n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894;
    wire n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
    wire n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910;
    wire n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918;
    wire n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926;
    wire n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934;
    wire n2935, n2936, n2937, n2938, n2939, n2940;
    not g0(n2488 ,n6[13]);
    not g1(n2487 ,n6[11]);
    not g2(n2486 ,n6[7]);
    not g3(n2485 ,n6[12]);
    not g4(n2484 ,n6[6]);
    not g5(n2483 ,n6[10]);
    not g6(n2482 ,n6[5]);
    not g7(n2481 ,n6[4]);
    not g8(n2480 ,n6[9]);
    not g9(n2479 ,n6[3]);
    not g10(n2478 ,n6[14]);
    not g11(n2477 ,n6[1]);
    not g12(n2476 ,n6[8]);
    not g13(n2475 ,n6[2]);
    xnor g14(n5[45] ,n2462 ,n7[45]);
    xnor g15(n3[47] ,n2474 ,n8[47]);
    xnor g16(n3[16] ,n2466 ,n8[16]);
    xnor g17(n4[16] ,n2466 ,n9[16]);
    xnor g18(n4[15] ,n2474 ,n9[15]);
    xnor g19(n3[15] ,n2474 ,n8[15]);
    xnor g20(n5[48] ,n2466 ,n7[48]);
    xnor g21(n5[47] ,n2474 ,n7[47]);
    xnor g22(n5[32] ,n2466 ,n7[32]);
    xnor g23(n5[31] ,n2474 ,n7[31]);
    xnor g24(n3[32] ,n2466 ,n8[32]);
    xnor g25(n4[48] ,n2466 ,n9[48]);
    xnor g26(n5[16] ,n2466 ,n7[16]);
    xnor g27(n5[15] ,n2474 ,n7[15]);
    xnor g28(n4[47] ,n2474 ,n9[47]);
    xnor g29(n3[31] ,n2474 ,n8[31]);
    xnor g30(n4[32] ,n2466 ,n9[32]);
    xnor g31(n4[31] ,n2474 ,n9[31]);
    xnor g32(n3[51] ,n2471 ,n8[51]);
    xnor g33(n3[28] ,n2468 ,n8[28]);
    xnor g34(n4[29] ,n2462 ,n9[29]);
    xnor g35(n4[28] ,n2468 ,n9[28]);
    xnor g36(n3[27] ,n2464 ,n8[27]);
    xnor g37(n4[27] ,n2464 ,n9[27]);
    xnor g38(n4[26] ,n2460 ,n9[26]);
    xnor g39(n3[26] ,n2460 ,n8[26]);
    xnor g40(n4[25] ,n2470 ,n9[25]);
    xnor g41(n4[24] ,n2467 ,n9[24]);
    xnor g42(n3[25] ,n2470 ,n8[25]);
    xnor g43(n4[23] ,n2465 ,n9[23]);
    xnor g44(n4[22] ,n2463 ,n9[22]);
    xnor g45(n3[23] ,n2465 ,n8[23]);
    xnor g46(n4[21] ,n2461 ,n9[21]);
    xnor g47(n4[20] ,n2459 ,n9[20]);
    xnor g48(n4[19] ,n2471 ,n9[19]);
    xnor g49(n4[18] ,n2469 ,n9[18]);
    xnor g50(n3[57] ,n2470 ,n8[57]);
    xnor g51(n3[22] ,n2463 ,n8[22]);
    xnor g52(n4[17] ,n2473 ,n9[17]);
    xnor g53(n3[24] ,n2467 ,n8[24]);
    xnor g54(n3[21] ,n2461 ,n8[21]);
    xnor g55(n4[14] ,n2472 ,n9[14]);
    xnor g56(n3[50] ,n2469 ,n8[50]);
    xnor g57(n3[20] ,n2459 ,n8[20]);
    xnor g58(n4[13] ,n2462 ,n9[13]);
    xnor g59(n4[12] ,n2468 ,n9[12]);
    xnor g60(n3[19] ,n2471 ,n8[19]);
    xnor g61(n4[11] ,n2464 ,n9[11]);
    xnor g62(n4[10] ,n2460 ,n9[10]);
    xnor g63(n3[18] ,n2469 ,n8[18]);
    xnor g64(n4[9] ,n2470 ,n9[9]);
    xnor g65(n4[8] ,n2467 ,n9[8]);
    xnor g66(n3[17] ,n2473 ,n8[17]);
    xnor g67(n4[7] ,n2465 ,n9[7]);
    xnor g68(n4[6] ,n2463 ,n9[6]);
    xnor g69(n3[60] ,n2468 ,n8[60]);
    xnor g70(n3[56] ,n2467 ,n8[56]);
    xnor g71(n4[5] ,n2461 ,n9[5]);
    xnor g72(n4[4] ,n2459 ,n9[4]);
    xnor g73(n3[49] ,n2473 ,n8[49]);
    xnor g74(n4[3] ,n2471 ,n9[3]);
    xnor g75(n4[2] ,n2469 ,n9[2]);
    xnor g76(n3[14] ,n2472 ,n8[14]);
    xnor g77(n4[1] ,n2473 ,n9[1]);
    xnor g78(n3[13] ,n2462 ,n8[13]);
    xnor g79(n5[62] ,n2472 ,n7[62]);
    xnor g80(n3[12] ,n2468 ,n8[12]);
    xnor g81(n3[11] ,n2464 ,n8[11]);
    xnor g82(n5[61] ,n2462 ,n7[61]);
    xnor g83(n5[60] ,n2468 ,n7[60]);
    xnor g84(n5[59] ,n2464 ,n7[59]);
    xnor g85(n5[58] ,n2460 ,n7[58]);
    xnor g86(n3[10] ,n2460 ,n8[10]);
    xnor g87(n5[57] ,n2470 ,n7[57]);
    xnor g88(n5[56] ,n2467 ,n7[56]);
    xnor g89(n3[9] ,n2470 ,n8[9]);
    xnor g90(n5[55] ,n2465 ,n7[55]);
    xnor g91(n5[54] ,n2463 ,n7[54]);
    xnor g92(n3[62] ,n2472 ,n8[62]);
    xnor g93(n3[7] ,n2465 ,n8[7]);
    xnor g94(n5[53] ,n2461 ,n7[53]);
    xnor g95(n5[52] ,n2459 ,n7[52]);
    xnor g96(n5[51] ,n2471 ,n7[51]);
    xnor g97(n5[50] ,n2469 ,n7[50]);
    xnor g98(n3[59] ,n2464 ,n8[59]);
    xnor g99(n3[6] ,n2463 ,n8[6]);
    xnor g100(n5[49] ,n2473 ,n7[49]);
    xnor g101(n3[8] ,n2467 ,n8[8]);
    xnor g102(n3[5] ,n2461 ,n8[5]);
    xnor g103(n5[46] ,n2472 ,n7[46]);
    xnor g104(n3[55] ,n2465 ,n8[55]);
    xnor g105(n3[4] ,n2459 ,n8[4]);
    xnor g106(n3[48] ,n2466 ,n8[48]);
    xnor g107(n4[30] ,n2472 ,n9[30]);
    xnor g108(n3[3] ,n2471 ,n8[3]);
    xnor g109(n5[43] ,n2464 ,n7[43]);
    xnor g110(n5[42] ,n2460 ,n7[42]);
    xnor g111(n3[2] ,n2469 ,n8[2]);
    xnor g112(n5[41] ,n2470 ,n7[41]);
    xnor g113(n5[40] ,n2467 ,n7[40]);
    xnor g114(n3[1] ,n2473 ,n8[1]);
    xnor g115(n5[39] ,n2465 ,n7[39]);
    xnor g116(n5[38] ,n2463 ,n7[38]);
    xnor g117(n5[37] ,n2461 ,n7[37]);
    xnor g118(n5[36] ,n2459 ,n7[36]);
    xnor g119(n5[35] ,n2471 ,n7[35]);
    xnor g120(n5[34] ,n2469 ,n7[34]);
    xnor g121(n3[61] ,n2462 ,n8[61]);
    xnor g122(n3[45] ,n2462 ,n8[45]);
    xnor g123(n5[33] ,n2473 ,n7[33]);
    xnor g124(n3[46] ,n2472 ,n8[46]);
    xnor g125(n4[62] ,n2472 ,n9[62]);
    xnor g126(n5[30] ,n2472 ,n7[30]);
    xnor g127(n3[43] ,n2464 ,n8[43]);
    xnor g128(n4[61] ,n2462 ,n9[61]);
    xnor g129(n5[29] ,n2462 ,n7[29]);
    xnor g130(n5[28] ,n2468 ,n7[28]);
    xnor g131(n4[60] ,n2468 ,n9[60]);
    xnor g132(n5[27] ,n2464 ,n7[27]);
    xnor g133(n5[26] ,n2460 ,n7[26]);
    xnor g134(n4[59] ,n2464 ,n9[59]);
    xnor g135(n5[25] ,n2470 ,n7[25]);
    xnor g136(n5[24] ,n2467 ,n7[24]);
    xnor g137(n4[58] ,n2460 ,n9[58]);
    xnor g138(n5[23] ,n2465 ,n7[23]);
    xnor g139(n5[22] ,n2463 ,n7[22]);
    xnor g140(n4[57] ,n2470 ,n9[57]);
    xnor g141(n5[21] ,n2461 ,n7[21]);
    xnor g142(n5[20] ,n2459 ,n7[20]);
    xnor g143(n4[56] ,n2467 ,n9[56]);
    xnor g144(n5[19] ,n2471 ,n7[19]);
    xnor g145(n5[18] ,n2469 ,n7[18]);
    xnor g146(n3[44] ,n2468 ,n8[44]);
    xnor g147(n3[41] ,n2470 ,n8[41]);
    xnor g148(n5[17] ,n2473 ,n7[17]);
    xnor g149(n4[55] ,n2465 ,n9[55]);
    xnor g150(n3[42] ,n2460 ,n8[42]);
    xnor g151(n4[54] ,n2463 ,n9[54]);
    xnor g152(n5[14] ,n2472 ,n7[14]);
    xnor g153(n3[40] ,n2467 ,n8[40]);
    xnor g154(n4[53] ,n2461 ,n9[53]);
    xnor g155(n5[13] ,n2462 ,n7[13]);
    xnor g156(n5[12] ,n2468 ,n7[12]);
    xnor g157(n4[52] ,n2459 ,n9[52]);
    xnor g158(n5[11] ,n2464 ,n7[11]);
    xnor g159(n5[10] ,n2460 ,n7[10]);
    xnor g160(n3[39] ,n2465 ,n8[39]);
    xnor g161(n4[51] ,n2471 ,n9[51]);
    xnor g162(n5[9] ,n2470 ,n7[9]);
    xnor g163(n5[8] ,n2467 ,n7[8]);
    xnor g164(n4[50] ,n2469 ,n9[50]);
    xnor g165(n5[7] ,n2465 ,n7[7]);
    xnor g166(n5[6] ,n2463 ,n7[6]);
    xnor g167(n3[54] ,n2463 ,n8[54]);
    xnor g168(n3[38] ,n2463 ,n8[38]);
    xnor g169(n5[5] ,n2461 ,n7[5]);
    xnor g170(n5[4] ,n2459 ,n7[4]);
    xnor g171(n4[49] ,n2473 ,n9[49]);
    xnor g172(n5[3] ,n2471 ,n7[3]);
    xnor g173(n5[2] ,n2469 ,n7[2]);
    xnor g174(n3[53] ,n2461 ,n8[53]);
    xnor g175(n3[37] ,n2461 ,n8[37]);
    xnor g176(n5[1] ,n2473 ,n7[1]);
    xnor g177(n4[46] ,n2472 ,n9[46]);
    xnor g178(n3[36] ,n2459 ,n8[36]);
    xnor g179(n3[35] ,n2471 ,n8[35]);
    xnor g180(n4[45] ,n2462 ,n9[45]);
    xnor g181(n4[44] ,n2468 ,n9[44]);
    xnor g182(n4[43] ,n2464 ,n9[43]);
    xnor g183(n4[42] ,n2460 ,n9[42]);
    xnor g184(n3[34] ,n2469 ,n8[34]);
    xnor g185(n4[41] ,n2470 ,n9[41]);
    xnor g186(n4[40] ,n2467 ,n9[40]);
    xnor g187(n3[33] ,n2473 ,n8[33]);
    xnor g188(n4[39] ,n2465 ,n9[39]);
    xnor g189(n4[38] ,n2463 ,n9[38]);
    xnor g190(n3[52] ,n2459 ,n8[52]);
    xnor g191(n4[37] ,n2461 ,n9[37]);
    xnor g192(n4[36] ,n2459 ,n9[36]);
    xnor g193(n4[35] ,n2471 ,n9[35]);
    xnor g194(n4[34] ,n2469 ,n9[34]);
    xnor g195(n3[30] ,n2472 ,n8[30]);
    xnor g196(n4[33] ,n2473 ,n9[33]);
    xnor g197(n3[58] ,n2460 ,n8[58]);
    xnor g198(n3[29] ,n2462 ,n8[29]);
    xnor g199(n5[44] ,n2468 ,n7[44]);
    xnor g200(n4[0] ,n2457 ,n9[0]);
    xnor g201(n5[63] ,n2458 ,n7[63]);
    xnor g202(n3[0] ,n2457 ,n8[0]);
    xnor g203(n4[63] ,n2458 ,n9[63]);
    xnor g204(n3[63] ,n2458 ,n8[63]);
    xnor g205(n5[0] ,n2457 ,n7[0]);
    xnor g206(n2474 ,n10[47] ,n2448);
    xnor g207(n2473 ,n10[49] ,n2445);
    xnor g208(n2472 ,n10[62] ,n2441);
    xnor g209(n2471 ,n10[51] ,n2456);
    xnor g210(n2470 ,n10[57] ,n2442);
    xnor g211(n2469 ,n10[50] ,n2443);
    xnor g212(n2468 ,n10[60] ,n2444);
    xnor g213(n2467 ,n10[56] ,n2446);
    xnor g214(n2466 ,n10[48] ,n2447);
    xnor g215(n2465 ,n10[55] ,n2449);
    xnor g216(n2464 ,n10[59] ,n2450);
    xnor g217(n2463 ,n10[54] ,n2451);
    xnor g218(n2462 ,n10[61] ,n2452);
    xnor g219(n2461 ,n10[53] ,n2453);
    xnor g220(n2460 ,n10[58] ,n2454);
    xnor g221(n2459 ,n10[52] ,n2455);
    xnor g222(n2458 ,n10[47] ,n2433);
    xnor g223(n2457 ,n10[48] ,n2432);
    xnor g224(n2867 ,n2405 ,n2868);
    xnor g225(n2721 ,n2414 ,n2[40]);
    xnor g226(n2722 ,n2418 ,n2[41]);
    xnor g227(n2723 ,n2421 ,n2[42]);
    xnor g228(n2724 ,n2407 ,n2[43]);
    xnor g229(n2725 ,n2415 ,n2[44]);
    xnor g230(n2726 ,n2410 ,n2[45]);
    xnor g231(n2564 ,n2[75] ,n2407);
    xnor g232(n2729 ,n2420 ,n2[48]);
    xnor g233(n2731 ,n2409 ,n2[50]);
    xnor g234(n2732 ,n2416 ,n2[51]);
    xnor g235(n2733 ,n2408 ,n2[52]);
    xnor g236(n2734 ,n2417 ,n2[53]);
    xnor g237(n2735 ,n2411 ,n2[54]);
    xnor g238(n2736 ,n2419 ,n2[55]);
    xnor g239(n2737 ,n2414 ,n2[56]);
    xnor g240(n2837 ,n2413 ,n2838);
    xnor g241(n2712 ,n2413 ,n2[31]);
    xnor g242(n2744 ,n2[63] ,n2413);
    xnor g243(n2728 ,n2413 ,n2[47]);
    xnor g244(n2568 ,n2[79] ,n2413);
    xnor g245(n2696 ,n2413 ,n2[15]);
    xnor g246(n2616 ,n2[127] ,n2413);
    xnor g247(n2600 ,n2[111] ,n2413);
    xnor g248(n2584 ,n2[95] ,n2413);
    xnor g249(n2933 ,n2413 ,n2934);
    xnor g250(n2901 ,n2413 ,n2902);
    xnor g251(n2869 ,n2413 ,n2870);
    xnor g252(n2841 ,n2406 ,n2842);
    xnor g253(n2835 ,n2405 ,n2836);
    xnor g254(n2809 ,n2810 ,n2406);
    xnor g255(n2743 ,n2[62] ,n2405);
    xnor g256(n2730 ,n2406 ,n2[49]);
    xnor g257(n2727 ,n2405 ,n2[46]);
    xnor g258(n2714 ,n2406 ,n2[33]);
    xnor g259(n2711 ,n2405 ,n2[30]);
    xnor g260(n2615 ,n2[126] ,n2405);
    xnor g261(n2698 ,n2406 ,n2[17]);
    xnor g262(n2695 ,n2405 ,n2[14]);
    xnor g263(n2682 ,n2406 ,n2[1]);
    xnor g264(n2602 ,n2[113] ,n2406);
    xnor g265(n2599 ,n2[110] ,n2405);
    xnor g266(n2586 ,n2[97] ,n2406);
    xnor g267(n2583 ,n2[94] ,n2405);
    xnor g268(n2570 ,n2[81] ,n2406);
    xnor g269(n2567 ,n2[78] ,n2405);
    xnor g270(n2554 ,n2[65] ,n2406);
    xnor g271(n2931 ,n2405 ,n2932);
    xnor g272(n2905 ,n2406 ,n2906);
    xnor g273(n2899 ,n2405 ,n2900);
    xnor g274(n2873 ,n2406 ,n2874);
    xnor g275(n2738 ,n2418 ,n2[57]);
    xnor g276(n2865 ,n2410 ,n2866);
    xnor g277(n2863 ,n2415 ,n2864);
    xnor g278(n2603 ,n2[114] ,n2409);
    xnor g279(n2861 ,n2407 ,n2862);
    xnor g280(n2859 ,n2421 ,n2860);
    xnor g281(n2857 ,n2418 ,n2858);
    xnor g282(n2855 ,n2414 ,n2856);
    xnor g283(n2853 ,n2419 ,n2854);
    xnor g284(n2851 ,n2411 ,n2852);
    xnor g285(n2849 ,n2417 ,n2850);
    xnor g286(n2605 ,n2[116] ,n2408);
    xnor g287(n2847 ,n2408 ,n2848);
    xnor g288(n2845 ,n2416 ,n2846);
    xnor g289(n2843 ,n2409 ,n2844);
    xnor g290(n2839 ,n2420 ,n2840);
    xnor g291(n2833 ,n2410 ,n2834);
    xnor g292(n2831 ,n2415 ,n2832);
    xnor g293(n2829 ,n2407 ,n2830);
    xnor g294(n2827 ,n2421 ,n2828);
    xnor g295(n2825 ,n2418 ,n2826);
    xnor g296(n2823 ,n2414 ,n2824);
    xnor g297(n2821 ,n2419 ,n2822);
    xnor g298(n2819 ,n2411 ,n2820);
    xnor g299(n2607 ,n2[118] ,n2411);
    xnor g300(n2817 ,n2417 ,n2818);
    xnor g301(n2561 ,n2[72] ,n2414);
    xnor g302(n2815 ,n2408 ,n2816);
    xnor g303(n2713 ,n2420 ,n2[32]);
    xnor g304(n2813 ,n2416 ,n2814);
    xnor g305(n2560 ,n2[71] ,n2419);
    xnor g306(n2811 ,n2409 ,n2812);
    xnor g307(n2742 ,n2[61] ,n2410);
    xnor g308(n2741 ,n2[60] ,n2415);
    xnor g309(n2740 ,n2407 ,n2[59]);
    xnor g310(n2739 ,n2421 ,n2[58]);
    nor g311(n2456 ,n2479 ,n2426);
    nor g312(n2455 ,n2481 ,n2437);
    nor g313(n2454 ,n2483 ,n2439);
    nor g314(n2453 ,n2482 ,n2424);
    nor g315(n2452 ,n2488 ,n2431);
    nor g316(n2451 ,n2484 ,n2428);
    nor g317(n2450 ,n2487 ,n2429);
    nor g318(n2449 ,n2486 ,n2438);
    nor g319(n2448 ,n2422 ,n2436);
    nor g320(n2447 ,n2412 ,n2434);
    nor g321(n2446 ,n2476 ,n2423);
    nor g322(n2445 ,n2477 ,n2425);
    nor g323(n2444 ,n2485 ,n2427);
    nor g324(n2443 ,n2475 ,n2435);
    nor g325(n2442 ,n2480 ,n2440);
    nor g326(n2441 ,n2478 ,n2430);
    xnor g327(n2720 ,n2419 ,n2[39]);
    xnor g328(n2719 ,n2411 ,n2[38]);
    xnor g329(n2718 ,n2417 ,n2[37]);
    xnor g330(n2717 ,n2408 ,n2[36]);
    xnor g331(n2716 ,n2416 ,n2[35]);
    xnor g332(n2715 ,n2409 ,n2[34]);
    xnor g333(n2710 ,n2410 ,n2[29]);
    xnor g334(n2709 ,n2415 ,n2[28]);
    xnor g335(n2708 ,n2407 ,n2[27]);
    xnor g336(n2707 ,n2421 ,n2[26]);
    xnor g337(n2706 ,n2418 ,n2[25]);
    xnor g338(n2705 ,n2414 ,n2[24]);
    xnor g339(n2704 ,n2419 ,n2[23]);
    xnor g340(n2703 ,n2411 ,n2[22]);
    xnor g341(n2702 ,n2417 ,n2[21]);
    xnor g342(n2701 ,n2408 ,n2[20]);
    xnor g343(n2569 ,n2[80] ,n2420);
    xnor g344(n2700 ,n2416 ,n2[19]);
    xnor g345(n2697 ,n2420 ,n2[16]);
    xnor g346(n2694 ,n2410 ,n2[13]);
    xnor g347(n2693 ,n2415 ,n2[12]);
    xnor g348(n2692 ,n2407 ,n2[11]);
    xnor g349(n2691 ,n2421 ,n2[10]);
    xnor g350(n2690 ,n2418 ,n2[9]);
    xnor g351(n2689 ,n2414 ,n2[8]);
    xnor g352(n2681 ,n2[0] ,n2420);
    xnor g353(n2688 ,n2419 ,n2[7]);
    xnor g354(n2687 ,n2411 ,n2[6]);
    xnor g355(n2571 ,n2[82] ,n2409);
    xnor g356(n2686 ,n2417 ,n2[5]);
    xnor g357(n2685 ,n2408 ,n2[4]);
    xnor g358(n2573 ,n2[84] ,n2408);
    xnor g359(n2684 ,n2416 ,n2[3]);
    xnor g360(n2683 ,n2409 ,n2[2]);
    xnor g361(n2572 ,n2[83] ,n2416);
    xnor g362(n2614 ,n2[125] ,n2410);
    xnor g363(n2613 ,n2[124] ,n2415);
    xnor g364(n2612 ,n2[123] ,n2407);
    xnor g365(n2611 ,n2[122] ,n2421);
    xnor g366(n2610 ,n2[121] ,n2418);
    xnor g367(n2609 ,n2[120] ,n2414);
    xnor g368(n2608 ,n2[119] ,n2419);
    xnor g369(n2606 ,n2[117] ,n2417);
    xnor g370(n2604 ,n2[115] ,n2416);
    xnor g371(n2601 ,n2[112] ,n2420);
    xnor g372(n2576 ,n2[87] ,n2419);
    xnor g373(n2598 ,n2[109] ,n2410);
    xnor g374(n2594 ,n2[105] ,n2418);
    xnor g375(n2591 ,n2[102] ,n2411);
    xnor g376(n2590 ,n2[101] ,n2417);
    xnor g377(n2589 ,n2[100] ,n2408);
    xnor g378(n2585 ,n2[96] ,n2420);
    xnor g379(n2582 ,n2[93] ,n2410);
    xnor g380(n2581 ,n2[92] ,n2415);
    xnor g381(n2555 ,n2[66] ,n2409);
    xnor g382(n2579 ,n2[90] ,n2421);
    xnor g383(n2578 ,n2[89] ,n2418);
    xnor g384(n2577 ,n2[88] ,n2414);
    xnor g385(n2556 ,n2[67] ,n2416);
    xnor g386(n2575 ,n2[86] ,n2411);
    xnor g387(n2580 ,n2[91] ,n2407);
    xnor g388(n2574 ,n2[85] ,n2417);
    xnor g389(n2566 ,n2[77] ,n2410);
    xnor g390(n2565 ,n2[76] ,n2415);
    xnor g391(n2563 ,n2[74] ,n2421);
    xnor g392(n2562 ,n2[73] ,n2418);
    xnor g393(n2559 ,n2[70] ,n2411);
    xnor g394(n2558 ,n2[69] ,n2417);
    xnor g395(n2557 ,n2[68] ,n2408);
    xnor g396(n2553 ,n2[64] ,n2420);
    xnor g397(n2587 ,n2[98] ,n2409);
    xnor g398(n2588 ,n2[99] ,n2416);
    xnor g399(n2699 ,n2409 ,n2[18]);
    xnor g400(n2592 ,n2[103] ,n2419);
    xnor g401(n2929 ,n2410 ,n2930);
    xnor g402(n2927 ,n2415 ,n2928);
    xnor g403(n2925 ,n2407 ,n2926);
    xnor g404(n2595 ,n2[106] ,n2421);
    xnor g405(n2923 ,n2421 ,n2924);
    xnor g406(n2921 ,n2418 ,n2922);
    xnor g407(n2593 ,n2[104] ,n2414);
    xnor g408(n2919 ,n2414 ,n2920);
    xnor g409(n2917 ,n2419 ,n2918);
    xnor g410(n2915 ,n2411 ,n2916);
    xnor g411(n2913 ,n2417 ,n2914);
    xnor g412(n2911 ,n2408 ,n2912);
    xnor g413(n2909 ,n2416 ,n2910);
    xnor g414(n2907 ,n2409 ,n2908);
    xnor g415(n2903 ,n2420 ,n2904);
    xnor g416(n2897 ,n2410 ,n2898);
    xnor g417(n2895 ,n2415 ,n2896);
    xnor g418(n2893 ,n2407 ,n2894);
    xnor g419(n2891 ,n2421 ,n2892);
    xnor g420(n2889 ,n2418 ,n2890);
    xnor g421(n2887 ,n2414 ,n2888);
    xnor g422(n2885 ,n2419 ,n2886);
    xnor g423(n2596 ,n2[107] ,n2407);
    xnor g424(n2883 ,n2411 ,n2884);
    xnor g425(n2881 ,n2417 ,n2882);
    xnor g426(n2879 ,n2408 ,n2880);
    xnor g427(n2877 ,n2416 ,n2878);
    xnor g428(n2875 ,n2409 ,n2876);
    xnor g429(n2597 ,n2[108] ,n2415);
    xnor g430(n2871 ,n2420 ,n2872);
    not g431(n11[41] ,n2440);
    not g432(n11[42] ,n2439);
    not g433(n11[39] ,n2438);
    not g434(n11[36] ,n2437);
    not g435(n11[31] ,n2436);
    not g436(n11[34] ,n2435);
    not g437(n11[32] ,n2434);
    nor g438(n2440 ,n10[58] ,n10[56]);
    nor g439(n2433 ,n2405 ,n2422);
    nor g440(n2439 ,n10[59] ,n10[57]);
    nor g441(n2438 ,n10[56] ,n10[54]);
    nor g442(n2437 ,n10[53] ,n10[51]);
    nor g443(n2436 ,n10[62] ,n10[48]);
    nor g444(n2435 ,n10[51] ,n10[49]);
    nor g445(n2434 ,n10[47] ,n10[49]);
    nor g446(n2432 ,n2406 ,n2412);
    not g447(n11[45] ,n2431);
    not g448(n11[46] ,n2430);
    not g449(n11[43] ,n2429);
    not g450(n11[38] ,n2428);
    not g451(n11[44] ,n2427);
    not g452(n11[35] ,n2426);
    not g453(n11[33] ,n2425);
    not g454(n11[37] ,n2424);
    not g455(n11[40] ,n2423);
    nor g456(n2431 ,n10[62] ,n10[60]);
    nor g457(n2430 ,n10[47] ,n10[61]);
    nor g458(n2429 ,n10[60] ,n10[58]);
    nor g459(n2428 ,n10[55] ,n10[53]);
    nor g460(n2427 ,n10[61] ,n10[59]);
    nor g461(n2426 ,n10[52] ,n10[50]);
    nor g462(n2425 ,n10[50] ,n10[48]);
    nor g463(n2424 ,n10[54] ,n10[52]);
    nor g464(n2423 ,n10[57] ,n10[55]);
    not g465(n2422 ,n6[15]);
    not g466(n2421 ,n10[58]);
    not g467(n2420 ,n10[48]);
    not g468(n2419 ,n10[55]);
    not g469(n2418 ,n10[57]);
    not g470(n2417 ,n10[53]);
    not g471(n2416 ,n10[51]);
    not g472(n2415 ,n10[60]);
    not g473(n2414 ,n10[56]);
    not g474(n2413 ,n10[47]);
    not g475(n2412 ,n6[0]);
    not g476(n2411 ,n10[54]);
    not g477(n2410 ,n10[61]);
    not g478(n2409 ,n10[50]);
    not g479(n2408 ,n10[52]);
    not g480(n2407 ,n10[59]);
    not g481(n2406 ,n10[49]);
    not g482(n2405 ,n10[62]);
    dff g483(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n7[0]));
    dff g484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2217), .Q(n7[1]));
    dff g485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n7[2]));
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n7[3]));
    dff g487(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2182), .Q(n7[4]));
    dff g488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n7[5]));
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n7[6]));
    dff g490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n7[7]));
    dff g491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2163), .Q(n7[8]));
    dff g492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2159), .Q(n7[9]));
    dff g493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2337), .Q(n7[10]));
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2330), .Q(n7[11]));
    dff g495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2335), .Q(n7[12]));
    dff g496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2332), .Q(n7[13]));
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2323), .Q(n7[14]));
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2322), .Q(n7[15]));
    dff g499(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2316), .Q(n7[16]));
    dff g500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2312), .Q(n7[17]));
    dff g501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2311), .Q(n7[18]));
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2305), .Q(n7[19]));
    dff g503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2308), .Q(n7[20]));
    dff g504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2302), .Q(n7[21]));
    dff g505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2298), .Q(n7[22]));
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2296), .Q(n7[23]));
    dff g507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2294), .Q(n7[24]));
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2282), .Q(n7[25]));
    dff g509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2289), .Q(n7[26]));
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2285), .Q(n7[27]));
    dff g511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2280), .Q(n7[28]));
    dff g512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2278), .Q(n7[29]));
    dff g513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2273), .Q(n7[30]));
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2270), .Q(n7[31]));
    dff g515(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n7[32]));
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2267), .Q(n7[33]));
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2265), .Q(n7[34]));
    dff g518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2261), .Q(n7[35]));
    dff g519(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2259), .Q(n7[36]));
    dff g520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2256), .Q(n7[37]));
    dff g521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2253), .Q(n7[38]));
    dff g522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2251), .Q(n7[39]));
    dff g523(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2248), .Q(n7[40]));
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2243), .Q(n7[41]));
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2241), .Q(n7[42]));
    dff g526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2239), .Q(n7[43]));
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2235), .Q(n7[44]));
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2230), .Q(n7[45]));
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2228), .Q(n7[46]));
    dff g530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2226), .Q(n7[47]));
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2224), .Q(n7[48]));
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2223), .Q(n7[49]));
    dff g533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2279), .Q(n7[50]));
    dff g534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2286), .Q(n7[51]));
    dff g535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2222), .Q(n7[52]));
    dff g536(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2221), .Q(n7[53]));
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2220), .Q(n7[54]));
    dff g538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2219), .Q(n7[55]));
    dff g539(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2218), .Q(n7[56]));
    dff g540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2215), .Q(n7[57]));
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2214), .Q(n7[58]));
    dff g542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2216), .Q(n7[59]));
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2213), .Q(n7[60]));
    dff g544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2212), .Q(n7[61]));
    dff g545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2211), .Q(n7[62]));
    dff g546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2210), .Q(n7[63]));
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2209), .Q(n8[0]));
    dff g548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2208), .Q(n8[1]));
    dff g549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2207), .Q(n8[2]));
    dff g550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2206), .Q(n8[3]));
    dff g551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2205), .Q(n8[4]));
    dff g552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2204), .Q(n8[5]));
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2201), .Q(n8[6]));
    dff g554(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2203), .Q(n8[7]));
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2202), .Q(n8[8]));
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2200), .Q(n8[9]));
    dff g557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2199), .Q(n8[10]));
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2198), .Q(n8[11]));
    dff g559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2197), .Q(n8[12]));
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2195), .Q(n8[13]));
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2196), .Q(n8[14]));
    dff g562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2194), .Q(n8[15]));
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n8[16]));
    dff g564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n8[17]));
    dff g565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2191), .Q(n8[18]));
    dff g566(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2189), .Q(n8[19]));
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n8[20]));
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n8[21]));
    dff g569(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n8[22]));
    dff g570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n8[23]));
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2183), .Q(n8[24]));
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2181), .Q(n8[25]));
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2180), .Q(n8[26]));
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n8[27]));
    dff g575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n8[28]));
    dff g576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n8[29]));
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n8[30]));
    dff g578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n8[31]));
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n8[32]));
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n8[33]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n8[34]));
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n8[35]));
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n8[36]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n8[37]));
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2164), .Q(n8[38]));
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2162), .Q(n8[39]));
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2161), .Q(n8[40]));
    dff g588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2160), .Q(n8[41]));
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2158), .Q(n8[42]));
    dff g590(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2157), .Q(n8[43]));
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2269), .Q(n8[44]));
    dff g592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2342), .Q(n8[45]));
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2343), .Q(n8[46]));
    dff g594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2341), .Q(n8[47]));
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2340), .Q(n8[48]));
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2339), .Q(n8[49]));
    dff g597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2338), .Q(n8[50]));
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2336), .Q(n8[51]));
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2334), .Q(n8[52]));
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2333), .Q(n8[53]));
    dff g601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2331), .Q(n8[54]));
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2329), .Q(n8[55]));
    dff g603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2328), .Q(n8[56]));
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2327), .Q(n8[57]));
    dff g605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2326), .Q(n8[58]));
    dff g606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2325), .Q(n8[59]));
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2324), .Q(n8[60]));
    dff g608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2321), .Q(n8[61]));
    dff g609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2320), .Q(n8[62]));
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2319), .Q(n8[63]));
    dff g611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2318), .Q(n9[0]));
    dff g612(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2317), .Q(n9[1]));
    dff g613(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2315), .Q(n9[2]));
    dff g614(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2314), .Q(n9[3]));
    dff g615(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2313), .Q(n9[4]));
    dff g616(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2310), .Q(n9[5]));
    dff g617(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2309), .Q(n9[6]));
    dff g618(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2307), .Q(n9[7]));
    dff g619(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2306), .Q(n9[8]));
    dff g620(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2304), .Q(n9[9]));
    dff g621(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2303), .Q(n9[10]));
    dff g622(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2301), .Q(n9[11]));
    dff g623(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2300), .Q(n9[12]));
    dff g624(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2299), .Q(n9[13]));
    dff g625(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2297), .Q(n9[14]));
    dff g626(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2295), .Q(n9[15]));
    dff g627(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2293), .Q(n9[16]));
    dff g628(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2292), .Q(n9[17]));
    dff g629(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2291), .Q(n9[18]));
    dff g630(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2290), .Q(n9[19]));
    dff g631(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2288), .Q(n9[20]));
    dff g632(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2287), .Q(n9[21]));
    dff g633(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2284), .Q(n9[22]));
    dff g634(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2283), .Q(n9[23]));
    dff g635(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2281), .Q(n9[24]));
    dff g636(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2277), .Q(n9[25]));
    dff g637(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2276), .Q(n9[26]));
    dff g638(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2275), .Q(n9[27]));
    dff g639(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2274), .Q(n9[28]));
    dff g640(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2272), .Q(n9[29]));
    dff g641(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2271), .Q(n9[30]));
    dff g642(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2344), .Q(n9[31]));
    dff g643(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n9[32]));
    dff g644(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n9[33]));
    dff g645(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2156), .Q(n9[34]));
    dff g646(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2268), .Q(n9[35]));
    dff g647(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2266), .Q(n9[36]));
    dff g648(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2264), .Q(n9[37]));
    dff g649(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2263), .Q(n9[38]));
    dff g650(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2262), .Q(n9[39]));
    dff g651(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2260), .Q(n9[40]));
    dff g652(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2258), .Q(n9[41]));
    dff g653(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2257), .Q(n9[42]));
    dff g654(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2255), .Q(n9[43]));
    dff g655(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2254), .Q(n9[44]));
    dff g656(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2252), .Q(n9[45]));
    dff g657(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2250), .Q(n9[46]));
    dff g658(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2249), .Q(n9[47]));
    dff g659(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2247), .Q(n9[48]));
    dff g660(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2246), .Q(n9[49]));
    dff g661(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2245), .Q(n9[50]));
    dff g662(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2244), .Q(n9[51]));
    dff g663(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2242), .Q(n9[52]));
    dff g664(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2240), .Q(n9[53]));
    dff g665(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2238), .Q(n9[54]));
    dff g666(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2237), .Q(n9[55]));
    dff g667(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2236), .Q(n9[56]));
    dff g668(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2234), .Q(n9[57]));
    dff g669(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2233), .Q(n9[58]));
    dff g670(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2232), .Q(n9[59]));
    dff g671(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2231), .Q(n9[60]));
    dff g672(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2229), .Q(n9[61]));
    dff g673(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2227), .Q(n9[62]));
    dff g674(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2225), .Q(n9[63]));
    dff g675(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2383), .Q(n6[0]));
    dff g676(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2384), .Q(n6[1]));
    dff g677(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2385), .Q(n6[2]));
    dff g678(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2386), .Q(n6[3]));
    dff g679(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2387), .Q(n6[4]));
    dff g680(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2388), .Q(n6[5]));
    dff g681(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2389), .Q(n6[6]));
    dff g682(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2390), .Q(n6[7]));
    dff g683(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n6[8]));
    dff g684(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n6[9]));
    dff g685(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2393), .Q(n6[10]));
    dff g686(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n6[11]));
    dff g687(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2395), .Q(n6[12]));
    dff g688(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2396), .Q(n6[13]));
    dff g689(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2397), .Q(n6[14]));
    dff g690(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2398), .Q(n6[15]));
    dff g691(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n12[0]));
    dff g692(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n12[1]));
    dff g693(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n12[2]));
    dff g694(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2401), .Q(n13[0]));
    dff g695(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2404), .Q(n13[1]));
    dff g696(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2400), .Q(n13[2]));
    nor g697(n2404 ,n1 ,n2403);
    nor g698(n2403 ,n1522 ,n2402);
    nor g699(n2402 ,n1477 ,n2399);
    nor g700(n2401 ,n1 ,n2399);
    nor g701(n2400 ,n1 ,n2382);
    or g702(n2398 ,n2346 ,n2345);
    or g703(n2397 ,n2348 ,n2347);
    or g704(n2396 ,n2350 ,n2349);
    or g705(n2395 ,n2352 ,n2351);
    or g706(n2394 ,n2354 ,n2353);
    or g707(n2393 ,n2356 ,n2355);
    or g708(n2392 ,n2358 ,n2357);
    or g709(n2391 ,n2360 ,n2359);
    or g710(n2390 ,n2362 ,n2361);
    or g711(n2389 ,n2364 ,n2363);
    or g712(n2388 ,n2375 ,n2365);
    or g713(n2387 ,n2374 ,n2366);
    or g714(n2386 ,n2376 ,n2367);
    or g715(n2385 ,n2373 ,n2368);
    or g716(n2384 ,n2372 ,n2369);
    or g717(n2383 ,n2371 ,n2370);
    or g718(n2382 ,n13[2] ,n2381);
    or g719(n2399 ,n1496 ,n2380);
    not g720(n2381 ,n2380);
    or g721(n2379 ,n1877 ,n2075);
    or g722(n2378 ,n1879 ,n2076);
    or g723(n2377 ,n1876 ,n2078);
    nor g724(n2376 ,n1481 ,n2056);
    nor g725(n2375 ,n1480 ,n2056);
    nor g726(n2374 ,n1485 ,n2056);
    nor g727(n2373 ,n1474 ,n2056);
    nor g728(n2372 ,n1483 ,n2056);
    nor g729(n2371 ,n1486 ,n2056);
    nor g730(n2370 ,n1262 ,n2155);
    nor g731(n2369 ,n1270 ,n2155);
    nor g732(n2368 ,n1267 ,n2155);
    nor g733(n2367 ,n1266 ,n2155);
    nor g734(n2366 ,n1276 ,n2155);
    nor g735(n2365 ,n1268 ,n2155);
    nor g736(n2364 ,n1475 ,n2056);
    nor g737(n2363 ,n1271 ,n2155);
    nor g738(n2362 ,n1487 ,n2056);
    nor g739(n2361 ,n1273 ,n2155);
    nor g740(n2360 ,n1484 ,n2056);
    nor g741(n2359 ,n1264 ,n2155);
    nor g742(n2358 ,n1482 ,n2056);
    nor g743(n2357 ,n1265 ,n2155);
    nor g744(n2356 ,n1478 ,n2056);
    nor g745(n2355 ,n1277 ,n2155);
    nor g746(n2354 ,n1471 ,n2056);
    nor g747(n2353 ,n1275 ,n2155);
    nor g748(n2352 ,n1476 ,n2056);
    nor g749(n2351 ,n1272 ,n2155);
    nor g750(n2350 ,n1473 ,n2056);
    nor g751(n2349 ,n1263 ,n2155);
    nor g752(n2348 ,n1472 ,n2056);
    nor g753(n2347 ,n1269 ,n2155);
    nor g754(n2346 ,n1479 ,n2056);
    nor g755(n2345 ,n1274 ,n2155);
    or g756(n2344 ,n1939 ,n2077);
    or g757(n2343 ,n1954 ,n2150);
    or g758(n2342 ,n1956 ,n2151);
    or g759(n2341 ,n1953 ,n2148);
    or g760(n2340 ,n1951 ,n2147);
    or g761(n2339 ,n1949 ,n2146);
    or g762(n2338 ,n1947 ,n2145);
    or g763(n2337 ,n1948 ,n2153);
    or g764(n2336 ,n1946 ,n2144);
    or g765(n2335 ,n1944 ,n2143);
    or g766(n2334 ,n1943 ,n2142);
    or g767(n2333 ,n1942 ,n2141);
    or g768(n2332 ,n1937 ,n2139);
    or g769(n2331 ,n1940 ,n2140);
    or g770(n2330 ,n1950 ,n2149);
    or g771(n2329 ,n1938 ,n2138);
    or g772(n2328 ,n1936 ,n2137);
    or g773(n2327 ,n1935 ,n2136);
    or g774(n2326 ,n1934 ,n2134);
    or g775(n2325 ,n1752 ,n2133);
    or g776(n2324 ,n1930 ,n2132);
    or g777(n2323 ,n1932 ,n2135);
    or g778(n2322 ,n1928 ,n2130);
    or g779(n2321 ,n1929 ,n2131);
    or g780(n2320 ,n1927 ,n2129);
    or g781(n2319 ,n1926 ,n2128);
    or g782(n2318 ,n1924 ,n2127);
    or g783(n2317 ,n1922 ,n2126);
    or g784(n2316 ,n1923 ,n2125);
    or g785(n2315 ,n1786 ,n2124);
    or g786(n2314 ,n1921 ,n2122);
    or g787(n2313 ,n1919 ,n2121);
    or g788(n2312 ,n1920 ,n2123);
    or g789(n2311 ,n1807 ,n2120);
    or g790(n2310 ,n1918 ,n2119);
    or g791(n2309 ,n1917 ,n2117);
    or g792(n2308 ,n1912 ,n2113);
    or g793(n2307 ,n1916 ,n2115);
    or g794(n2306 ,n1914 ,n2114);
    or g795(n2305 ,n1915 ,n2116);
    or g796(n2304 ,n1913 ,n2112);
    or g797(n2303 ,n1911 ,n2111);
    or g798(n2302 ,n1910 ,n2109);
    or g799(n2301 ,n1909 ,n2110);
    or g800(n2300 ,n1907 ,n2107);
    or g801(n2299 ,n1905 ,n2106);
    or g802(n2298 ,n1906 ,n2108);
    or g803(n2297 ,n1903 ,n2154);
    or g804(n2296 ,n1901 ,n2101);
    or g805(n2295 ,n1863 ,n2103);
    or g806(n2294 ,n1899 ,n2099);
    or g807(n2293 ,n1900 ,n2102);
    or g808(n2292 ,n1898 ,n2100);
    or g809(n2291 ,n1890 ,n2098);
    or g810(n2290 ,n1894 ,n2097);
    or g811(n2289 ,n1887 ,n2094);
    or g812(n2288 ,n1892 ,n2095);
    or g813(n2287 ,n1891 ,n2093);
    or g814(n2286 ,n1897 ,n2104);
    or g815(n2285 ,n1889 ,n2089);
    or g816(n2284 ,n1895 ,n2092);
    or g817(n2283 ,n1888 ,n2091);
    or g818(n2282 ,n1893 ,n2096);
    or g819(n2281 ,n1902 ,n2090);
    or g820(n2280 ,n1885 ,n2086);
    or g821(n2279 ,n1881 ,n2080);
    or g822(n2278 ,n1884 ,n2084);
    or g823(n2277 ,n1886 ,n2088);
    or g824(n2276 ,n1955 ,n2087);
    or g825(n2275 ,n1883 ,n2085);
    or g826(n2274 ,n1882 ,n2083);
    or g827(n2273 ,n1931 ,n2082);
    or g828(n2272 ,n1880 ,n2081);
    or g829(n2271 ,n1945 ,n2079);
    or g830(n2270 ,n1941 ,n2070);
    nor g831(n2380 ,n1477 ,n1961);
    or g832(n2269 ,n1904 ,n2152);
    or g833(n2268 ,n1874 ,n2072);
    or g834(n2267 ,n1873 ,n2073);
    or g835(n2266 ,n1872 ,n2071);
    or g836(n2265 ,n1820 ,n2069);
    or g837(n2264 ,n1819 ,n2068);
    or g838(n2263 ,n1870 ,n2067);
    or g839(n2262 ,n1869 ,n2027);
    or g840(n2261 ,n1871 ,n2064);
    or g841(n2260 ,n1816 ,n2065);
    or g842(n2259 ,n1867 ,n2063);
    or g843(n2258 ,n1868 ,n2062);
    or g844(n2257 ,n1866 ,n2061);
    or g845(n2256 ,n1865 ,n2059);
    or g846(n2255 ,n1864 ,n2060);
    or g847(n2254 ,n1862 ,n2058);
    or g848(n2253 ,n1861 ,n2054);
    or g849(n2252 ,n1860 ,n2105);
    or g850(n2251 ,n1858 ,n2051);
    or g851(n2250 ,n1859 ,n2006);
    or g852(n2249 ,n1764 ,n2053);
    or g853(n2248 ,n1855 ,n2049);
    or g854(n2247 ,n1856 ,n2052);
    or g855(n2246 ,n1778 ,n2050);
    or g856(n2245 ,n1812 ,n2048);
    or g857(n2244 ,n1852 ,n2047);
    or g858(n2243 ,n1853 ,n2045);
    or g859(n2242 ,n1794 ,n2046);
    or g860(n2241 ,n1804 ,n2044);
    or g861(n2240 ,n1814 ,n2043);
    or g862(n2239 ,n1831 ,n2039);
    or g863(n2238 ,n1832 ,n2042);
    or g864(n2237 ,n1830 ,n2041);
    or g865(n2236 ,n1817 ,n2040);
    or g866(n2235 ,n1826 ,n2034);
    or g867(n2234 ,n1827 ,n2038);
    or g868(n2233 ,n1821 ,n2036);
    or g869(n2232 ,n1825 ,n2035);
    or g870(n2231 ,n1823 ,n2033);
    or g871(n2230 ,n1824 ,n2037);
    or g872(n2229 ,n1828 ,n2031);
    or g873(n2228 ,n1818 ,n2032);
    or g874(n2227 ,n1748 ,n2030);
    or g875(n2226 ,n1857 ,n2029);
    or g876(n2225 ,n1854 ,n2057);
    or g877(n2224 ,n1822 ,n2066);
    or g878(n2223 ,n1878 ,n2028);
    or g879(n2222 ,n1957 ,n2026);
    or g880(n2221 ,n1908 ,n2118);
    or g881(n2220 ,n1925 ,n2025);
    or g882(n2219 ,n1933 ,n2024);
    or g883(n2218 ,n1952 ,n2023);
    or g884(n2217 ,n1788 ,n2002);
    or g885(n2216 ,n1813 ,n2020);
    or g886(n2215 ,n1815 ,n2021);
    or g887(n2214 ,n1896 ,n2022);
    or g888(n2213 ,n1811 ,n2019);
    or g889(n2212 ,n1810 ,n2018);
    or g890(n2211 ,n1809 ,n2017);
    or g891(n2210 ,n1808 ,n2016);
    or g892(n2209 ,n1806 ,n2015);
    or g893(n2208 ,n1805 ,n2014);
    or g894(n2207 ,n1803 ,n2013);
    or g895(n2206 ,n1802 ,n2012);
    or g896(n2205 ,n1801 ,n2011);
    or g897(n2204 ,n1800 ,n2010);
    or g898(n2203 ,n1798 ,n2007);
    or g899(n2202 ,n1797 ,n2055);
    or g900(n2201 ,n1799 ,n2008);
    or g901(n2200 ,n1796 ,n2005);
    or g902(n2199 ,n1795 ,n2004);
    or g903(n2198 ,n1793 ,n2003);
    or g904(n2197 ,n1792 ,n2001);
    or g905(n2196 ,n1790 ,n1999);
    or g906(n2195 ,n1791 ,n2000);
    or g907(n2194 ,n1789 ,n1998);
    or g908(n2193 ,n1787 ,n1997);
    or g909(n2192 ,n1785 ,n1996);
    or g910(n2191 ,n1784 ,n1995);
    or g911(n2190 ,n1783 ,n1991);
    or g912(n2189 ,n1782 ,n1994);
    or g913(n2188 ,n1781 ,n1993);
    or g914(n2187 ,n1780 ,n1992);
    or g915(n2186 ,n1779 ,n1990);
    or g916(n2185 ,n1776 ,n1989);
    or g917(n2184 ,n1777 ,n1988);
    or g918(n2183 ,n1775 ,n1987);
    or g919(n2182 ,n1772 ,n1984);
    or g920(n2181 ,n1774 ,n1986);
    or g921(n2180 ,n1773 ,n1985);
    or g922(n2179 ,n1771 ,n1983);
    or g923(n2178 ,n1770 ,n1982);
    or g924(n2177 ,n1744 ,n2009);
    or g925(n2176 ,n1768 ,n1980);
    or g926(n2175 ,n1769 ,n1981);
    or g927(n2174 ,n1767 ,n1979);
    or g928(n2173 ,n1766 ,n1977);
    or g929(n2172 ,n1765 ,n1976);
    or g930(n2171 ,n1763 ,n1975);
    or g931(n2170 ,n1761 ,n1974);
    or g932(n2169 ,n1759 ,n1972);
    or g933(n2168 ,n1760 ,n1973);
    or g934(n2167 ,n1762 ,n1978);
    or g935(n2166 ,n1829 ,n1971);
    or g936(n2165 ,n1758 ,n1970);
    or g937(n2164 ,n1757 ,n1969);
    or g938(n2163 ,n1755 ,n1968);
    or g939(n2162 ,n1756 ,n1967);
    or g940(n2161 ,n1754 ,n1966);
    or g941(n2160 ,n1753 ,n1965);
    or g942(n2159 ,n1750 ,n1963);
    or g943(n2158 ,n1751 ,n1964);
    or g944(n2157 ,n1749 ,n1962);
    or g945(n2156 ,n1875 ,n2074);
    nor g946(n2154 ,n1683 ,n1849);
    nor g947(n2153 ,n1733 ,n1836);
    nor g948(n2152 ,n1732 ,n1838);
    nor g949(n2151 ,n1673 ,n1834);
    nor g950(n2150 ,n1728 ,n1849);
    nor g951(n2149 ,n1724 ,n1837);
    nor g952(n2148 ,n1727 ,n1848);
    nor g953(n2147 ,n1726 ,n1847);
    nor g954(n2146 ,n1685 ,n1846);
    nor g955(n2145 ,n1723 ,n1845);
    nor g956(n2144 ,n1721 ,n1844);
    nor g957(n2143 ,n1718 ,n1838);
    nor g958(n2142 ,n1719 ,n1843);
    nor g959(n2141 ,n1702 ,n1842);
    nor g960(n2140 ,n1710 ,n1841);
    nor g961(n2139 ,n1716 ,n1834);
    nor g962(n2138 ,n1720 ,n1840);
    nor g963(n2137 ,n1715 ,n1839);
    nor g964(n2136 ,n1713 ,n1835);
    nor g965(n2135 ,n1712 ,n1849);
    nor g966(n2134 ,n1558 ,n1836);
    nor g967(n2133 ,n1711 ,n1837);
    nor g968(n2132 ,n1709 ,n1838);
    nor g969(n2131 ,n1554 ,n1834);
    nor g970(n2130 ,n1707 ,n1848);
    nor g971(n2129 ,n1599 ,n1849);
    nor g972(n2128 ,n1706 ,n1848);
    nor g973(n2127 ,n1704 ,n1847);
    nor g974(n2126 ,n1703 ,n1846);
    nor g975(n2125 ,n1581 ,n1847);
    nor g976(n2124 ,n1701 ,n1845);
    nor g977(n2123 ,n1698 ,n1846);
    nor g978(n2122 ,n1699 ,n1844);
    nor g979(n2121 ,n1696 ,n1843);
    nor g980(n2120 ,n1635 ,n1845);
    nor g981(n2119 ,n1604 ,n1842);
    nor g982(n2118 ,n1730 ,n1842);
    nor g983(n2117 ,n1695 ,n1841);
    nor g984(n2116 ,n1691 ,n1844);
    nor g985(n2115 ,n1596 ,n1840);
    nor g986(n2114 ,n1690 ,n1839);
    nor g987(n2113 ,n1741 ,n1843);
    nor g988(n2112 ,n1689 ,n1835);
    nor g989(n2111 ,n1657 ,n1836);
    nor g990(n2110 ,n1687 ,n1837);
    nor g991(n2109 ,n1648 ,n1842);
    nor g992(n2108 ,n1684 ,n1841);
    nor g993(n2107 ,n1686 ,n1838);
    nor g994(n2106 ,n1653 ,n1834);
    nor g995(n2105 ,n1547 ,n1834);
    nor g996(n2104 ,n1677 ,n1844);
    nor g997(n2103 ,n1682 ,n1848);
    nor g998(n2102 ,n1662 ,n1847);
    nor g999(n2101 ,n1669 ,n1840);
    nor g1000(n2100 ,n1665 ,n1846);
    nor g1001(n2099 ,n1639 ,n1839);
    nor g1002(n2098 ,n1681 ,n1845);
    nor g1003(n2097 ,n1679 ,n1844);
    nor g1004(n2096 ,n1680 ,n1835);
    nor g1005(n2095 ,n1678 ,n1843);
    nor g1006(n2094 ,n1654 ,n1836);
    nor g1007(n2093 ,n1675 ,n1842);
    nor g1008(n2092 ,n1692 ,n1841);
    nor g1009(n2091 ,n1731 ,n1840);
    nor g1010(n2090 ,n1660 ,n1839);
    nor g1011(n2089 ,n1676 ,n1837);
    nor g1012(n2088 ,n1688 ,n1835);
    nor g1013(n2087 ,n1705 ,n1836);
    nor g1014(n2086 ,n1644 ,n1838);
    nor g1015(n2085 ,n1697 ,n1837);
    nor g1016(n2084 ,n1700 ,n1834);
    nor g1017(n2083 ,n1552 ,n1838);
    nor g1018(n2082 ,n1672 ,n1849);
    nor g1019(n2081 ,n1708 ,n1834);
    nor g1020(n2080 ,n1632 ,n1845);
    nor g1021(n2079 ,n1671 ,n1849);
    nor g1022(n2078 ,n1622 ,n1847);
    nor g1023(n2077 ,n1670 ,n1848);
    nor g1024(n2076 ,n1725 ,n1847);
    nor g1025(n2075 ,n1623 ,n1846);
    nor g1026(n2074 ,n1666 ,n1845);
    nor g1027(n2073 ,n1629 ,n1846);
    nor g1028(n2072 ,n1627 ,n1844);
    nor g1029(n2071 ,n1630 ,n1843);
    nor g1030(n2070 ,n1667 ,n1848);
    nor g1031(n2069 ,n1664 ,n1845);
    nor g1032(n2068 ,n1631 ,n1842);
    nor g1033(n2067 ,n1668 ,n1841);
    nor g1034(n2066 ,n1625 ,n1847);
    nor g1035(n2065 ,n1619 ,n1839);
    nor g1036(n2064 ,n1663 ,n1844);
    nor g1037(n2063 ,n1633 ,n1843);
    nor g1038(n2062 ,n1628 ,n1835);
    nor g1039(n2061 ,n1637 ,n1836);
    nor g1040(n2060 ,n1614 ,n1837);
    nor g1041(n2059 ,n1574 ,n1842);
    nor g1042(n2058 ,n1573 ,n1838);
    nor g1043(n2057 ,n1640 ,n1848);
    or g1044(n2155 ,n1 ,n1851);
    nor g1045(n2055 ,n1592 ,n1839);
    nor g1046(n2054 ,n1656 ,n1841);
    nor g1047(n2053 ,n1655 ,n1848);
    nor g1048(n2052 ,n1582 ,n1847);
    nor g1049(n2051 ,n1563 ,n1840);
    nor g1050(n2050 ,n1568 ,n1846);
    nor g1051(n2049 ,n1571 ,n1839);
    nor g1052(n2048 ,n1652 ,n1845);
    nor g1053(n2047 ,n1584 ,n1844);
    nor g1054(n2046 ,n1594 ,n1843);
    nor g1055(n2045 ,n1651 ,n1835);
    nor g1056(n2044 ,n1610 ,n1836);
    nor g1057(n2043 ,n1600 ,n1842);
    nor g1058(n2042 ,n1612 ,n1841);
    nor g1059(n2041 ,n1634 ,n1840);
    nor g1060(n2040 ,n1620 ,n1839);
    nor g1061(n2039 ,n1647 ,n1837);
    nor g1062(n2038 ,n1645 ,n1835);
    nor g1063(n2037 ,n1642 ,n1834);
    nor g1064(n2036 ,n1638 ,n1836);
    nor g1065(n2035 ,n1643 ,n1837);
    nor g1066(n2034 ,n1717 ,n1838);
    nor g1067(n2033 ,n1650 ,n1838);
    nor g1068(n2032 ,n1608 ,n1849);
    nor g1069(n2031 ,n1624 ,n1834);
    nor g1070(n2030 ,n1658 ,n1849);
    nor g1071(n2029 ,n1557 ,n1848);
    nor g1072(n2028 ,n1674 ,n1846);
    nor g1073(n2027 ,n1626 ,n1840);
    nor g1074(n2026 ,n1694 ,n1843);
    nor g1075(n2025 ,n1714 ,n1841);
    nor g1076(n2024 ,n1722 ,n1840);
    nor g1077(n2023 ,n1729 ,n1839);
    nor g1078(n2022 ,n1616 ,n1836);
    nor g1079(n2021 ,n1617 ,n1835);
    nor g1080(n2020 ,n1615 ,n1837);
    nor g1081(n2019 ,n1613 ,n1838);
    nor g1082(n2018 ,n1611 ,n1834);
    nor g1083(n2017 ,n1609 ,n1849);
    nor g1084(n2016 ,n1607 ,n1848);
    nor g1085(n2015 ,n1605 ,n1847);
    nor g1086(n2014 ,n1603 ,n1846);
    nor g1087(n2013 ,n1602 ,n1845);
    nor g1088(n2012 ,n1601 ,n1844);
    nor g1089(n2011 ,n1598 ,n1843);
    nor g1090(n2010 ,n1597 ,n1842);
    nor g1091(n2009 ,n1588 ,n1847);
    nor g1092(n2008 ,n1595 ,n1841);
    nor g1093(n2007 ,n1593 ,n1840);
    nor g1094(n2006 ,n1559 ,n1849);
    nor g1095(n2005 ,n1591 ,n1835);
    nor g1096(n2004 ,n1590 ,n1836);
    nor g1097(n2003 ,n1589 ,n1837);
    nor g1098(n2002 ,n1578 ,n1846);
    nor g1099(n2001 ,n1587 ,n1838);
    nor g1100(n2000 ,n1586 ,n1834);
    nor g1101(n1999 ,n1585 ,n1849);
    nor g1102(n1998 ,n1583 ,n1848);
    nor g1103(n1997 ,n1580 ,n1847);
    nor g1104(n1996 ,n1579 ,n1846);
    nor g1105(n1995 ,n1576 ,n1845);
    nor g1106(n1994 ,n1575 ,n1844);
    nor g1107(n1993 ,n1544 ,n1843);
    nor g1108(n1992 ,n1549 ,n1842);
    nor g1109(n1991 ,n1572 ,n1845);
    nor g1110(n1990 ,n1553 ,n1841);
    nor g1111(n1989 ,n1569 ,n1844);
    nor g1112(n1988 ,n1570 ,n1840);
    nor g1113(n1987 ,n1566 ,n1839);
    nor g1114(n1986 ,n1567 ,n1835);
    nor g1115(n1985 ,n1565 ,n1836);
    nor g1116(n1984 ,n1564 ,n1843);
    nor g1117(n1983 ,n1577 ,n1837);
    nor g1118(n1982 ,n1562 ,n1838);
    nor g1119(n1981 ,n1561 ,n1834);
    nor g1120(n1980 ,n1560 ,n1842);
    nor g1121(n1979 ,n1606 ,n1849);
    nor g1122(n1978 ,n1636 ,n1841);
    nor g1123(n1977 ,n1618 ,n1848);
    nor g1124(n1976 ,n1621 ,n1847);
    nor g1125(n1975 ,n1641 ,n1846);
    nor g1126(n1974 ,n1556 ,n1845);
    nor g1127(n1973 ,n1555 ,n1844);
    nor g1128(n1972 ,n1649 ,n1840);
    nor g1129(n1971 ,n1646 ,n1843);
    nor g1130(n1970 ,n1551 ,n1842);
    nor g1131(n1969 ,n1550 ,n1841);
    nor g1132(n1968 ,n1659 ,n1839);
    nor g1133(n1967 ,n1548 ,n1840);
    nor g1134(n1966 ,n1661 ,n1839);
    nor g1135(n1965 ,n1546 ,n1835);
    nor g1136(n1964 ,n1545 ,n1836);
    nor g1137(n1963 ,n1543 ,n1835);
    nor g1138(n1962 ,n1693 ,n1837);
    nor g1139(n1961 ,n13[0] ,n1747);
    nor g1140(n1960 ,n1 ,n1833);
    nor g1141(n1959 ,n1 ,n1746);
    nor g1142(n1958 ,n1 ,n1745);
    or g1143(n2056 ,n1 ,n1850);
    nor g1144(n1957 ,n1317 ,n1257);
    nor g1145(n1956 ,n1390 ,n1257);
    nor g1146(n1955 ,n1394 ,n1259);
    nor g1147(n1954 ,n1457 ,n1259);
    nor g1148(n1953 ,n1403 ,n1742);
    nor g1149(n1952 ,n1320 ,n1259);
    nor g1150(n1951 ,n1404 ,n1257);
    nor g1151(n1950 ,n1443 ,n1261);
    nor g1152(n1949 ,n1306 ,n1257);
    nor g1153(n1948 ,n1315 ,n1742);
    nor g1154(n1947 ,n1327 ,n1257);
    nor g1155(n1946 ,n1336 ,n1742);
    nor g1156(n1945 ,n1389 ,n1257);
    nor g1157(n1944 ,n1417 ,n1742);
    nor g1158(n1943 ,n1399 ,n1257);
    nor g1159(n1942 ,n1461 ,n1742);
    nor g1160(n1941 ,n1431 ,n1261);
    nor g1161(n1940 ,n1339 ,n1261);
    nor g1162(n1939 ,n1362 ,n1742);
    nor g1163(n1938 ,n1360 ,n1261);
    nor g1164(n1937 ,n1374 ,n1261);
    nor g1165(n1936 ,n1326 ,n1258);
    nor g1166(n1935 ,n1385 ,n1258);
    nor g1167(n1934 ,n1429 ,n1261);
    nor g1168(n1933 ,n1463 ,n1259);
    nor g1169(n1932 ,n1303 ,n1261);
    nor g1170(n1931 ,n1418 ,n1261);
    nor g1171(n1930 ,n1288 ,n1261);
    nor g1172(n1929 ,n1381 ,n1261);
    nor g1173(n1928 ,n1464 ,n1261);
    nor g1174(n1927 ,n1450 ,n1261);
    nor g1175(n1926 ,n1296 ,n1742);
    nor g1176(n1925 ,n1344 ,n1742);
    nor g1177(n1924 ,n1291 ,n1258);
    nor g1178(n1923 ,n1446 ,n1261);
    nor g1179(n1922 ,n1345 ,n1742);
    nor g1180(n1921 ,n1414 ,n1258);
    nor g1181(n1920 ,n1365 ,n1261);
    nor g1182(n1919 ,n1433 ,n1261);
    nor g1183(n1918 ,n1314 ,n1259);
    nor g1184(n1917 ,n1427 ,n1259);
    nor g1185(n1916 ,n1434 ,n1742);
    nor g1186(n1915 ,n1329 ,n1259);
    nor g1187(n1914 ,n1411 ,n1259);
    nor g1188(n1913 ,n1386 ,n1259);
    nor g1189(n1912 ,n1405 ,n1259);
    nor g1190(n1911 ,n1293 ,n1742);
    nor g1191(n1910 ,n1467 ,n1259);
    nor g1192(n1909 ,n1321 ,n1261);
    nor g1193(n1908 ,n1368 ,n1258);
    nor g1194(n1907 ,n1307 ,n1742);
    nor g1195(n1906 ,n1330 ,n1261);
    nor g1196(n1905 ,n1366 ,n1261);
    nor g1197(n1904 ,n1338 ,n1261);
    nor g1198(n1903 ,n1323 ,n1261);
    nor g1199(n1902 ,n1351 ,n1261);
    nor g1200(n1901 ,n1449 ,n1258);
    nor g1201(n1900 ,n1343 ,n1742);
    nor g1202(n1899 ,n1350 ,n1261);
    nor g1203(n1898 ,n1424 ,n1742);
    nor g1204(n1897 ,n1313 ,n1257);
    nor g1205(n1896 ,n1286 ,n1742);
    nor g1206(n1895 ,n1419 ,n1257);
    nor g1207(n1894 ,n1309 ,n1257);
    nor g1208(n1893 ,n1451 ,n1261);
    nor g1209(n1892 ,n1388 ,n1258);
    nor g1210(n1891 ,n1395 ,n1256);
    nor g1211(n1890 ,n1462 ,n1256);
    nor g1212(n1889 ,n1332 ,n1258);
    nor g1213(n1888 ,n1357 ,n1256);
    nor g1214(n1887 ,n1319 ,n1256);
    nor g1215(n1886 ,n1287 ,n1256);
    nor g1216(n1885 ,n1453 ,n1258);
    nor g1217(n1884 ,n1422 ,n1258);
    nor g1218(n1883 ,n1420 ,n1256);
    nor g1219(n1882 ,n1391 ,n1258);
    nor g1220(n1881 ,n1283 ,n1258);
    nor g1221(n1880 ,n1376 ,n1256);
    nor g1222(n1879 ,n1406 ,n1258);
    nor g1223(n1878 ,n1356 ,n1259);
    nor g1224(n1877 ,n1324 ,n1257);
    nor g1225(n1876 ,n1387 ,n1259);
    nor g1226(n1875 ,n1466 ,n1256);
    nor g1227(n1874 ,n1282 ,n1257);
    nor g1228(n1873 ,n1361 ,n1256);
    nor g1229(n1872 ,n1410 ,n1257);
    nor g1230(n1871 ,n1397 ,n1257);
    nor g1231(n1870 ,n1382 ,n1258);
    nor g1232(n1869 ,n1348 ,n1256);
    nor g1233(n1868 ,n1440 ,n1257);
    nor g1234(n1867 ,n1415 ,n1259);
    nor g1235(n1866 ,n1445 ,n1256);
    nor g1236(n1865 ,n1305 ,n1258);
    nor g1237(n1864 ,n1448 ,n1258);
    nor g1238(n1863 ,n1423 ,n1258);
    nor g1239(n1862 ,n1349 ,n1256);
    nor g1240(n1861 ,n1363 ,n1256);
    nor g1241(n1860 ,n1458 ,n1258);
    nor g1242(n1859 ,n1377 ,n1261);
    nor g1243(n1858 ,n1400 ,n1742);
    nor g1244(n1857 ,n1281 ,n1742);
    nor g1245(n1856 ,n1468 ,n1257);
    nor g1246(n1855 ,n1358 ,n1257);
    nor g1247(n1854 ,n1353 ,n1256);
    nor g1248(n1853 ,n1301 ,n1257);
    nor g1249(n1852 ,n1294 ,n1259);
    not g1250(n1851 ,n1850);
    xnor g1251(n1833 ,n1521 ,n12[0]);
    nor g1252(n1832 ,n1398 ,n1259);
    nor g1253(n1831 ,n1342 ,n1259);
    nor g1254(n1830 ,n1396 ,n1742);
    nor g1255(n1829 ,n1364 ,n1261);
    nor g1256(n1828 ,n1373 ,n1257);
    nor g1257(n1827 ,n1370 ,n1261);
    nor g1258(n1826 ,n1347 ,n1261);
    nor g1259(n1825 ,n1421 ,n1742);
    nor g1260(n1824 ,n1331 ,n1742);
    nor g1261(n1823 ,n1413 ,n1259);
    nor g1262(n1822 ,n1444 ,n1259);
    nor g1263(n1821 ,n1289 ,n1742);
    nor g1264(n1820 ,n1393 ,n1259);
    nor g1265(n1819 ,n1300 ,n1259);
    nor g1266(n1818 ,n1432 ,n1261);
    nor g1267(n1817 ,n1383 ,n1742);
    nor g1268(n1816 ,n1340 ,n1261);
    nor g1269(n1815 ,n1469 ,n1259);
    nor g1270(n1814 ,n1335 ,n1258);
    nor g1271(n1813 ,n1308 ,n1261);
    nor g1272(n1812 ,n1302 ,n1742);
    nor g1273(n1811 ,n1341 ,n1742);
    nor g1274(n1810 ,n1470 ,n1257);
    nor g1275(n1809 ,n1384 ,n1261);
    nor g1276(n1808 ,n1447 ,n1261);
    nor g1277(n1807 ,n1392 ,n1259);
    nor g1278(n1806 ,n1459 ,n1257);
    nor g1279(n1805 ,n1298 ,n1257);
    nor g1280(n1804 ,n1279 ,n1256);
    nor g1281(n1803 ,n1426 ,n1258);
    nor g1282(n1802 ,n1337 ,n1258);
    nor g1283(n1801 ,n1452 ,n1258);
    nor g1284(n1800 ,n1454 ,n1258);
    nor g1285(n1799 ,n1402 ,n1258);
    nor g1286(n1798 ,n1354 ,n1257);
    nor g1287(n1797 ,n1346 ,n1258);
    nor g1288(n1796 ,n1430 ,n1258);
    nor g1289(n1795 ,n1465 ,n1256);
    nor g1290(n1794 ,n1299 ,n1258);
    nor g1291(n1793 ,n1416 ,n1261);
    nor g1292(n1792 ,n1378 ,n1256);
    nor g1293(n1791 ,n1285 ,n1256);
    nor g1294(n1790 ,n1428 ,n1257);
    nor g1295(n1789 ,n1437 ,n1259);
    nor g1296(n1788 ,n1297 ,n1742);
    nor g1297(n1787 ,n1290 ,n1257);
    nor g1298(n1786 ,n1439 ,n1742);
    nor g1299(n1785 ,n1379 ,n1259);
    nor g1300(n1784 ,n1408 ,n1259);
    nor g1301(n1783 ,n1380 ,n1259);
    nor g1302(n1782 ,n1367 ,n1258);
    nor g1303(n1781 ,n1441 ,n1261);
    nor g1304(n1780 ,n1412 ,n1261);
    nor g1305(n1779 ,n1435 ,n1257);
    nor g1306(n1778 ,n1401 ,n1259);
    nor g1307(n1777 ,n1334 ,n1259);
    nor g1308(n1776 ,n1460 ,n1257);
    nor g1309(n1775 ,n1436 ,n1256);
    nor g1310(n1774 ,n1371 ,n1257);
    nor g1311(n1773 ,n1318 ,n1258);
    nor g1312(n1772 ,n1455 ,n1256);
    nor g1313(n1771 ,n1407 ,n1256);
    nor g1314(n1770 ,n1409 ,n1256);
    nor g1315(n1769 ,n1355 ,n1256);
    nor g1316(n1768 ,n1375 ,n1742);
    nor g1317(n1767 ,n1352 ,n1261);
    nor g1318(n1766 ,n1292 ,n1742);
    nor g1319(n1765 ,n1312 ,n1742);
    nor g1320(n1764 ,n1322 ,n1742);
    nor g1321(n1763 ,n1425 ,n1261);
    nor g1322(n1762 ,n1372 ,n1742);
    nor g1323(n1761 ,n1316 ,n1257);
    nor g1324(n1760 ,n1438 ,n1257);
    nor g1325(n1759 ,n1304 ,n1259);
    nor g1326(n1758 ,n1284 ,n1256);
    nor g1327(n1757 ,n1278 ,n1742);
    nor g1328(n1756 ,n1280 ,n1261);
    nor g1329(n1755 ,n1328 ,n1261);
    nor g1330(n1754 ,n1295 ,n1259);
    nor g1331(n1753 ,n1359 ,n1258);
    nor g1332(n1752 ,n1369 ,n1258);
    nor g1333(n1751 ,n1325 ,n1261);
    nor g1334(n1750 ,n1333 ,n1259);
    nor g1335(n1749 ,n1456 ,n1258);
    nor g1336(n1748 ,n1442 ,n1257);
    nor g1337(n1747 ,n1737 ,n1736);
    nor g1338(n1746 ,n1738 ,n1735);
    nor g1339(n1745 ,n1739 ,n1740);
    nor g1340(n1744 ,n1518 ,n1257);
    nor g1341(n1850 ,n1500 ,n1734);
    or g1342(n1849 ,n1509 ,n1743);
    or g1343(n1848 ,n1511 ,n1743);
    or g1344(n1847 ,n1516 ,n1743);
    or g1345(n1846 ,n1504 ,n1743);
    or g1346(n1845 ,n1503 ,n1743);
    or g1347(n1844 ,n1502 ,n1743);
    or g1348(n1843 ,n1505 ,n1743);
    or g1349(n1842 ,n1512 ,n1743);
    or g1350(n1841 ,n1507 ,n1743);
    or g1351(n1840 ,n1506 ,n1743);
    or g1352(n1839 ,n1508 ,n1743);
    or g1353(n1838 ,n1513 ,n1743);
    or g1354(n1837 ,n1515 ,n1743);
    or g1355(n1836 ,n1510 ,n1743);
    or g1356(n1835 ,n1517 ,n1743);
    or g1357(n1834 ,n1514 ,n1743);
    not g1358(n1742 ,n1260);
    not g1359(n1259 ,n1260);
    not g1360(n1260 ,n1261);
    not g1361(n1257 ,n1260);
    not g1362(n1256 ,n1260);
    not g1363(n1258 ,n1260);
    nor g1364(n1741 ,n7[20] ,n1533);
    nor g1365(n1740 ,n1311 ,n1520);
    nor g1366(n1739 ,n1490 ,n1521);
    nor g1367(n1738 ,n1488 ,n1521);
    or g1368(n1737 ,n1519 ,n1526);
    or g1369(n1736 ,n1525 ,n1524);
    nor g1370(n1735 ,n1310 ,n1520);
    or g1371(n1734 ,n12[2] ,n1520);
    nor g1372(n1733 ,n7[10] ,n1536);
    nor g1373(n1732 ,n8[44] ,n1539);
    nor g1374(n1731 ,n9[23] ,n1529);
    nor g1375(n1730 ,n7[53] ,n1531);
    nor g1376(n1729 ,n7[56] ,n1537);
    nor g1377(n1728 ,n8[46] ,n1541);
    nor g1378(n1727 ,n8[47] ,n1540);
    nor g1379(n1726 ,n8[48] ,n1534);
    nor g1380(n1725 ,n9[32] ,n1534);
    nor g1381(n1724 ,n7[11] ,n1527);
    nor g1382(n1723 ,n8[50] ,n1530);
    nor g1383(n1722 ,n7[55] ,n1529);
    nor g1384(n1721 ,n8[51] ,n1532);
    nor g1385(n1720 ,n8[55] ,n1529);
    nor g1386(n1719 ,n8[52] ,n1533);
    nor g1387(n1718 ,n7[12] ,n1539);
    nor g1388(n1717 ,n7[44] ,n1539);
    nor g1389(n1716 ,n7[13] ,n1542);
    nor g1390(n1715 ,n8[56] ,n1537);
    nor g1391(n1714 ,n7[54] ,n1535);
    nor g1392(n1713 ,n8[57] ,n1538);
    nor g1393(n1712 ,n7[14] ,n1541);
    nor g1394(n1711 ,n8[59] ,n1527);
    nor g1395(n1710 ,n8[54] ,n1535);
    nor g1396(n1709 ,n8[60] ,n1539);
    nor g1397(n1708 ,n9[29] ,n1542);
    nor g1398(n1707 ,n7[15] ,n1540);
    nor g1399(n1706 ,n8[63] ,n1540);
    nor g1400(n1705 ,n9[26] ,n1536);
    nor g1401(n1704 ,n9[0] ,n1534);
    nor g1402(n1703 ,n9[1] ,n1528);
    nor g1403(n1702 ,n8[53] ,n1531);
    nor g1404(n1701 ,n9[2] ,n1530);
    nor g1405(n1700 ,n7[29] ,n1542);
    nor g1406(n1699 ,n9[3] ,n1532);
    nor g1407(n1698 ,n7[17] ,n1528);
    nor g1408(n1697 ,n9[27] ,n1527);
    nor g1409(n1696 ,n9[4] ,n1533);
    nor g1410(n1695 ,n9[6] ,n1535);
    nor g1411(n1694 ,n7[52] ,n1533);
    nor g1412(n1693 ,n8[43] ,n1527);
    nor g1413(n1692 ,n9[22] ,n1535);
    nor g1414(n1691 ,n7[19] ,n1532);
    nor g1415(n1690 ,n9[8] ,n1537);
    nor g1416(n1689 ,n9[9] ,n1538);
    nor g1417(n1688 ,n9[25] ,n1538);
    nor g1418(n1687 ,n9[11] ,n1527);
    nor g1419(n1686 ,n9[12] ,n1539);
    nor g1420(n1685 ,n8[49] ,n1528);
    nor g1421(n1684 ,n7[22] ,n1535);
    nor g1422(n1683 ,n9[14] ,n1541);
    nor g1423(n1682 ,n9[15] ,n1540);
    nor g1424(n1681 ,n9[18] ,n1530);
    nor g1425(n1680 ,n7[25] ,n1538);
    nor g1426(n1679 ,n9[19] ,n1532);
    nor g1427(n1678 ,n9[20] ,n1533);
    nor g1428(n1677 ,n7[51] ,n1532);
    nor g1429(n1676 ,n7[27] ,n1527);
    nor g1430(n1675 ,n9[21] ,n1531);
    nor g1431(n1674 ,n7[49] ,n1528);
    nor g1432(n1673 ,n8[45] ,n1542);
    nor g1433(n1672 ,n7[30] ,n1541);
    nor g1434(n1671 ,n9[30] ,n1541);
    nor g1435(n1670 ,n9[31] ,n1540);
    nor g1436(n1669 ,n7[23] ,n1529);
    nor g1437(n1668 ,n9[38] ,n1535);
    nor g1438(n1667 ,n7[31] ,n1540);
    nor g1439(n1666 ,n9[34] ,n1530);
    nor g1440(n1665 ,n9[17] ,n1528);
    nor g1441(n1664 ,n7[34] ,n1530);
    nor g1442(n1663 ,n7[35] ,n1532);
    nor g1443(n1662 ,n9[16] ,n1534);
    nor g1444(n1661 ,n8[40] ,n1537);
    nor g1445(n1660 ,n9[24] ,n1537);
    nor g1446(n1659 ,n7[8] ,n1537);
    nor g1447(n1658 ,n9[62] ,n1541);
    nor g1448(n1657 ,n9[10] ,n1536);
    nor g1449(n1656 ,n7[38] ,n1535);
    nor g1450(n1655 ,n9[47] ,n1540);
    nor g1451(n1654 ,n7[26] ,n1536);
    nor g1452(n1653 ,n9[13] ,n1542);
    nor g1453(n1652 ,n9[50] ,n1530);
    nor g1454(n1651 ,n7[41] ,n1538);
    nor g1455(n1650 ,n9[60] ,n1539);
    nor g1456(n1649 ,n7[7] ,n1529);
    nor g1457(n1648 ,n7[21] ,n1531);
    nor g1458(n1647 ,n7[43] ,n1527);
    nor g1459(n1646 ,n8[36] ,n1533);
    nor g1460(n1645 ,n9[57] ,n1538);
    nor g1461(n1644 ,n7[28] ,n1539);
    or g1462(n1743 ,n1 ,n1522);
    or g1463(n1261 ,n1 ,n1523);
    nor g1464(n1643 ,n9[59] ,n1527);
    nor g1465(n1642 ,n7[45] ,n1542);
    nor g1466(n1641 ,n8[33] ,n1528);
    nor g1467(n1640 ,n9[63] ,n1540);
    nor g1468(n1639 ,n7[24] ,n1537);
    nor g1469(n1638 ,n9[58] ,n1536);
    nor g1470(n1637 ,n9[42] ,n1536);
    nor g1471(n1636 ,n7[6] ,n1535);
    nor g1472(n1635 ,n7[18] ,n1530);
    nor g1473(n1634 ,n9[55] ,n1529);
    nor g1474(n1633 ,n7[36] ,n1533);
    nor g1475(n1632 ,n7[50] ,n1530);
    nor g1476(n1631 ,n9[37] ,n1531);
    nor g1477(n1630 ,n9[36] ,n1533);
    nor g1478(n1629 ,n7[33] ,n1528);
    nor g1479(n1628 ,n9[41] ,n1538);
    nor g1480(n1627 ,n9[35] ,n1532);
    nor g1481(n1626 ,n9[39] ,n1529);
    nor g1482(n1625 ,n7[48] ,n1534);
    nor g1483(n1624 ,n9[61] ,n1542);
    nor g1484(n1623 ,n9[33] ,n1528);
    nor g1485(n1622 ,n7[32] ,n1534);
    nor g1486(n1621 ,n8[32] ,n1534);
    nor g1487(n1620 ,n9[56] ,n1537);
    nor g1488(n1619 ,n9[40] ,n1537);
    nor g1489(n1618 ,n8[31] ,n1540);
    nor g1490(n1617 ,n7[57] ,n1538);
    nor g1491(n1616 ,n7[58] ,n1536);
    nor g1492(n1615 ,n7[59] ,n1527);
    nor g1493(n1614 ,n9[43] ,n1527);
    nor g1494(n1613 ,n7[60] ,n1539);
    nor g1495(n1612 ,n9[54] ,n1535);
    nor g1496(n1611 ,n7[61] ,n1542);
    nor g1497(n1610 ,n7[42] ,n1536);
    nor g1498(n1609 ,n7[62] ,n1541);
    nor g1499(n1608 ,n7[46] ,n1541);
    nor g1500(n1607 ,n7[63] ,n1540);
    nor g1501(n1606 ,n8[30] ,n1541);
    nor g1502(n1605 ,n8[0] ,n1534);
    nor g1503(n1604 ,n9[5] ,n1531);
    nor g1504(n1603 ,n8[1] ,n1528);
    nor g1505(n1602 ,n8[2] ,n1530);
    nor g1506(n1601 ,n8[3] ,n1532);
    nor g1507(n1600 ,n9[53] ,n1531);
    nor g1508(n1599 ,n8[62] ,n1541);
    nor g1509(n1598 ,n8[4] ,n1533);
    nor g1510(n1597 ,n8[5] ,n1531);
    nor g1511(n1596 ,n9[7] ,n1529);
    nor g1512(n1595 ,n8[6] ,n1535);
    nor g1513(n1594 ,n9[52] ,n1533);
    nor g1514(n1593 ,n8[7] ,n1529);
    nor g1515(n1592 ,n8[8] ,n1537);
    nor g1516(n1591 ,n8[9] ,n1538);
    nor g1517(n1590 ,n8[10] ,n1536);
    nor g1518(n1589 ,n8[11] ,n1527);
    nor g1519(n1588 ,n7[0] ,n1534);
    nor g1520(n1587 ,n8[12] ,n1539);
    nor g1521(n1586 ,n8[13] ,n1542);
    nor g1522(n1585 ,n8[14] ,n1541);
    nor g1523(n1584 ,n9[51] ,n1532);
    nor g1524(n1583 ,n8[15] ,n1540);
    nor g1525(n1582 ,n9[48] ,n1534);
    nor g1526(n1581 ,n7[16] ,n1534);
    nor g1527(n1580 ,n8[16] ,n1534);
    nor g1528(n1579 ,n8[17] ,n1528);
    nor g1529(n1578 ,n7[1] ,n1528);
    nor g1530(n1577 ,n8[27] ,n1527);
    nor g1531(n1576 ,n8[18] ,n1530);
    nor g1532(n1575 ,n8[19] ,n1532);
    nor g1533(n1574 ,n7[37] ,n1531);
    nor g1534(n1573 ,n9[44] ,n1539);
    nor g1535(n1572 ,n7[2] ,n1530);
    nor g1536(n1571 ,n7[40] ,n1537);
    nor g1537(n1570 ,n8[23] ,n1529);
    nor g1538(n1569 ,n7[3] ,n1532);
    nor g1539(n1568 ,n9[49] ,n1528);
    nor g1540(n1567 ,n8[25] ,n1538);
    nor g1541(n1566 ,n8[24] ,n1537);
    nor g1542(n1565 ,n8[26] ,n1536);
    nor g1543(n1564 ,n7[4] ,n1533);
    nor g1544(n1563 ,n7[39] ,n1529);
    nor g1545(n1562 ,n8[28] ,n1539);
    nor g1546(n1561 ,n8[29] ,n1542);
    nor g1547(n1560 ,n7[5] ,n1531);
    nor g1548(n1559 ,n9[46] ,n1541);
    nor g1549(n1558 ,n8[58] ,n1536);
    nor g1550(n1557 ,n7[47] ,n1540);
    nor g1551(n1556 ,n8[34] ,n1530);
    nor g1552(n1555 ,n8[35] ,n1532);
    nor g1553(n1554 ,n8[61] ,n1542);
    nor g1554(n1553 ,n8[22] ,n1535);
    nor g1555(n1552 ,n9[28] ,n1539);
    nor g1556(n1551 ,n8[37] ,n1531);
    nor g1557(n1550 ,n8[38] ,n1535);
    nor g1558(n1549 ,n8[21] ,n1531);
    nor g1559(n1548 ,n8[39] ,n1529);
    nor g1560(n1547 ,n9[45] ,n1542);
    nor g1561(n1546 ,n8[41] ,n1538);
    nor g1562(n1545 ,n8[42] ,n1536);
    nor g1563(n1544 ,n8[20] ,n1533);
    nor g1564(n1543 ,n7[9] ,n1538);
    or g1565(n1526 ,n1498 ,n1495);
    or g1566(n1525 ,n1499 ,n1497);
    or g1567(n1524 ,n1492 ,n1491);
    nor g1568(n1542 ,n1473 ,n1501);
    nor g1569(n1541 ,n1472 ,n1501);
    nor g1570(n1540 ,n1479 ,n1501);
    nor g1571(n1539 ,n1476 ,n1501);
    nor g1572(n1538 ,n1482 ,n1501);
    nor g1573(n1537 ,n1484 ,n1501);
    nor g1574(n1536 ,n1478 ,n1501);
    nor g1575(n1535 ,n1475 ,n1501);
    nor g1576(n1534 ,n1486 ,n1501);
    nor g1577(n1533 ,n1485 ,n1501);
    nor g1578(n1532 ,n1481 ,n1501);
    nor g1579(n1531 ,n1480 ,n1501);
    nor g1580(n1530 ,n1474 ,n1501);
    nor g1581(n1529 ,n1487 ,n1501);
    nor g1582(n1528 ,n1483 ,n1501);
    nor g1583(n1527 ,n1471 ,n1501);
    not g1584(n1523 ,n1522);
    not g1585(n1520 ,n1521);
    or g1586(n1519 ,n1493 ,n1494);
    xnor g1587(n1518 ,n2745 ,n10[48]);
    nor g1588(n1517 ,n10[57] ,n1501);
    nor g1589(n1516 ,n10[48] ,n1501);
    nor g1590(n1515 ,n10[59] ,n1501);
    nor g1591(n1514 ,n10[61] ,n1501);
    nor g1592(n1513 ,n10[60] ,n1501);
    nor g1593(n1512 ,n10[53] ,n1501);
    nor g1594(n1511 ,n10[47] ,n1501);
    nor g1595(n1510 ,n10[58] ,n1501);
    nor g1596(n1509 ,n10[62] ,n1501);
    nor g1597(n1508 ,n10[56] ,n1501);
    nor g1598(n1507 ,n10[54] ,n1501);
    nor g1599(n1506 ,n10[55] ,n1501);
    nor g1600(n1505 ,n10[52] ,n1501);
    nor g1601(n1504 ,n10[49] ,n1501);
    nor g1602(n1503 ,n10[50] ,n1501);
    nor g1603(n1502 ,n10[51] ,n1501);
    nor g1604(n1522 ,n13[1] ,n1501);
    nor g1605(n1521 ,n13[1] ,n1496);
    or g1606(n1500 ,n12[0] ,n12[1]);
    or g1607(n1499 ,n6[8] ,n6[9]);
    or g1608(n1498 ,n6[4] ,n6[5]);
    or g1609(n1497 ,n6[10] ,n6[11]);
    or g1610(n1501 ,n1489 ,n13[2]);
    or g1611(n1495 ,n6[6] ,n6[7]);
    or g1612(n1494 ,n6[2] ,n6[3]);
    or g1613(n1493 ,n6[0] ,n6[1]);
    or g1614(n1492 ,n6[12] ,n6[13]);
    or g1615(n1491 ,n6[14] ,n6[15]);
    or g1616(n1496 ,n13[0] ,n13[2]);
    not g1617(n1490 ,n12[2]);
    not g1618(n1489 ,n13[0]);
    not g1619(n1488 ,n12[1]);
    not g1620(n1487 ,n6[7]);
    not g1621(n1486 ,n6[0]);
    not g1622(n1485 ,n6[4]);
    not g1623(n1484 ,n6[8]);
    not g1624(n1483 ,n6[1]);
    not g1625(n1482 ,n6[9]);
    not g1626(n1481 ,n6[3]);
    not g1627(n1480 ,n6[5]);
    not g1628(n1479 ,n6[15]);
    not g1629(n1478 ,n6[10]);
    not g1630(n1477 ,n13[1]);
    not g1631(n1476 ,n6[12]);
    not g1632(n1475 ,n6[6]);
    not g1633(n1474 ,n6[2]);
    not g1634(n1473 ,n6[13]);
    not g1635(n1472 ,n6[14]);
    not g1636(n1471 ,n6[11]);
    not g1637(n1470 ,n2806);
    not g1638(n1469 ,n2802);
    not g1639(n1468 ,n2537);
    not g1640(n1467 ,n2766);
    not g1641(n1466 ,n2523);
    not g1642(n1465 ,n2627);
    not g1643(n1464 ,n2760);
    not g1644(n1463 ,n2800);
    not g1645(n1462 ,n2507);
    not g1646(n1461 ,n2670);
    not g1647(n1460 ,n2748);
    not g1648(n1459 ,n2617);
    not g1649(n1458 ,n2534);
    not g1650(n1457 ,n2663);
    not g1651(n1456 ,n2660);
    not g1652(n1455 ,n2749);
    not g1653(n1454 ,n2622);
    not g1654(n1453 ,n2773);
    not g1655(n1452 ,n2621);
    not g1656(n1451 ,n2770);
    not g1657(n1450 ,n2679);
    not g1658(n1449 ,n2768);
    not g1659(n1448 ,n2532);
    not g1660(n1447 ,n2808);
    not g1661(n1446 ,n2761);
    not g1662(n1445 ,n2531);
    not g1663(n1444 ,n2793);
    not g1664(n1443 ,n2756);
    not g1665(n1442 ,n2551);
    not g1666(n1441 ,n2637);
    not g1667(n1440 ,n2530);
    not g1668(n1439 ,n2491);
    not g1669(n1438 ,n2652);
    not g1670(n1437 ,n2632);
    not g1671(n1436 ,n2641);
    not g1672(n1435 ,n2639);
    not g1673(n1434 ,n2496);
    not g1674(n1433 ,n2493);
    not g1675(n1432 ,n2791);
    not g1676(n1431 ,n2776);
    not g1677(n1430 ,n2626);
    not g1678(n1429 ,n2675);
    not g1679(n1428 ,n2631);
    not g1680(n1427 ,n2495);
    not g1681(n1426 ,n2619);
    not g1682(n1425 ,n2650);
    not g1683(n1424 ,n2506);
    not g1684(n1423 ,n2504);
    not g1685(n1422 ,n2774);
    not g1686(n1421 ,n2548);
    not g1687(n1420 ,n2516);
    not g1688(n1419 ,n2511);
    not g1689(n1418 ,n2775);
    not g1690(n1417 ,n2757);
    not g1691(n1416 ,n2628);
    not g1692(n1415 ,n2781);
    not g1693(n1414 ,n2492);
    not g1694(n1413 ,n2549);
    not g1695(n1412 ,n2638);
    not g1696(n1411 ,n2497);
    not g1697(n1410 ,n2525);
    not g1698(n1409 ,n2645);
    not g1699(n1408 ,n2635);
    not g1700(n1407 ,n2644);
    not g1701(n1406 ,n2521);
    not g1702(n1405 ,n2765);
    not g1703(n1404 ,n2665);
    not g1704(n1403 ,n2664);
    not g1705(n1402 ,n2623);
    not g1706(n1401 ,n2538);
    not g1707(n1400 ,n2784);
    not g1708(n1399 ,n2669);
    not g1709(n1398 ,n2543);
    not g1710(n1397 ,n2780);
    not g1711(n1396 ,n2544);
    not g1712(n1395 ,n2510);
    not g1713(n1394 ,n2515);
    not g1714(n1393 ,n2779);
    not g1715(n1392 ,n2763);
    not g1716(n1391 ,n2517);
    not g1717(n1390 ,n2662);
    not g1718(n1389 ,n2519);
    not g1719(n1388 ,n2509);
    not g1720(n1387 ,n2777);
    not g1721(n1386 ,n2498);
    not g1722(n1385 ,n2674);
    not g1723(n1384 ,n2807);
    not g1724(n1383 ,n2545);
    not g1725(n1382 ,n2527);
    not g1726(n1381 ,n2678);
    not g1727(n1380 ,n2747);
    not g1728(n1379 ,n2634);
    not g1729(n1378 ,n2629);
    not g1730(n1377 ,n2535);
    not g1731(n1376 ,n2518);
    not g1732(n1375 ,n2750);
    not g1733(n1374 ,n2758);
    not g1734(n1373 ,n2550);
    not g1735(n1372 ,n2751);
    not g1736(n1371 ,n2642);
    not g1737(n1370 ,n2546);
    not g1738(n1369 ,n2676);
    not g1739(n1368 ,n2798);
    not g1740(n1367 ,n2636);
    not g1741(n1366 ,n2502);
    not g1742(n1365 ,n2762);
    not g1743(n1364 ,n2653);
    not g1744(n1363 ,n2783);
    not g1745(n1362 ,n2520);
    not g1746(n1361 ,n2778);
    not g1747(n1360 ,n2672);
    not g1748(n1359 ,n2658);
    not g1749(n1358 ,n2785);
    not g1750(n1357 ,n2512);
    not g1751(n1356 ,n2794);
    not g1752(n1355 ,n2646);
    not g1753(n1354 ,n2624);
    not g1754(n1353 ,n2552);
    not g1755(n1352 ,n2647);
    not g1756(n1351 ,n2513);
    not g1757(n1350 ,n2769);
    not g1758(n1349 ,n2533);
    not g1759(n1348 ,n2528);
    not g1760(n1347 ,n2789);
    not g1761(n1346 ,n2625);
    not g1762(n1345 ,n2490);
    not g1763(n1344 ,n2799);
    not g1764(n1343 ,n2505);
    not g1765(n1342 ,n2788);
    not g1766(n1341 ,n2805);
    not g1767(n1340 ,n2529);
    not g1768(n1339 ,n2671);
    not g1769(n1338 ,n2661);
    not g1770(n1337 ,n2620);
    not g1771(n1336 ,n2668);
    not g1772(n1335 ,n2542);
    not g1773(n1334 ,n2640);
    not g1774(n1333 ,n2754);
    not g1775(n1332 ,n2772);
    not g1776(n1331 ,n2790);
    not g1777(n1330 ,n2767);
    not g1778(n1329 ,n2764);
    not g1779(n1328 ,n2753);
    not g1780(n1327 ,n2667);
    not g1781(n1326 ,n2673);
    not g1782(n1325 ,n2659);
    not g1783(n1324 ,n2522);
    not g1784(n1323 ,n2503);
    not g1785(n1322 ,n2536);
    not g1786(n1321 ,n2500);
    not g1787(n1320 ,n2801);
    not g1788(n1319 ,n2771);
    not g1789(n1318 ,n2643);
    not g1790(n1317 ,n2797);
    not g1791(n1316 ,n2651);
    not g1792(n1315 ,n2755);
    not g1793(n1314 ,n2494);
    not g1794(n1313 ,n2796);
    not g1795(n1312 ,n2649);
    not g1796(n1311 ,n2935);
    not g1797(n1310 ,n2936);
    not g1798(n1309 ,n2508);
    not g1799(n1308 ,n2804);
    not g1800(n1307 ,n2501);
    not g1801(n1306 ,n2666);
    not g1802(n1305 ,n2782);
    not g1803(n1304 ,n2752);
    not g1804(n1303 ,n2759);
    not g1805(n1302 ,n2539);
    not g1806(n1301 ,n2786);
    not g1807(n1300 ,n2526);
    not g1808(n1299 ,n2541);
    not g1809(n1298 ,n2618);
    not g1810(n1297 ,n2746);
    not g1811(n1296 ,n2680);
    not g1812(n1295 ,n2657);
    not g1813(n1294 ,n2540);
    not g1814(n1293 ,n2499);
    not g1815(n1292 ,n2648);
    not g1816(n1291 ,n2489);
    not g1817(n1290 ,n2633);
    not g1818(n1289 ,n2547);
    not g1819(n1288 ,n2677);
    not g1820(n1287 ,n2514);
    not g1821(n1286 ,n2803);
    not g1822(n1285 ,n2630);
    not g1823(n1284 ,n2654);
    not g1824(n1283 ,n2795);
    not g1825(n1282 ,n2524);
    not g1826(n1281 ,n2792);
    not g1827(n1280 ,n2656);
    not g1828(n1279 ,n2787);
    not g1829(n1278 ,n2655);
    not g1830(n1277 ,n10[58]);
    not g1831(n1276 ,n10[52]);
    not g1832(n1275 ,n10[59]);
    not g1833(n1274 ,n10[47]);
    not g1834(n1273 ,n10[55]);
    not g1835(n1272 ,n10[60]);
    not g1836(n1271 ,n10[54]);
    not g1837(n1270 ,n10[49]);
    not g1838(n1269 ,n10[62]);
    not g1839(n1268 ,n10[53]);
    not g1840(n1267 ,n10[50]);
    not g1841(n1266 ,n10[51]);
    not g1842(n1265 ,n10[57]);
    not g1843(n1264 ,n10[56]);
    not g1844(n1263 ,n10[61]);
    not g1845(n1262 ,n10[48]);
    xor g1846(n2680 ,n2744 ,n399);
    nor g1847(n2679 ,n398 ,n399);
    nor g1848(n399 ,n94 ,n397);
    nor g1849(n398 ,n2743 ,n396);
    nor g1850(n2678 ,n395 ,n396);
    not g1851(n397 ,n396);
    nor g1852(n396 ,n55 ,n394);
    nor g1853(n395 ,n2742 ,n393);
    xnor g1854(n2677 ,n2741 ,n392);
    not g1855(n394 ,n393);
    nor g1856(n393 ,n93 ,n392);
    nor g1857(n392 ,n213 ,n391);
    xor g1858(n2676 ,n258 ,n390);
    nor g1859(n391 ,n143 ,n390);
    nor g1860(n390 ,n194 ,n389);
    xor g1861(n2675 ,n264 ,n388);
    nor g1862(n389 ,n102 ,n388);
    nor g1863(n388 ,n181 ,n387);
    xor g1864(n2674 ,n259 ,n386);
    nor g1865(n387 ,n144 ,n386);
    nor g1866(n386 ,n162 ,n385);
    xor g1867(n2673 ,n257 ,n384);
    nor g1868(n385 ,n103 ,n384);
    nor g1869(n384 ,n160 ,n383);
    xor g1870(n2672 ,n255 ,n382);
    nor g1871(n383 ,n107 ,n382);
    nor g1872(n382 ,n182 ,n381);
    xor g1873(n2671 ,n254 ,n380);
    nor g1874(n381 ,n139 ,n380);
    nor g1875(n380 ,n179 ,n379);
    xor g1876(n2670 ,n252 ,n378);
    nor g1877(n379 ,n125 ,n378);
    nor g1878(n378 ,n172 ,n377);
    xor g1879(n2669 ,n251 ,n376);
    nor g1880(n377 ,n123 ,n376);
    nor g1881(n376 ,n158 ,n375);
    xor g1882(n2668 ,n250 ,n374);
    nor g1883(n375 ,n152 ,n374);
    nor g1884(n374 ,n196 ,n373);
    xor g1885(n2667 ,n249 ,n372);
    nor g1886(n373 ,n145 ,n372);
    nor g1887(n372 ,n193 ,n371);
    xor g1888(n2666 ,n248 ,n370);
    nor g1889(n371 ,n104 ,n370);
    nor g1890(n370 ,n200 ,n369);
    xor g1891(n2665 ,n226 ,n368);
    nor g1892(n369 ,n108 ,n368);
    nor g1893(n368 ,n210 ,n367);
    xor g1894(n2664 ,n225 ,n366);
    nor g1895(n367 ,n154 ,n366);
    nor g1896(n366 ,n206 ,n365);
    xor g1897(n2663 ,n224 ,n364);
    nor g1898(n365 ,n131 ,n364);
    nor g1899(n364 ,n203 ,n363);
    xor g1900(n2662 ,n222 ,n362);
    nor g1901(n363 ,n96 ,n362);
    nor g1902(n362 ,n201 ,n361);
    xor g1903(n2661 ,n220 ,n360);
    nor g1904(n361 ,n97 ,n360);
    nor g1905(n360 ,n170 ,n359);
    xor g1906(n2660 ,n246 ,n358);
    nor g1907(n359 ,n101 ,n358);
    nor g1908(n358 ,n165 ,n357);
    xor g1909(n2659 ,n245 ,n356);
    nor g1910(n357 ,n149 ,n356);
    nor g1911(n356 ,n161 ,n355);
    xor g1912(n2658 ,n244 ,n354);
    nor g1913(n355 ,n98 ,n354);
    nor g1914(n354 ,n157 ,n353);
    xor g1915(n2657 ,n243 ,n352);
    nor g1916(n353 ,n113 ,n352);
    nor g1917(n352 ,n155 ,n351);
    xor g1918(n2656 ,n242 ,n350);
    nor g1919(n351 ,n153 ,n350);
    nor g1920(n350 ,n184 ,n349);
    xor g1921(n2655 ,n240 ,n348);
    nor g1922(n349 ,n141 ,n348);
    nor g1923(n348 ,n156 ,n347);
    xor g1924(n2654 ,n239 ,n346);
    nor g1925(n347 ,n132 ,n346);
    nor g1926(n346 ,n192 ,n345);
    xor g1927(n2653 ,n238 ,n344);
    nor g1928(n345 ,n100 ,n344);
    nor g1929(n344 ,n189 ,n343);
    xor g1930(n2652 ,n236 ,n342);
    nor g1931(n343 ,n106 ,n342);
    nor g1932(n342 ,n178 ,n341);
    xor g1933(n2651 ,n235 ,n340);
    nor g1934(n341 ,n119 ,n340);
    nor g1935(n340 ,n197 ,n339);
    xor g1936(n2650 ,n233 ,n338);
    nor g1937(n339 ,n138 ,n338);
    nor g1938(n338 ,n205 ,n337);
    xor g1939(n2649 ,n218 ,n336);
    nor g1940(n337 ,n112 ,n336);
    nor g1941(n336 ,n209 ,n335);
    xor g1942(n2648 ,n217 ,n334);
    nor g1943(n335 ,n137 ,n334);
    nor g1944(n334 ,n208 ,n333);
    xor g1945(n2647 ,n216 ,n332);
    nor g1946(n333 ,n116 ,n332);
    nor g1947(n332 ,n207 ,n331);
    xor g1948(n2646 ,n230 ,n330);
    nor g1949(n331 ,n120 ,n330);
    nor g1950(n330 ,n204 ,n329);
    xor g1951(n2645 ,n229 ,n328);
    nor g1952(n329 ,n127 ,n328);
    nor g1953(n328 ,n180 ,n327);
    xor g1954(n2644 ,n274 ,n326);
    nor g1955(n327 ,n118 ,n326);
    nor g1956(n326 ,n177 ,n325);
    xor g1957(n2643 ,n273 ,n324);
    nor g1958(n325 ,n114 ,n324);
    nor g1959(n324 ,n175 ,n323);
    xor g1960(n2642 ,n272 ,n322);
    nor g1961(n323 ,n147 ,n322);
    nor g1962(n322 ,n174 ,n321);
    xor g1963(n2641 ,n231 ,n320);
    nor g1964(n321 ,n130 ,n320);
    nor g1965(n320 ,n173 ,n319);
    xor g1966(n2640 ,n232 ,n318);
    nor g1967(n319 ,n126 ,n318);
    nor g1968(n318 ,n171 ,n317);
    xor g1969(n2639 ,n234 ,n316);
    nor g1970(n317 ,n133 ,n316);
    nor g1971(n316 ,n169 ,n315);
    xor g1972(n2638 ,n270 ,n314);
    nor g1973(n315 ,n115 ,n314);
    nor g1974(n314 ,n166 ,n313);
    xor g1975(n2637 ,n271 ,n312);
    nor g1976(n313 ,n142 ,n312);
    nor g1977(n312 ,n164 ,n311);
    xor g1978(n2636 ,n241 ,n310);
    nor g1979(n311 ,n150 ,n310);
    nor g1980(n310 ,n163 ,n309);
    xor g1981(n2635 ,n269 ,n308);
    nor g1982(n309 ,n128 ,n308);
    nor g1983(n308 ,n159 ,n307);
    xor g1984(n2634 ,n267 ,n306);
    nor g1985(n307 ,n117 ,n306);
    nor g1986(n306 ,n199 ,n305);
    xor g1987(n2633 ,n219 ,n304);
    nor g1988(n305 ,n124 ,n304);
    nor g1989(n304 ,n211 ,n303);
    xor g1990(n2632 ,n221 ,n302);
    nor g1991(n303 ,n146 ,n302);
    nor g1992(n302 ,n198 ,n301);
    xor g1993(n2631 ,n227 ,n300);
    nor g1994(n301 ,n129 ,n300);
    nor g1995(n300 ,n212 ,n299);
    xor g1996(n2630 ,n228 ,n298);
    nor g1997(n299 ,n121 ,n298);
    nor g1998(n298 ,n202 ,n297);
    xor g1999(n2629 ,n223 ,n296);
    nor g2000(n297 ,n109 ,n296);
    nor g2001(n296 ,n183 ,n295);
    xor g2002(n2628 ,n261 ,n294);
    nor g2003(n295 ,n99 ,n294);
    nor g2004(n294 ,n195 ,n293);
    xor g2005(n2627 ,n247 ,n292);
    nor g2006(n293 ,n148 ,n292);
    nor g2007(n292 ,n168 ,n291);
    xor g2008(n2626 ,n237 ,n290);
    nor g2009(n291 ,n135 ,n290);
    nor g2010(n290 ,n190 ,n289);
    xor g2011(n2625 ,n253 ,n288);
    nor g2012(n289 ,n134 ,n288);
    nor g2013(n288 ,n191 ,n287);
    xor g2014(n2624 ,n265 ,n286);
    nor g2015(n287 ,n95 ,n286);
    nor g2016(n286 ,n167 ,n285);
    xor g2017(n2623 ,n256 ,n284);
    nor g2018(n285 ,n111 ,n284);
    nor g2019(n284 ,n188 ,n283);
    xor g2020(n2622 ,n268 ,n282);
    nor g2021(n283 ,n105 ,n282);
    nor g2022(n282 ,n185 ,n281);
    xor g2023(n2621 ,n266 ,n280);
    nor g2024(n281 ,n151 ,n280);
    nor g2025(n280 ,n186 ,n279);
    xor g2026(n2620 ,n263 ,n278);
    nor g2027(n279 ,n136 ,n278);
    nor g2028(n278 ,n176 ,n277);
    xor g2029(n2619 ,n260 ,n276);
    nor g2030(n277 ,n110 ,n276);
    xnor g2031(n2618 ,n262 ,n214);
    nor g2032(n276 ,n187 ,n275);
    nor g2033(n2617 ,n214 ,n140);
    nor g2034(n275 ,n215 ,n122);
    xnor g2035(n274 ,n11[43] ,n2708);
    xnor g2036(n273 ,n11[42] ,n2707);
    xnor g2037(n272 ,n11[41] ,n2706);
    xnor g2038(n271 ,n11[36] ,n2701);
    xnor g2039(n270 ,n11[37] ,n2702);
    xnor g2040(n269 ,n11[34] ,n2699);
    xnor g2041(n268 ,n11[37] ,n2686);
    xnor g2042(n267 ,n11[33] ,n2698);
    xnor g2043(n266 ,n11[36] ,n2685);
    xnor g2044(n265 ,n11[39] ,n2688);
    xnor g2045(n264 ,n11[42] ,n2739);
    xnor g2046(n263 ,n11[35] ,n2684);
    xnor g2047(n262 ,n11[33] ,n2682);
    xnor g2048(n261 ,n11[43] ,n2692);
    xnor g2049(n260 ,n11[34] ,n2683);
    xnor g2050(n259 ,n11[41] ,n2738);
    xnor g2051(n258 ,n11[43] ,n2740);
    xnor g2052(n257 ,n11[40] ,n2737);
    xnor g2053(n256 ,n11[38] ,n2687);
    xnor g2054(n255 ,n11[39] ,n2736);
    xnor g2055(n254 ,n11[38] ,n2735);
    xnor g2056(n253 ,n11[40] ,n2689);
    xnor g2057(n252 ,n11[37] ,n2734);
    xnor g2058(n251 ,n11[36] ,n2733);
    xnor g2059(n250 ,n11[35] ,n2732);
    xnor g2060(n249 ,n11[34] ,n2731);
    xnor g2061(n248 ,n11[33] ,n2730);
    xnor g2062(n247 ,n11[42] ,n2691);
    xnor g2063(n246 ,n11[43] ,n2724);
    xnor g2064(n245 ,n11[42] ,n2723);
    xnor g2065(n244 ,n11[41] ,n2722);
    xnor g2066(n243 ,n11[40] ,n2721);
    xnor g2067(n242 ,n11[39] ,n2720);
    xnor g2068(n241 ,n11[35] ,n2700);
    xnor g2069(n240 ,n11[38] ,n2719);
    xnor g2070(n239 ,n11[37] ,n2718);
    xnor g2071(n238 ,n11[36] ,n2717);
    xnor g2072(n237 ,n11[41] ,n2690);
    xnor g2073(n236 ,n11[35] ,n2716);
    xnor g2074(n235 ,n11[34] ,n2715);
    xnor g2075(n234 ,n11[38] ,n2703);
    xnor g2076(n233 ,n11[33] ,n2714);
    xnor g2077(n232 ,n11[39] ,n2704);
    xnor g2078(n231 ,n11[40] ,n2705);
    xnor g2079(n230 ,n11[45] ,n2710);
    xnor g2080(n229 ,n11[44] ,n2709);
    xnor g2081(n228 ,n11[45] ,n2694);
    xnor g2082(n227 ,n11[46] ,n2695);
    xnor g2083(n226 ,n11[32] ,n2729);
    xnor g2084(n225 ,n11[31] ,n2728);
    xnor g2085(n224 ,n11[46] ,n2727);
    xnor g2086(n223 ,n11[44] ,n2693);
    xnor g2087(n222 ,n11[45] ,n2726);
    xnor g2088(n221 ,n11[31] ,n2696);
    xnor g2089(n220 ,n11[44] ,n2725);
    xnor g2090(n219 ,n11[32] ,n2697);
    xnor g2091(n218 ,n11[32] ,n2713);
    xnor g2092(n217 ,n11[31] ,n2712);
    xnor g2093(n216 ,n11[46] ,n2711);
    not g2094(n215 ,n214);
    nor g2095(n213 ,n70 ,n60);
    nor g2096(n212 ,n77 ,n21);
    nor g2097(n211 ,n72 ,n19);
    nor g2098(n210 ,n28 ,n19);
    nor g2099(n209 ,n65 ,n19);
    nor g2100(n208 ,n48 ,n64);
    nor g2101(n207 ,n27 ,n21);
    nor g2102(n206 ,n69 ,n64);
    nor g2103(n205 ,n79 ,n20);
    nor g2104(n204 ,n49 ,n63);
    nor g2105(n203 ,n66 ,n21);
    nor g2106(n202 ,n91 ,n63);
    nor g2107(n201 ,n43 ,n63);
    nor g2108(n200 ,n40 ,n20);
    nor g2109(n199 ,n36 ,n20);
    nor g2110(n198 ,n44 ,n64);
    nor g2111(n197 ,n25 ,n57);
    nor g2112(n196 ,n76 ,n59);
    nor g2113(n195 ,n35 ,n56);
    nor g2114(n194 ,n83 ,n56);
    nor g2115(n193 ,n75 ,n57);
    nor g2116(n192 ,n68 ,n58);
    nor g2117(n191 ,n46 ,n16);
    nor g2118(n190 ,n45 ,n62);
    nor g2119(n189 ,n47 ,n61);
    nor g2120(n188 ,n85 ,n18);
    nor g2121(n187 ,n67 ,n57);
    nor g2122(n186 ,n74 ,n61);
    nor g2123(n185 ,n84 ,n58);
    nor g2124(n184 ,n52 ,n15);
    nor g2125(n183 ,n89 ,n60);
    nor g2126(n182 ,n71 ,n15);
    nor g2127(n181 ,n50 ,n17);
    nor g2128(n180 ,n88 ,n60);
    nor g2129(n179 ,n26 ,n18);
    nor g2130(n178 ,n51 ,n59);
    nor g2131(n177 ,n32 ,n56);
    nor g2132(n176 ,n23 ,n59);
    nor g2133(n175 ,n22 ,n17);
    nor g2134(n174 ,n31 ,n62);
    nor g2135(n173 ,n81 ,n16);
    nor g2136(n172 ,n34 ,n58);
    nor g2137(n171 ,n87 ,n15);
    nor g2138(n170 ,n29 ,n60);
    nor g2139(n169 ,n41 ,n18);
    nor g2140(n168 ,n92 ,n17);
    nor g2141(n167 ,n39 ,n15);
    nor g2142(n166 ,n37 ,n58);
    nor g2143(n165 ,n82 ,n56);
    nor g2144(n164 ,n86 ,n61);
    nor g2145(n163 ,n78 ,n59);
    nor g2146(n162 ,n73 ,n62);
    nor g2147(n161 ,n80 ,n17);
    nor g2148(n160 ,n90 ,n16);
    nor g2149(n159 ,n42 ,n57);
    nor g2150(n158 ,n38 ,n61);
    nor g2151(n157 ,n24 ,n62);
    nor g2152(n156 ,n33 ,n18);
    nor g2153(n155 ,n30 ,n16);
    nor g2154(n214 ,n54 ,n53);
    nor g2155(n154 ,n2728 ,n11[31]);
    nor g2156(n153 ,n2720 ,n11[39]);
    nor g2157(n152 ,n2732 ,n11[35]);
    nor g2158(n151 ,n2685 ,n11[36]);
    nor g2159(n150 ,n2700 ,n11[35]);
    nor g2160(n149 ,n2723 ,n11[42]);
    nor g2161(n148 ,n2691 ,n11[42]);
    nor g2162(n147 ,n2706 ,n11[41]);
    nor g2163(n146 ,n2696 ,n11[31]);
    nor g2164(n145 ,n2731 ,n11[34]);
    nor g2165(n144 ,n2738 ,n11[41]);
    nor g2166(n143 ,n2740 ,n11[43]);
    nor g2167(n142 ,n2701 ,n11[36]);
    nor g2168(n141 ,n2719 ,n11[38]);
    nor g2169(n140 ,n2681 ,n10[49]);
    nor g2170(n139 ,n2735 ,n11[38]);
    nor g2171(n138 ,n2714 ,n11[33]);
    nor g2172(n137 ,n2712 ,n11[31]);
    nor g2173(n136 ,n2684 ,n11[35]);
    nor g2174(n135 ,n2690 ,n11[41]);
    nor g2175(n134 ,n2689 ,n11[40]);
    nor g2176(n133 ,n2703 ,n11[38]);
    nor g2177(n132 ,n2718 ,n11[37]);
    nor g2178(n131 ,n2727 ,n11[46]);
    nor g2179(n130 ,n2705 ,n11[40]);
    nor g2180(n129 ,n2695 ,n11[46]);
    nor g2181(n128 ,n2699 ,n11[34]);
    nor g2182(n127 ,n2709 ,n11[44]);
    nor g2183(n126 ,n2704 ,n11[39]);
    nor g2184(n125 ,n2734 ,n11[37]);
    nor g2185(n124 ,n2697 ,n11[32]);
    nor g2186(n123 ,n2733 ,n11[36]);
    nor g2187(n122 ,n2682 ,n11[33]);
    nor g2188(n121 ,n2694 ,n11[45]);
    nor g2189(n120 ,n2710 ,n11[45]);
    nor g2190(n119 ,n2715 ,n11[34]);
    nor g2191(n118 ,n2708 ,n11[43]);
    nor g2192(n117 ,n2698 ,n11[33]);
    nor g2193(n116 ,n2711 ,n11[46]);
    nor g2194(n115 ,n2702 ,n11[37]);
    nor g2195(n114 ,n2707 ,n11[42]);
    nor g2196(n113 ,n2721 ,n11[40]);
    nor g2197(n112 ,n2713 ,n11[32]);
    nor g2198(n111 ,n2687 ,n11[38]);
    nor g2199(n110 ,n2683 ,n11[34]);
    nor g2200(n109 ,n2693 ,n11[44]);
    nor g2201(n108 ,n2729 ,n11[32]);
    nor g2202(n107 ,n2736 ,n11[39]);
    nor g2203(n106 ,n2716 ,n11[35]);
    nor g2204(n105 ,n2686 ,n11[37]);
    nor g2205(n104 ,n2730 ,n11[33]);
    nor g2206(n103 ,n2737 ,n11[40]);
    nor g2207(n102 ,n2739 ,n11[42]);
    nor g2208(n101 ,n2724 ,n11[43]);
    nor g2209(n100 ,n2717 ,n11[36]);
    nor g2210(n99 ,n2692 ,n11[43]);
    nor g2211(n98 ,n2722 ,n11[41]);
    nor g2212(n97 ,n2725 ,n11[44]);
    nor g2213(n96 ,n2726 ,n11[45]);
    nor g2214(n95 ,n2688 ,n11[39]);
    not g2215(n94 ,n2743);
    not g2216(n93 ,n2741);
    not g2217(n92 ,n2690);
    not g2218(n91 ,n2693);
    not g2219(n90 ,n2736);
    not g2220(n89 ,n2692);
    not g2221(n88 ,n2708);
    not g2222(n87 ,n2703);
    not g2223(n86 ,n2700);
    not g2224(n85 ,n2686);
    not g2225(n84 ,n2685);
    not g2226(n83 ,n2739);
    not g2227(n82 ,n2723);
    not g2228(n81 ,n2704);
    not g2229(n80 ,n2722);
    not g2230(n79 ,n2713);
    not g2231(n78 ,n2699);
    not g2232(n77 ,n2694);
    not g2233(n76 ,n2731);
    not g2234(n75 ,n2730);
    not g2235(n74 ,n2684);
    not g2236(n73 ,n2737);
    not g2237(n72 ,n2696);
    not g2238(n71 ,n2735);
    not g2239(n70 ,n2740);
    not g2240(n69 ,n2727);
    not g2241(n68 ,n2717);
    not g2242(n67 ,n2682);
    not g2243(n66 ,n2726);
    not g2244(n65 ,n2712);
    not g2245(n64 ,n11[46]);
    not g2246(n63 ,n11[44]);
    not g2247(n62 ,n11[40]);
    not g2248(n61 ,n11[35]);
    not g2249(n60 ,n11[43]);
    not g2250(n59 ,n11[34]);
    not g2251(n58 ,n11[36]);
    not g2252(n57 ,n11[33]);
    not g2253(n56 ,n11[42]);
    not g2254(n55 ,n2742);
    not g2255(n54 ,n2681);
    not g2256(n53 ,n10[49]);
    not g2257(n52 ,n2719);
    not g2258(n51 ,n2715);
    not g2259(n50 ,n2738);
    not g2260(n49 ,n2709);
    not g2261(n48 ,n2711);
    not g2262(n47 ,n2716);
    not g2263(n46 ,n2688);
    not g2264(n45 ,n2689);
    not g2265(n44 ,n2695);
    not g2266(n43 ,n2725);
    not g2267(n42 ,n2698);
    not g2268(n41 ,n2702);
    not g2269(n40 ,n2729);
    not g2270(n39 ,n2687);
    not g2271(n38 ,n2732);
    not g2272(n37 ,n2701);
    not g2273(n36 ,n2697);
    not g2274(n35 ,n2691);
    not g2275(n34 ,n2733);
    not g2276(n33 ,n2718);
    not g2277(n32 ,n2707);
    not g2278(n31 ,n2705);
    not g2279(n30 ,n2720);
    not g2280(n29 ,n2724);
    not g2281(n28 ,n2728);
    not g2282(n27 ,n2710);
    not g2283(n26 ,n2734);
    not g2284(n25 ,n2714);
    not g2285(n24 ,n2721);
    not g2286(n23 ,n2683);
    not g2287(n22 ,n2706);
    not g2288(n21 ,n11[45]);
    not g2289(n20 ,n11[32]);
    not g2290(n19 ,n11[31]);
    not g2291(n18 ,n11[37]);
    not g2292(n17 ,n11[41]);
    not g2293(n16 ,n11[39]);
    not g2294(n15 ,n11[38]);
    xnor g2295(n2552 ,n2616 ,n729);
    nor g2296(n729 ,n526 ,n728);
    xor g2297(n2551 ,n593 ,n727);
    nor g2298(n728 ,n593 ,n727);
    nor g2299(n727 ,n484 ,n726);
    xor g2300(n2550 ,n603 ,n725);
    nor g2301(n726 ,n603 ,n725);
    nor g2302(n725 ,n517 ,n724);
    xor g2303(n2549 ,n565 ,n723);
    nor g2304(n724 ,n565 ,n723);
    nor g2305(n723 ,n493 ,n722);
    xor g2306(n2548 ,n590 ,n721);
    nor g2307(n722 ,n590 ,n721);
    nor g2308(n721 ,n530 ,n720);
    xor g2309(n2547 ,n587 ,n719);
    nor g2310(n720 ,n587 ,n719);
    nor g2311(n719 ,n490 ,n718);
    xor g2312(n2546 ,n569 ,n717);
    nor g2313(n718 ,n569 ,n717);
    nor g2314(n717 ,n497 ,n716);
    xor g2315(n2545 ,n554 ,n715);
    nor g2316(n716 ,n554 ,n715);
    nor g2317(n715 ,n485 ,n714);
    xor g2318(n2544 ,n575 ,n713);
    nor g2319(n714 ,n575 ,n713);
    nor g2320(n713 ,n482 ,n712);
    xor g2321(n2543 ,n604 ,n711);
    nor g2322(n712 ,n604 ,n711);
    nor g2323(n711 ,n527 ,n710);
    xor g2324(n2542 ,n592 ,n709);
    nor g2325(n710 ,n592 ,n709);
    nor g2326(n709 ,n519 ,n708);
    xor g2327(n2541 ,n579 ,n707);
    nor g2328(n708 ,n579 ,n707);
    nor g2329(n707 ,n491 ,n706);
    xor g2330(n2540 ,n570 ,n705);
    nor g2331(n706 ,n570 ,n705);
    nor g2332(n705 ,n504 ,n704);
    xor g2333(n2539 ,n564 ,n703);
    nor g2334(n704 ,n564 ,n703);
    nor g2335(n703 ,n489 ,n702);
    xor g2336(n2538 ,n555 ,n701);
    nor g2337(n702 ,n555 ,n701);
    nor g2338(n701 ,n483 ,n700);
    xor g2339(n2537 ,n551 ,n699);
    nor g2340(n700 ,n551 ,n699);
    nor g2341(n699 ,n536 ,n698);
    xor g2342(n2536 ,n544 ,n697);
    nor g2343(n698 ,n544 ,n697);
    nor g2344(n697 ,n541 ,n696);
    xor g2345(n2535 ,n559 ,n695);
    nor g2346(n696 ,n559 ,n695);
    nor g2347(n695 ,n492 ,n694);
    xor g2348(n2534 ,n556 ,n693);
    nor g2349(n694 ,n556 ,n693);
    nor g2350(n693 ,n533 ,n692);
    xor g2351(n2533 ,n601 ,n691);
    nor g2352(n692 ,n601 ,n691);
    nor g2353(n691 ,n534 ,n690);
    xor g2354(n2532 ,n597 ,n689);
    nor g2355(n690 ,n597 ,n689);
    nor g2356(n689 ,n542 ,n688);
    xor g2357(n2531 ,n589 ,n687);
    nor g2358(n688 ,n589 ,n687);
    nor g2359(n687 ,n521 ,n686);
    xor g2360(n2530 ,n585 ,n685);
    nor g2361(n686 ,n585 ,n685);
    nor g2362(n685 ,n518 ,n684);
    xor g2363(n2529 ,n580 ,n683);
    nor g2364(n684 ,n580 ,n683);
    nor g2365(n683 ,n479 ,n682);
    xor g2366(n2528 ,n576 ,n681);
    nor g2367(n682 ,n576 ,n681);
    nor g2368(n681 ,n512 ,n680);
    xor g2369(n2527 ,n573 ,n679);
    nor g2370(n680 ,n573 ,n679);
    nor g2371(n679 ,n507 ,n678);
    xor g2372(n2526 ,n545 ,n677);
    nor g2373(n678 ,n545 ,n677);
    nor g2374(n677 ,n503 ,n676);
    xor g2375(n2525 ,n567 ,n675);
    nor g2376(n676 ,n567 ,n675);
    nor g2377(n675 ,n500 ,n674);
    xor g2378(n2524 ,n563 ,n673);
    nor g2379(n674 ,n563 ,n673);
    nor g2380(n673 ,n488 ,n672);
    xor g2381(n2523 ,n561 ,n671);
    nor g2382(n672 ,n561 ,n671);
    nor g2383(n671 ,n496 ,n670);
    xor g2384(n2522 ,n557 ,n669);
    nor g2385(n670 ,n557 ,n669);
    nor g2386(n669 ,n487 ,n668);
    xor g2387(n2521 ,n547 ,n667);
    nor g2388(n668 ,n547 ,n667);
    nor g2389(n667 ,n538 ,n666);
    xor g2390(n2520 ,n577 ,n665);
    nor g2391(n666 ,n577 ,n665);
    nor g2392(n665 ,n537 ,n664);
    xor g2393(n2519 ,n582 ,n663);
    nor g2394(n664 ,n582 ,n663);
    nor g2395(n663 ,n522 ,n662);
    xor g2396(n2518 ,n595 ,n661);
    nor g2397(n662 ,n595 ,n661);
    nor g2398(n661 ,n480 ,n660);
    xor g2399(n2517 ,n548 ,n659);
    nor g2400(n660 ,n548 ,n659);
    nor g2401(n659 ,n486 ,n658);
    xor g2402(n2516 ,n549 ,n657);
    nor g2403(n658 ,n549 ,n657);
    nor g2404(n657 ,n513 ,n656);
    xor g2405(n2515 ,n552 ,n655);
    nor g2406(n656 ,n552 ,n655);
    nor g2407(n655 ,n494 ,n654);
    xor g2408(n2514 ,n553 ,n653);
    nor g2409(n654 ,n553 ,n653);
    nor g2410(n653 ,n535 ,n652);
    xor g2411(n2513 ,n550 ,n651);
    nor g2412(n652 ,n550 ,n651);
    nor g2413(n651 ,n495 ,n650);
    xor g2414(n2512 ,n574 ,n649);
    nor g2415(n650 ,n574 ,n649);
    nor g2416(n649 ,n532 ,n648);
    xor g2417(n2511 ,n602 ,n647);
    nor g2418(n648 ,n602 ,n647);
    nor g2419(n647 ,n531 ,n646);
    xor g2420(n2510 ,n599 ,n645);
    nor g2421(n646 ,n599 ,n645);
    nor g2422(n645 ,n529 ,n644);
    xor g2423(n2509 ,n596 ,n643);
    nor g2424(n644 ,n596 ,n643);
    nor g2425(n643 ,n528 ,n642);
    xor g2426(n2508 ,n594 ,n641);
    nor g2427(n642 ,n594 ,n641);
    nor g2428(n641 ,n525 ,n640);
    xor g2429(n2507 ,n591 ,n639);
    nor g2430(n640 ,n591 ,n639);
    nor g2431(n639 ,n523 ,n638);
    xor g2432(n2506 ,n588 ,n637);
    nor g2433(n638 ,n588 ,n637);
    nor g2434(n637 ,n520 ,n636);
    xor g2435(n2505 ,n586 ,n635);
    nor g2436(n636 ,n586 ,n635);
    nor g2437(n635 ,n540 ,n634);
    xor g2438(n2504 ,n583 ,n633);
    nor g2439(n634 ,n583 ,n633);
    nor g2440(n633 ,n539 ,n632);
    xor g2441(n2503 ,n581 ,n631);
    nor g2442(n632 ,n581 ,n631);
    nor g2443(n631 ,n516 ,n630);
    xor g2444(n2502 ,n578 ,n629);
    nor g2445(n630 ,n578 ,n629);
    nor g2446(n629 ,n515 ,n628);
    xor g2447(n2501 ,n584 ,n627);
    nor g2448(n628 ,n584 ,n627);
    nor g2449(n627 ,n514 ,n626);
    xor g2450(n2500 ,n558 ,n625);
    nor g2451(n626 ,n558 ,n625);
    nor g2452(n625 ,n511 ,n624);
    xor g2453(n2499 ,n572 ,n623);
    nor g2454(n624 ,n572 ,n623);
    nor g2455(n623 ,n508 ,n622);
    xor g2456(n2498 ,n571 ,n621);
    nor g2457(n622 ,n571 ,n621);
    nor g2458(n621 ,n506 ,n620);
    xor g2459(n2497 ,n598 ,n619);
    nor g2460(n620 ,n598 ,n619);
    nor g2461(n619 ,n505 ,n618);
    xor g2462(n2496 ,n568 ,n617);
    nor g2463(n618 ,n568 ,n617);
    nor g2464(n617 ,n502 ,n616);
    xor g2465(n2495 ,n600 ,n615);
    nor g2466(n616 ,n600 ,n615);
    nor g2467(n615 ,n501 ,n614);
    xor g2468(n2494 ,n566 ,n613);
    nor g2469(n614 ,n566 ,n613);
    nor g2470(n613 ,n499 ,n612);
    xor g2471(n2493 ,n546 ,n611);
    nor g2472(n612 ,n546 ,n611);
    nor g2473(n611 ,n498 ,n610);
    xor g2474(n2492 ,n562 ,n609);
    nor g2475(n610 ,n562 ,n609);
    nor g2476(n609 ,n524 ,n608);
    xnor g2477(n2491 ,n560 ,n606);
    nor g2478(n608 ,n560 ,n607);
    not g2479(n607 ,n606);
    nor g2480(n606 ,n481 ,n605);
    xnor g2481(n2490 ,n543 ,n510);
    nor g2482(n605 ,n510 ,n543);
    nor g2483(n2489 ,n510 ,n509);
    xnor g2484(n604 ,n2607 ,n11[39]);
    xnor g2485(n603 ,n2614 ,n11[46]);
    xnor g2486(n602 ,n2575 ,n11[39]);
    xnor g2487(n601 ,n2597 ,n11[45]);
    xnor g2488(n600 ,n2559 ,n11[39]);
    xnor g2489(n599 ,n2574 ,n11[38]);
    xnor g2490(n598 ,n2561 ,n11[41]);
    xnor g2491(n597 ,n2596 ,n11[44]);
    xnor g2492(n596 ,n2573 ,n11[37]);
    xnor g2493(n595 ,n2582 ,n11[46]);
    xnor g2494(n594 ,n2572 ,n11[36]);
    xnor g2495(n593 ,n2615 ,n10[62]);
    xnor g2496(n592 ,n2606 ,n11[38]);
    xnor g2497(n591 ,n2571 ,n11[35]);
    xnor g2498(n590 ,n2612 ,n11[44]);
    xnor g2499(n589 ,n2595 ,n11[43]);
    xnor g2500(n588 ,n2570 ,n11[34]);
    xnor g2501(n587 ,n2611 ,n11[43]);
    xnor g2502(n586 ,n2569 ,n11[33]);
    xnor g2503(n585 ,n2594 ,n11[42]);
    xnor g2504(n584 ,n2565 ,n11[45]);
    xnor g2505(n583 ,n2568 ,n11[32]);
    xnor g2506(n582 ,n2583 ,n11[31]);
    xnor g2507(n581 ,n2567 ,n11[31]);
    xnor g2508(n580 ,n2593 ,n11[41]);
    xnor g2509(n579 ,n2605 ,n11[37]);
    xnor g2510(n578 ,n2566 ,n11[46]);
    xnor g2511(n577 ,n2584 ,n11[32]);
    xnor g2512(n576 ,n2592 ,n11[40]);
    xnor g2513(n575 ,n2608 ,n11[40]);
    xnor g2514(n574 ,n2576 ,n11[40]);
    xnor g2515(n573 ,n2591 ,n11[39]);
    xnor g2516(n572 ,n2563 ,n11[43]);
    xnor g2517(n571 ,n2562 ,n11[42]);
    xnor g2518(n570 ,n2604 ,n11[36]);
    xnor g2519(n569 ,n2610 ,n11[42]);
    xnor g2520(n568 ,n2560 ,n11[40]);
    xnor g2521(n567 ,n2589 ,n11[37]);
    xnor g2522(n566 ,n2558 ,n11[38]);
    xnor g2523(n565 ,n2613 ,n11[45]);
    xnor g2524(n564 ,n2603 ,n11[35]);
    xnor g2525(n563 ,n2588 ,n11[36]);
    xnor g2526(n562 ,n2556 ,n11[36]);
    xnor g2527(n561 ,n2587 ,n11[35]);
    xnor g2528(n560 ,n2555 ,n11[35]);
    xnor g2529(n559 ,n2599 ,n11[31]);
    xnor g2530(n558 ,n2564 ,n11[44]);
    xnor g2531(n557 ,n2586 ,n11[34]);
    xnor g2532(n556 ,n2598 ,n11[46]);
    xnor g2533(n555 ,n2602 ,n11[34]);
    xnor g2534(n554 ,n2609 ,n11[41]);
    xnor g2535(n553 ,n2578 ,n11[42]);
    xnor g2536(n552 ,n2579 ,n11[43]);
    xnor g2537(n551 ,n2601 ,n11[33]);
    xnor g2538(n550 ,n2577 ,n11[41]);
    xnor g2539(n549 ,n2580 ,n11[44]);
    xnor g2540(n548 ,n2581 ,n11[45]);
    xnor g2541(n547 ,n2585 ,n11[33]);
    xnor g2542(n546 ,n2557 ,n11[37]);
    xnor g2543(n545 ,n2590 ,n11[38]);
    xnor g2544(n544 ,n2600 ,n11[32]);
    xnor g2545(n543 ,n2554 ,n11[34]);
    nor g2546(n542 ,n475 ,n439);
    nor g2547(n541 ,n427 ,n406);
    nor g2548(n540 ,n458 ,n447);
    nor g2549(n539 ,n436 ,n406);
    nor g2550(n538 ,n478 ,n447);
    nor g2551(n537 ,n449 ,n406);
    nor g2552(n536 ,n456 ,n447);
    nor g2553(n535 ,n466 ,n405);
    nor g2554(n534 ,n471 ,n443);
    nor g2555(n533 ,n464 ,n404);
    nor g2556(n532 ,n417 ,n400);
    nor g2557(n531 ,n429 ,n441);
    nor g2558(n530 ,n414 ,n439);
    nor g2559(n529 ,n430 ,n440);
    nor g2560(n528 ,n453 ,n442);
    nor g2561(n527 ,n463 ,n441);
    nor g2562(n526 ,n409 ,n468);
    nor g2563(n525 ,n425 ,n446);
    nor g2564(n524 ,n413 ,n446);
    nor g2565(n523 ,n473 ,n401);
    nor g2566(n522 ,n437 ,n403);
    nor g2567(n521 ,n412 ,n402);
    nor g2568(n520 ,n416 ,n445);
    nor g2569(n519 ,n422 ,n440);
    nor g2570(n518 ,n469 ,n405);
    nor g2571(n517 ,n410 ,n404);
    nor g2572(n516 ,n455 ,n403);
    nor g2573(n515 ,n452 ,n404);
    nor g2574(n514 ,n460 ,n443);
    nor g2575(n513 ,n420 ,n439);
    nor g2576(n512 ,n448 ,n400);
    nor g2577(n511 ,n434 ,n439);
    nor g2578(n509 ,n2553 ,n11[33]);
    nor g2579(n508 ,n477 ,n402);
    nor g2580(n507 ,n421 ,n441);
    nor g2581(n506 ,n451 ,n405);
    nor g2582(n505 ,n474 ,n444);
    nor g2583(n504 ,n415 ,n446);
    nor g2584(n503 ,n426 ,n440);
    nor g2585(n502 ,n467 ,n400);
    nor g2586(n501 ,n462 ,n441);
    nor g2587(n500 ,n433 ,n442);
    nor g2588(n499 ,n450 ,n440);
    nor g2589(n498 ,n457 ,n442);
    nor g2590(n497 ,n408 ,n405);
    nor g2591(n496 ,n418 ,n401);
    nor g2592(n495 ,n407 ,n444);
    nor g2593(n494 ,n435 ,n402);
    nor g2594(n493 ,n419 ,n443);
    nor g2595(n492 ,n459 ,n403);
    nor g2596(n491 ,n424 ,n442);
    nor g2597(n490 ,n476 ,n402);
    nor g2598(n489 ,n470 ,n401);
    nor g2599(n488 ,n432 ,n446);
    nor g2600(n487 ,n428 ,n445);
    nor g2601(n486 ,n461 ,n443);
    nor g2602(n485 ,n423 ,n444);
    nor g2603(n484 ,n472 ,n403);
    nor g2604(n483 ,n438 ,n445);
    nor g2605(n482 ,n431 ,n400);
    nor g2606(n481 ,n2554 ,n11[34]);
    nor g2607(n480 ,n454 ,n404);
    nor g2608(n479 ,n465 ,n444);
    nor g2609(n510 ,n411 ,n445);
    not g2610(n478 ,n2584);
    not g2611(n477 ,n2562);
    not g2612(n476 ,n2610);
    not g2613(n475 ,n2595);
    not g2614(n474 ,n2560);
    not g2615(n473 ,n2570);
    not g2616(n472 ,n2614);
    not g2617(n471 ,n2596);
    not g2618(n470 ,n2602);
    not g2619(n469 ,n2593);
    not g2620(n468 ,n10[62]);
    not g2621(n467 ,n2559);
    not g2622(n466 ,n2577);
    not g2623(n465 ,n2592);
    not g2624(n464 ,n2597);
    not g2625(n463 ,n2606);
    not g2626(n462 ,n2558);
    not g2627(n461 ,n2580);
    not g2628(n460 ,n2564);
    not g2629(n459 ,n2598);
    not g2630(n458 ,n2568);
    not g2631(n457 ,n2556);
    not g2632(n456 ,n2600);
    not g2633(n455 ,n2566);
    not g2634(n454 ,n2581);
    not g2635(n453 ,n2572);
    not g2636(n452 ,n2565);
    not g2637(n451 ,n2561);
    not g2638(n450 ,n2557);
    not g2639(n449 ,n2583);
    not g2640(n448 ,n2591);
    not g2641(n447 ,n11[32]);
    not g2642(n446 ,n11[35]);
    not g2643(n445 ,n11[33]);
    not g2644(n444 ,n11[40]);
    not g2645(n443 ,n11[44]);
    not g2646(n442 ,n11[36]);
    not g2647(n441 ,n11[38]);
    not g2648(n440 ,n11[37]);
    not g2649(n439 ,n11[43]);
    not g2650(n438 ,n2601);
    not g2651(n437 ,n2582);
    not g2652(n436 ,n2567);
    not g2653(n435 ,n2578);
    not g2654(n434 ,n2563);
    not g2655(n433 ,n2588);
    not g2656(n432 ,n2587);
    not g2657(n431 ,n2607);
    not g2658(n430 ,n2573);
    not g2659(n429 ,n2574);
    not g2660(n428 ,n2585);
    not g2661(n427 ,n2599);
    not g2662(n426 ,n2589);
    not g2663(n425 ,n2571);
    not g2664(n424 ,n2604);
    not g2665(n423 ,n2608);
    not g2666(n422 ,n2605);
    not g2667(n421 ,n2590);
    not g2668(n420 ,n2579);
    not g2669(n419 ,n2612);
    not g2670(n418 ,n2586);
    not g2671(n417 ,n2575);
    not g2672(n416 ,n2569);
    not g2673(n415 ,n2603);
    not g2674(n414 ,n2611);
    not g2675(n413 ,n2555);
    not g2676(n412 ,n2594);
    not g2677(n411 ,n2553);
    not g2678(n410 ,n2613);
    not g2679(n409 ,n2615);
    not g2680(n408 ,n2609);
    not g2681(n407 ,n2576);
    not g2682(n406 ,n11[31]);
    not g2683(n405 ,n11[41]);
    not g2684(n404 ,n11[45]);
    not g2685(n403 ,n11[46]);
    not g2686(n402 ,n11[42]);
    not g2687(n401 ,n11[34]);
    not g2688(n400 ,n11[39]);
    xnor g2689(n2934 ,n798 ,n986);
    nor g2690(n986 ,n771 ,n985);
    xnor g2691(n2932 ,n814 ,n984);
    nor g2692(n985 ,n814 ,n984);
    nor g2693(n984 ,n760 ,n983);
    xnor g2694(n2930 ,n835 ,n982);
    nor g2695(n983 ,n835 ,n982);
    nor g2696(n982 ,n789 ,n981);
    xnor g2697(n2928 ,n817 ,n980);
    nor g2698(n981 ,n817 ,n980);
    nor g2699(n980 ,n763 ,n979);
    xnor g2700(n2926 ,n822 ,n978);
    nor g2701(n979 ,n822 ,n978);
    nor g2702(n978 ,n775 ,n977);
    xnor g2703(n2924 ,n844 ,n976);
    nor g2704(n977 ,n844 ,n976);
    nor g2705(n976 ,n756 ,n975);
    xnor g2706(n2922 ,n827 ,n974);
    nor g2707(n975 ,n827 ,n974);
    nor g2708(n974 ,n790 ,n973);
    xnor g2709(n2920 ,n816 ,n972);
    nor g2710(n973 ,n816 ,n972);
    nor g2711(n972 ,n736 ,n971);
    xnor g2712(n2918 ,n855 ,n970);
    nor g2713(n971 ,n855 ,n970);
    nor g2714(n970 ,n755 ,n969);
    xnor g2715(n2916 ,n809 ,n968);
    nor g2716(n969 ,n809 ,n968);
    nor g2717(n968 ,n782 ,n967);
    xnor g2718(n2914 ,n850 ,n966);
    nor g2719(n967 ,n850 ,n966);
    nor g2720(n966 ,n767 ,n965);
    xnor g2721(n2912 ,n845 ,n964);
    nor g2722(n965 ,n845 ,n964);
    nor g2723(n964 ,n759 ,n963);
    xnor g2724(n2910 ,n839 ,n962);
    nor g2725(n963 ,n839 ,n962);
    nor g2726(n962 ,n751 ,n961);
    xnor g2727(n2908 ,n831 ,n960);
    nor g2728(n961 ,n831 ,n960);
    nor g2729(n960 ,n747 ,n959);
    xnor g2730(n2906 ,n820 ,n958);
    nor g2731(n959 ,n820 ,n958);
    nor g2732(n958 ,n741 ,n957);
    xnor g2733(n2904 ,n829 ,n956);
    nor g2734(n957 ,n829 ,n956);
    nor g2735(n956 ,n734 ,n955);
    xnor g2736(n2902 ,n805 ,n954);
    nor g2737(n955 ,n805 ,n954);
    nor g2738(n954 ,n777 ,n953);
    xnor g2739(n2900 ,n800 ,n952);
    nor g2740(n953 ,n800 ,n952);
    nor g2741(n952 ,n795 ,n951);
    xnor g2742(n2898 ,n802 ,n950);
    nor g2743(n951 ,n802 ,n950);
    nor g2744(n950 ,n776 ,n949);
    xnor g2745(n2896 ,n808 ,n948);
    nor g2746(n949 ,n808 ,n948);
    nor g2747(n948 ,n783 ,n947);
    xnor g2748(n2894 ,n857 ,n946);
    nor g2749(n947 ,n857 ,n946);
    nor g2750(n946 ,n750 ,n945);
    xnor g2751(n2892 ,n853 ,n944);
    nor g2752(n945 ,n853 ,n944);
    nor g2753(n944 ,n769 ,n943);
    xnor g2754(n2890 ,n848 ,n942);
    nor g2755(n943 ,n848 ,n942);
    nor g2756(n942 ,n745 ,n941);
    xnor g2757(n2888 ,n818 ,n940);
    nor g2758(n941 ,n818 ,n940);
    nor g2759(n940 ,n761 ,n939);
    xnor g2760(n2886 ,n842 ,n938);
    nor g2761(n939 ,n842 ,n938);
    nor g2762(n938 ,n786 ,n937);
    xnor g2763(n2884 ,n838 ,n936);
    nor g2764(n937 ,n838 ,n936);
    nor g2765(n936 ,n753 ,n935);
    xnor g2766(n2882 ,n833 ,n934);
    nor g2767(n935 ,n833 ,n934);
    nor g2768(n934 ,n758 ,n933);
    xnor g2769(n2880 ,n830 ,n932);
    nor g2770(n933 ,n830 ,n932);
    nor g2771(n932 ,n773 ,n931);
    xnor g2772(n2878 ,n828 ,n930);
    nor g2773(n931 ,n828 ,n930);
    nor g2774(n930 ,n737 ,n929);
    xnor g2775(n2876 ,n824 ,n928);
    nor g2776(n929 ,n824 ,n928);
    nor g2777(n928 ,n743 ,n927);
    xnor g2778(n2874 ,n819 ,n926);
    nor g2779(n927 ,n819 ,n926);
    nor g2780(n926 ,n766 ,n925);
    xnor g2781(n2872 ,n812 ,n924);
    nor g2782(n925 ,n812 ,n924);
    nor g2783(n924 ,n792 ,n923);
    xnor g2784(n2870 ,n807 ,n922);
    nor g2785(n923 ,n807 ,n922);
    nor g2786(n922 ,n793 ,n921);
    xnor g2787(n2868 ,n804 ,n920);
    nor g2788(n921 ,n804 ,n920);
    nor g2789(n920 ,n735 ,n919);
    xnor g2790(n2866 ,n799 ,n918);
    nor g2791(n919 ,n799 ,n918);
    nor g2792(n918 ,n772 ,n917);
    xnor g2793(n2864 ,n801 ,n916);
    nor g2794(n917 ,n801 ,n916);
    nor g2795(n916 ,n787 ,n915);
    xnor g2796(n2862 ,n803 ,n914);
    nor g2797(n915 ,n803 ,n914);
    nor g2798(n914 ,n784 ,n913);
    xnor g2799(n2860 ,n806 ,n912);
    nor g2800(n913 ,n806 ,n912);
    nor g2801(n912 ,n764 ,n911);
    xnor g2802(n2858 ,n811 ,n910);
    nor g2803(n911 ,n811 ,n910);
    nor g2804(n910 ,n762 ,n909);
    xnor g2805(n2856 ,n810 ,n908);
    nor g2806(n909 ,n810 ,n908);
    nor g2807(n908 ,n738 ,n907);
    xnor g2808(n2854 ,n859 ,n906);
    nor g2809(n907 ,n859 ,n906);
    nor g2810(n906 ,n781 ,n905);
    xnor g2811(n2852 ,n856 ,n904);
    nor g2812(n905 ,n856 ,n904);
    nor g2813(n904 ,n778 ,n903);
    xnor g2814(n2850 ,n854 ,n902);
    nor g2815(n903 ,n854 ,n902);
    nor g2816(n902 ,n774 ,n901);
    xnor g2817(n2848 ,n852 ,n900);
    nor g2818(n901 ,n852 ,n900);
    nor g2819(n900 ,n770 ,n899);
    xnor g2820(n2846 ,n851 ,n898);
    nor g2821(n899 ,n851 ,n898);
    nor g2822(n898 ,n768 ,n897);
    xnor g2823(n2844 ,n849 ,n896);
    nor g2824(n897 ,n849 ,n896);
    nor g2825(n896 ,n749 ,n895);
    xnor g2826(n2842 ,n846 ,n894);
    nor g2827(n895 ,n846 ,n894);
    nor g2828(n894 ,n740 ,n893);
    xnor g2829(n2840 ,n825 ,n892);
    nor g2830(n893 ,n825 ,n892);
    nor g2831(n892 ,n742 ,n891);
    xnor g2832(n2838 ,n843 ,n890);
    nor g2833(n891 ,n843 ,n890);
    nor g2834(n890 ,n785 ,n889);
    xnor g2835(n2836 ,n841 ,n888);
    nor g2836(n889 ,n841 ,n888);
    nor g2837(n888 ,n757 ,n887);
    xnor g2838(n2834 ,n840 ,n886);
    nor g2839(n887 ,n840 ,n886);
    nor g2840(n886 ,n754 ,n885);
    xnor g2841(n2832 ,n837 ,n884);
    nor g2842(n885 ,n837 ,n884);
    nor g2843(n884 ,n788 ,n883);
    xnor g2844(n2830 ,n836 ,n882);
    nor g2845(n883 ,n836 ,n882);
    nor g2846(n882 ,n752 ,n881);
    xnor g2847(n2828 ,n834 ,n880);
    nor g2848(n881 ,n834 ,n880);
    nor g2849(n880 ,n765 ,n879);
    xnor g2850(n2826 ,n832 ,n878);
    nor g2851(n879 ,n832 ,n878);
    nor g2852(n878 ,n748 ,n877);
    xnor g2853(n2824 ,n847 ,n876);
    nor g2854(n877 ,n847 ,n876);
    nor g2855(n876 ,n779 ,n875);
    xnor g2856(n2822 ,n813 ,n874);
    nor g2857(n875 ,n813 ,n874);
    nor g2858(n874 ,n746 ,n873);
    xnor g2859(n2820 ,n858 ,n872);
    nor g2860(n873 ,n858 ,n872);
    nor g2861(n872 ,n744 ,n871);
    xnor g2862(n2818 ,n826 ,n870);
    nor g2863(n871 ,n826 ,n870);
    nor g2864(n870 ,n794 ,n869);
    xnor g2865(n2816 ,n823 ,n868);
    nor g2866(n869 ,n823 ,n868);
    nor g2867(n868 ,n791 ,n867);
    xor g2868(n2814 ,n821 ,n865);
    nor g2869(n867 ,n821 ,n866);
    not g2870(n866 ,n865);
    nor g2871(n865 ,n780 ,n864);
    xnor g2872(n2812 ,n860 ,n862);
    nor g2873(n864 ,n860 ,n863);
    not g2874(n863 ,n862);
    nor g2875(n862 ,n739 ,n861);
    xnor g2876(n2810 ,n815 ,n797);
    nor g2877(n861 ,n797 ,n815);
    nor g2878(n2745 ,n797 ,n796);
    xnor g2879(n860 ,n2[2] ,n2[66]);
    xnor g2880(n859 ,n2[23] ,n2[87]);
    xnor g2881(n858 ,n2[6] ,n2[70]);
    xnor g2882(n857 ,n2[43] ,n2[107]);
    xnor g2883(n856 ,n2[22] ,n2[86]);
    xnor g2884(n855 ,n2[55] ,n2[119]);
    xnor g2885(n854 ,n2[21] ,n2[85]);
    xnor g2886(n853 ,n2[42] ,n2[106]);
    xnor g2887(n852 ,n2[20] ,n2[84]);
    xnor g2888(n851 ,n2[19] ,n2[83]);
    xnor g2889(n850 ,n2[53] ,n2[117]);
    xnor g2890(n849 ,n2[18] ,n2[82]);
    xnor g2891(n848 ,n2[41] ,n2[105]);
    xnor g2892(n847 ,n2[8] ,n2[72]);
    xnor g2893(n846 ,n2[17] ,n2[81]);
    xnor g2894(n845 ,n2[52] ,n2[116]);
    xnor g2895(n844 ,n2[58] ,n2[122]);
    xnor g2896(n843 ,n2[15] ,n2[79]);
    xnor g2897(n842 ,n2[39] ,n2[103]);
    xnor g2898(n841 ,n2[14] ,n2[78]);
    xnor g2899(n840 ,n2[13] ,n2[77]);
    xnor g2900(n839 ,n2[51] ,n2[115]);
    xnor g2901(n838 ,n2[38] ,n2[102]);
    xnor g2902(n837 ,n2[12] ,n2[76]);
    xnor g2903(n836 ,n2[11] ,n2[75]);
    xnor g2904(n835 ,n2[61] ,n2[125]);
    xnor g2905(n834 ,n2[10] ,n2[74]);
    xnor g2906(n833 ,n2[37] ,n2[101]);
    xnor g2907(n832 ,n2[9] ,n2[73]);
    xnor g2908(n831 ,n2[50] ,n2[114]);
    xnor g2909(n830 ,n2[36] ,n2[100]);
    xnor g2910(n829 ,n2[48] ,n2[112]);
    xnor g2911(n828 ,n2[35] ,n2[99]);
    xnor g2912(n827 ,n2[57] ,n2[121]);
    xnor g2913(n826 ,n2[5] ,n2[69]);
    xnor g2914(n825 ,n2[16] ,n2[80]);
    xnor g2915(n824 ,n2[34] ,n2[98]);
    xnor g2916(n823 ,n2[4] ,n2[68]);
    xnor g2917(n822 ,n2[59] ,n2[123]);
    xnor g2918(n821 ,n2[3] ,n2[67]);
    xnor g2919(n820 ,n2[49] ,n2[113]);
    xnor g2920(n819 ,n2[33] ,n2[97]);
    xnor g2921(n818 ,n2[40] ,n2[104]);
    xnor g2922(n817 ,n2[60] ,n2[124]);
    xnor g2923(n816 ,n2[56] ,n2[120]);
    xnor g2924(n815 ,n2[1] ,n2[65]);
    xnor g2925(n814 ,n2[62] ,n2[126]);
    xnor g2926(n813 ,n2[7] ,n2[71]);
    xnor g2927(n812 ,n2[32] ,n2[96]);
    xnor g2928(n811 ,n2[25] ,n2[89]);
    xnor g2929(n810 ,n2[24] ,n2[88]);
    xnor g2930(n809 ,n2[54] ,n2[118]);
    xnor g2931(n808 ,n2[44] ,n2[108]);
    xnor g2932(n807 ,n2[31] ,n2[95]);
    xnor g2933(n806 ,n2[26] ,n2[90]);
    xnor g2934(n805 ,n2[47] ,n2[111]);
    xnor g2935(n804 ,n2[30] ,n2[94]);
    xnor g2936(n803 ,n2[27] ,n2[91]);
    xnor g2937(n802 ,n2[45] ,n2[109]);
    xnor g2938(n801 ,n2[28] ,n2[92]);
    xnor g2939(n800 ,n2[46] ,n2[110]);
    xnor g2940(n799 ,n2[29] ,n2[93]);
    xnor g2941(n798 ,n2[63] ,n2[127]);
    nor g2942(n796 ,n2[0] ,n2[64]);
    nor g2943(n795 ,n2[45] ,n2[109]);
    nor g2944(n794 ,n2[4] ,n2[68]);
    nor g2945(n793 ,n2[30] ,n2[94]);
    nor g2946(n792 ,n2[31] ,n2[95]);
    nor g2947(n791 ,n2[3] ,n2[67]);
    nor g2948(n790 ,n2[56] ,n2[120]);
    nor g2949(n789 ,n2[60] ,n2[124]);
    nor g2950(n788 ,n2[11] ,n2[75]);
    nor g2951(n787 ,n2[27] ,n2[91]);
    nor g2952(n786 ,n2[38] ,n2[102]);
    nor g2953(n785 ,n2[14] ,n2[78]);
    nor g2954(n784 ,n2[26] ,n2[90]);
    nor g2955(n783 ,n2[43] ,n2[107]);
    nor g2956(n782 ,n2[53] ,n2[117]);
    nor g2957(n781 ,n2[22] ,n2[86]);
    nor g2958(n780 ,n732 ,n731);
    nor g2959(n779 ,n2[7] ,n2[71]);
    nor g2960(n778 ,n2[21] ,n2[85]);
    nor g2961(n777 ,n2[46] ,n2[110]);
    nor g2962(n776 ,n2[44] ,n2[108]);
    nor g2963(n775 ,n2[58] ,n2[122]);
    nor g2964(n774 ,n2[20] ,n2[84]);
    nor g2965(n773 ,n2[35] ,n2[99]);
    nor g2966(n772 ,n2[28] ,n2[92]);
    nor g2967(n771 ,n2[62] ,n2[126]);
    nor g2968(n770 ,n2[19] ,n2[83]);
    nor g2969(n769 ,n2[41] ,n2[105]);
    nor g2970(n768 ,n2[18] ,n2[82]);
    nor g2971(n767 ,n2[52] ,n2[116]);
    nor g2972(n766 ,n2[32] ,n2[96]);
    nor g2973(n797 ,n733 ,n730);
    nor g2974(n765 ,n2[9] ,n2[73]);
    nor g2975(n764 ,n2[25] ,n2[89]);
    nor g2976(n763 ,n2[59] ,n2[123]);
    nor g2977(n762 ,n2[24] ,n2[88]);
    nor g2978(n761 ,n2[39] ,n2[103]);
    nor g2979(n760 ,n2[61] ,n2[125]);
    nor g2980(n759 ,n2[51] ,n2[115]);
    nor g2981(n758 ,n2[36] ,n2[100]);
    nor g2982(n757 ,n2[13] ,n2[77]);
    nor g2983(n756 ,n2[57] ,n2[121]);
    nor g2984(n755 ,n2[54] ,n2[118]);
    nor g2985(n754 ,n2[12] ,n2[76]);
    nor g2986(n753 ,n2[37] ,n2[101]);
    nor g2987(n752 ,n2[10] ,n2[74]);
    nor g2988(n751 ,n2[50] ,n2[114]);
    nor g2989(n750 ,n2[42] ,n2[106]);
    nor g2990(n749 ,n2[17] ,n2[81]);
    nor g2991(n748 ,n2[8] ,n2[72]);
    nor g2992(n747 ,n2[49] ,n2[113]);
    nor g2993(n746 ,n2[6] ,n2[70]);
    nor g2994(n745 ,n2[40] ,n2[104]);
    nor g2995(n744 ,n2[5] ,n2[69]);
    nor g2996(n743 ,n2[33] ,n2[97]);
    nor g2997(n742 ,n2[15] ,n2[79]);
    nor g2998(n741 ,n2[48] ,n2[112]);
    nor g2999(n740 ,n2[16] ,n2[80]);
    nor g3000(n739 ,n2[1] ,n2[65]);
    nor g3001(n738 ,n2[23] ,n2[87]);
    nor g3002(n737 ,n2[34] ,n2[98]);
    nor g3003(n736 ,n2[55] ,n2[119]);
    nor g3004(n735 ,n2[29] ,n2[93]);
    nor g3005(n734 ,n2[47] ,n2[111]);
    not g3006(n733 ,n2[0]);
    not g3007(n732 ,n2[2]);
    not g3008(n731 ,n2[66]);
    not g3009(n730 ,n2[64]);
    xnor g3010(n2808 ,n1062 ,n1251);
    nor g3011(n1251 ,n1000 ,n1250);
    xnor g3012(n2807 ,n1072 ,n1249);
    nor g3013(n1250 ,n1072 ,n1249);
    nor g3014(n1249 ,n1048 ,n1248);
    xnor g3015(n2806 ,n1088 ,n1247);
    nor g3016(n1248 ,n1088 ,n1247);
    nor g3017(n1247 ,n1021 ,n1246);
    xnor g3018(n2805 ,n1070 ,n1245);
    nor g3019(n1246 ,n1070 ,n1245);
    nor g3020(n1245 ,n1004 ,n1244);
    xnor g3021(n2804 ,n1116 ,n1243);
    nor g3022(n1244 ,n1116 ,n1243);
    nor g3023(n1243 ,n1027 ,n1242);
    xnor g3024(n2803 ,n1099 ,n1241);
    nor g3025(n1242 ,n1099 ,n1241);
    nor g3026(n1241 ,n1025 ,n1240);
    xnor g3027(n2802 ,n1093 ,n1239);
    nor g3028(n1240 ,n1093 ,n1239);
    nor g3029(n1239 ,n1008 ,n1238);
    xnor g3030(n2801 ,n1107 ,n1237);
    nor g3031(n1238 ,n1107 ,n1237);
    nor g3032(n1237 ,n1046 ,n1236);
    xnor g3033(n2800 ,n1082 ,n1235);
    nor g3034(n1236 ,n1082 ,n1235);
    nor g3035(n1235 ,n1051 ,n1234);
    xnor g3036(n2799 ,n1114 ,n1233);
    nor g3037(n1234 ,n1114 ,n1233);
    nor g3038(n1233 ,n1011 ,n1232);
    xnor g3039(n2798 ,n1103 ,n1231);
    nor g3040(n1232 ,n1103 ,n1231);
    nor g3041(n1231 ,n1034 ,n1230);
    xnor g3042(n2797 ,n1108 ,n1229);
    nor g3043(n1230 ,n1108 ,n1229);
    nor g3044(n1229 ,n1043 ,n1228);
    xnor g3045(n2796 ,n1090 ,n1227);
    nor g3046(n1228 ,n1090 ,n1227);
    nor g3047(n1227 ,n1022 ,n1226);
    xnor g3048(n2795 ,n1084 ,n1225);
    nor g3049(n1226 ,n1084 ,n1225);
    nor g3050(n1225 ,n1009 ,n1224);
    xnor g3051(n2794 ,n1064 ,n1223);
    nor g3052(n1224 ,n1064 ,n1223);
    nor g3053(n1223 ,n1042 ,n1222);
    xnor g3054(n2793 ,n1063 ,n1221);
    nor g3055(n1222 ,n1063 ,n1221);
    nor g3056(n1221 ,n1012 ,n1220);
    xnor g3057(n2792 ,n1078 ,n1219);
    nor g3058(n1220 ,n1078 ,n1219);
    nor g3059(n1219 ,n1015 ,n1218);
    xnor g3060(n2791 ,n1087 ,n1217);
    nor g3061(n1218 ,n1087 ,n1217);
    nor g3062(n1217 ,n1054 ,n1216);
    xnor g3063(n2790 ,n1079 ,n1215);
    nor g3064(n1216 ,n1079 ,n1215);
    nor g3065(n1215 ,n1049 ,n1214);
    xnor g3066(n2789 ,n1117 ,n1213);
    nor g3067(n1214 ,n1117 ,n1213);
    nor g3068(n1213 ,n1047 ,n1212);
    xnor g3069(n2788 ,n1112 ,n1211);
    nor g3070(n1212 ,n1112 ,n1211);
    nor g3071(n1211 ,n1045 ,n1210);
    xnor g3072(n2787 ,n1109 ,n1209);
    nor g3073(n1210 ,n1109 ,n1209);
    nor g3074(n1209 ,n1040 ,n1208);
    xnor g3075(n2786 ,n1106 ,n1207);
    nor g3076(n1208 ,n1106 ,n1207);
    nor g3077(n1207 ,n1016 ,n1206);
    xnor g3078(n2785 ,n1102 ,n1205);
    nor g3079(n1206 ,n1102 ,n1205);
    nor g3080(n1205 ,n1037 ,n1204);
    xnor g3081(n2784 ,n1098 ,n1203);
    nor g3082(n1204 ,n1098 ,n1203);
    nor g3083(n1203 ,n1001 ,n1202);
    xnor g3084(n2783 ,n1096 ,n1201);
    nor g3085(n1202 ,n1096 ,n1201);
    nor g3086(n1201 ,n1018 ,n1200);
    xnor g3087(n2782 ,n1077 ,n1199);
    nor g3088(n1200 ,n1077 ,n1199);
    nor g3089(n1199 ,n1024 ,n1198);
    xnor g3090(n2781 ,n1089 ,n1197);
    nor g3091(n1198 ,n1089 ,n1197);
    nor g3092(n1197 ,n1029 ,n1196);
    xnor g3093(n2780 ,n1086 ,n1195);
    nor g3094(n1196 ,n1086 ,n1195);
    nor g3095(n1195 ,n1030 ,n1194);
    xnor g3096(n2779 ,n1083 ,n1193);
    nor g3097(n1194 ,n1083 ,n1193);
    nor g3098(n1193 ,n1017 ,n1192);
    xnor g3099(n2778 ,n1066 ,n1191);
    nor g3100(n1192 ,n1066 ,n1191);
    nor g3101(n1191 ,n1052 ,n1190);
    xnor g3102(n2777 ,n1065 ,n1189);
    nor g3103(n1190 ,n1065 ,n1189);
    nor g3104(n1189 ,n1041 ,n1188);
    xnor g3105(n2776 ,n1074 ,n1187);
    nor g3106(n1188 ,n1074 ,n1187);
    nor g3107(n1187 ,n1013 ,n1186);
    xnor g3108(n2775 ,n1071 ,n1185);
    nor g3109(n1186 ,n1071 ,n1185);
    nor g3110(n1185 ,n1005 ,n1184);
    xnor g3111(n2774 ,n1073 ,n1183);
    nor g3112(n1184 ,n1073 ,n1183);
    nor g3113(n1183 ,n1006 ,n1182);
    xnor g3114(n2773 ,n1075 ,n1181);
    nor g3115(n1182 ,n1075 ,n1181);
    nor g3116(n1181 ,n1002 ,n1180);
    xnor g3117(n2772 ,n1081 ,n1179);
    nor g3118(n1180 ,n1081 ,n1179);
    nor g3119(n1179 ,n1055 ,n1178);
    xnor g3120(n2771 ,n1076 ,n1177);
    nor g3121(n1178 ,n1076 ,n1177);
    nor g3122(n1177 ,n1023 ,n1176);
    xnor g3123(n2770 ,n1091 ,n1175);
    nor g3124(n1176 ,n1091 ,n1175);
    nor g3125(n1175 ,n1033 ,n1174);
    xnor g3126(n2769 ,n1080 ,n1173);
    nor g3127(n1174 ,n1080 ,n1173);
    nor g3128(n1173 ,n1053 ,n1172);
    xnor g3129(n2768 ,n1119 ,n1171);
    nor g3130(n1172 ,n1119 ,n1171);
    nor g3131(n1171 ,n1050 ,n1170);
    xnor g3132(n2767 ,n1118 ,n1169);
    nor g3133(n1170 ,n1118 ,n1169);
    nor g3134(n1169 ,n1039 ,n1168);
    xnor g3135(n2766 ,n1115 ,n1167);
    nor g3136(n1168 ,n1115 ,n1167);
    nor g3137(n1167 ,n1014 ,n1166);
    xnor g3138(n2765 ,n1113 ,n1165);
    nor g3139(n1166 ,n1113 ,n1165);
    nor g3140(n1165 ,n1010 ,n1164);
    xnor g3141(n2764 ,n1111 ,n1163);
    nor g3142(n1164 ,n1111 ,n1163);
    nor g3143(n1163 ,n1044 ,n1162);
    xnor g3144(n2763 ,n1110 ,n1161);
    nor g3145(n1162 ,n1110 ,n1161);
    nor g3146(n1161 ,n1038 ,n1160);
    xnor g3147(n2762 ,n1068 ,n1159);
    nor g3148(n1160 ,n1068 ,n1159);
    nor g3149(n1159 ,n1019 ,n1158);
    xnor g3150(n2761 ,n1067 ,n1157);
    nor g3151(n1158 ,n1067 ,n1157);
    nor g3152(n1157 ,n999 ,n1156);
    xnor g3153(n2760 ,n1105 ,n1155);
    nor g3154(n1156 ,n1105 ,n1155);
    nor g3155(n1155 ,n1036 ,n1154);
    xnor g3156(n2759 ,n1104 ,n1153);
    nor g3157(n1154 ,n1104 ,n1153);
    nor g3158(n1153 ,n1003 ,n1152);
    xnor g3159(n2758 ,n1101 ,n1151);
    nor g3160(n1152 ,n1101 ,n1151);
    nor g3161(n1151 ,n1035 ,n1150);
    xor g3162(n2757 ,n1100 ,n1148);
    nor g3163(n1150 ,n1100 ,n1149);
    not g3164(n1149 ,n1148);
    nor g3165(n1148 ,n1056 ,n1147);
    xnor g3166(n2756 ,n1123 ,n1145);
    nor g3167(n1147 ,n1123 ,n1146);
    not g3168(n1146 ,n1145);
    nor g3169(n1145 ,n1032 ,n1144);
    xor g3170(n2755 ,n1097 ,n1142);
    nor g3171(n1144 ,n1097 ,n1143);
    not g3172(n1143 ,n1142);
    nor g3173(n1142 ,n1031 ,n1141);
    xnor g3174(n2754 ,n1094 ,n1139);
    nor g3175(n1141 ,n1094 ,n1140);
    not g3176(n1140 ,n1139);
    nor g3177(n1139 ,n1026 ,n1138);
    xnor g3178(n2753 ,n1095 ,n1137);
    nor g3179(n1138 ,n1095 ,n1137);
    nor g3180(n1137 ,n1007 ,n1136);
    xor g3181(n2752 ,n1092 ,n1134);
    nor g3182(n1136 ,n1092 ,n1135);
    not g3183(n1135 ,n1134);
    nor g3184(n1134 ,n1058 ,n1133);
    xor g3185(n2751 ,n1122 ,n1132);
    nor g3186(n1133 ,n1122 ,n1132);
    nor g3187(n1132 ,n1059 ,n1131);
    xor g3188(n2750 ,n1121 ,n1130);
    nor g3189(n1131 ,n1121 ,n1130);
    nor g3190(n1130 ,n1057 ,n1129);
    xnor g3191(n2749 ,n1120 ,n1127);
    nor g3192(n1129 ,n1120 ,n1128);
    not g3193(n1128 ,n1127);
    nor g3194(n1127 ,n1028 ,n1126);
    xnor g3195(n2748 ,n1085 ,n1125);
    nor g3196(n1126 ,n1085 ,n1125);
    nor g3197(n1125 ,n1020 ,n1124);
    xnor g3198(n2747 ,n1069 ,n1061);
    nor g3199(n1124 ,n1061 ,n1069);
    nor g3200(n2746 ,n1061 ,n1060);
    xnor g3201(n1123 ,n2829 ,n11[42]);
    xnor g3202(n1122 ,n2819 ,n11[37]);
    xnor g3203(n1121 ,n2817 ,n11[36]);
    xnor g3204(n1120 ,n2815 ,n11[35]);
    xnor g3205(n1119 ,n2853 ,n11[38]);
    xnor g3206(n1118 ,n2851 ,n11[37]);
    xnor g3207(n1117 ,n2895 ,n11[43]);
    xnor g3208(n1116 ,n2925 ,n11[42]);
    xnor g3209(n1115 ,n2849 ,n11[36]);
    xnor g3210(n1114 ,n2915 ,n11[37]);
    xnor g3211(n1113 ,n2847 ,n11[35]);
    xnor g3212(n1112 ,n2893 ,n11[42]);
    xnor g3213(n1111 ,n2845 ,n11[34]);
    xnor g3214(n1110 ,n2843 ,n11[33]);
    xnor g3215(n1109 ,n2891 ,n11[41]);
    xnor g3216(n1108 ,n2911 ,n11[35]);
    xnor g3217(n1107 ,n2919 ,n11[39]);
    xnor g3218(n1106 ,n2889 ,n11[40]);
    xnor g3219(n1105 ,n2837 ,n11[46]);
    xnor g3220(n1104 ,n2835 ,n11[45]);
    xnor g3221(n1103 ,n2913 ,n11[36]);
    xnor g3222(n1102 ,n2887 ,n11[39]);
    xnor g3223(n1101 ,n2833 ,n11[44]);
    xnor g3224(n1100 ,n2831 ,n11[43]);
    xnor g3225(n1099 ,n2923 ,n11[41]);
    xnor g3226(n1098 ,n2885 ,n11[38]);
    xnor g3227(n1097 ,n2827 ,n11[41]);
    xnor g3228(n1096 ,n2883 ,n11[37]);
    xnor g3229(n1095 ,n2823 ,n11[39]);
    xnor g3230(n1094 ,n2825 ,n11[40]);
    xnor g3231(n1093 ,n2921 ,n11[40]);
    xnor g3232(n1092 ,n2821 ,n11[38]);
    xnor g3233(n1091 ,n2857 ,n11[40]);
    xnor g3234(n1090 ,n2909 ,n11[34]);
    xnor g3235(n1089 ,n2879 ,n11[35]);
    xnor g3236(n1088 ,n2929 ,n11[44]);
    xnor g3237(n1087 ,n2899 ,n11[45]);
    xnor g3238(n1086 ,n2877 ,n11[34]);
    xnor g3239(n1085 ,n2813 ,n11[34]);
    xnor g3240(n1084 ,n2907 ,n11[33]);
    xnor g3241(n1083 ,n2875 ,n11[33]);
    xnor g3242(n1082 ,n2917 ,n11[38]);
    xnor g3243(n1081 ,n2861 ,n11[42]);
    xnor g3244(n1080 ,n2855 ,n11[39]);
    xnor g3245(n1079 ,n2897 ,n11[44]);
    xnor g3246(n1078 ,n2901 ,n11[46]);
    xnor g3247(n1077 ,n2881 ,n11[36]);
    xnor g3248(n1076 ,n2859 ,n11[41]);
    xnor g3249(n1075 ,n2863 ,n11[43]);
    xnor g3250(n1074 ,n2869 ,n11[46]);
    xnor g3251(n1073 ,n2865 ,n11[44]);
    xnor g3252(n1072 ,n2931 ,n11[45]);
    xnor g3253(n1071 ,n2867 ,n11[45]);
    xnor g3254(n1070 ,n2927 ,n11[43]);
    xnor g3255(n1069 ,n2811 ,n11[33]);
    xnor g3256(n1068 ,n2841 ,n11[32]);
    xnor g3257(n1067 ,n2839 ,n11[31]);
    xnor g3258(n1066 ,n2873 ,n11[32]);
    xnor g3259(n1065 ,n2871 ,n11[31]);
    xnor g3260(n1064 ,n2905 ,n11[32]);
    xnor g3261(n1063 ,n2903 ,n11[31]);
    xnor g3262(n1062 ,n11[46] ,n2933);
    nor g3263(n1060 ,n2809 ,n10[49]);
    nor g3264(n1059 ,n998 ,n989);
    nor g3265(n1058 ,n993 ,n987);
    nor g3266(n1057 ,n996 ,n988);
    nor g3267(n1056 ,n992 ,n995);
    nor g3268(n1055 ,n2859 ,n11[41]);
    nor g3269(n1054 ,n2897 ,n11[44]);
    nor g3270(n1053 ,n2853 ,n11[38]);
    nor g3271(n1052 ,n2871 ,n11[31]);
    nor g3272(n1051 ,n2915 ,n11[37]);
    nor g3273(n1050 ,n2851 ,n11[37]);
    nor g3274(n1049 ,n2895 ,n11[43]);
    nor g3275(n1048 ,n2929 ,n11[44]);
    nor g3276(n1047 ,n2893 ,n11[42]);
    nor g3277(n1046 ,n2917 ,n11[38]);
    nor g3278(n1045 ,n2891 ,n11[41]);
    nor g3279(n1044 ,n2843 ,n11[33]);
    nor g3280(n1043 ,n2909 ,n11[34]);
    nor g3281(n1042 ,n2903 ,n11[31]);
    nor g3282(n1041 ,n2869 ,n11[46]);
    nor g3283(n1040 ,n2889 ,n11[40]);
    nor g3284(n1039 ,n2849 ,n11[36]);
    nor g3285(n1038 ,n2841 ,n11[32]);
    nor g3286(n1037 ,n2885 ,n11[38]);
    nor g3287(n1036 ,n2835 ,n11[45]);
    nor g3288(n1035 ,n2831 ,n11[43]);
    nor g3289(n1034 ,n2911 ,n11[35]);
    nor g3290(n1033 ,n2855 ,n11[39]);
    nor g3291(n1032 ,n2827 ,n11[41]);
    nor g3292(n1031 ,n991 ,n994);
    nor g3293(n1061 ,n997 ,n990);
    nor g3294(n1030 ,n2875 ,n11[33]);
    nor g3295(n1029 ,n2877 ,n11[34]);
    nor g3296(n1028 ,n2813 ,n11[34]);
    nor g3297(n1027 ,n2923 ,n11[41]);
    nor g3298(n1026 ,n2823 ,n11[39]);
    nor g3299(n1025 ,n2921 ,n11[40]);
    nor g3300(n1024 ,n2879 ,n11[35]);
    nor g3301(n1023 ,n2857 ,n11[40]);
    nor g3302(n1022 ,n2907 ,n11[33]);
    nor g3303(n1021 ,n2927 ,n11[43]);
    nor g3304(n1020 ,n2811 ,n11[33]);
    nor g3305(n1019 ,n2839 ,n11[31]);
    nor g3306(n1018 ,n2881 ,n11[36]);
    nor g3307(n1017 ,n2873 ,n11[32]);
    nor g3308(n1016 ,n2887 ,n11[39]);
    nor g3309(n1015 ,n2899 ,n11[45]);
    nor g3310(n1014 ,n2847 ,n11[35]);
    nor g3311(n1013 ,n2867 ,n11[45]);
    nor g3312(n1012 ,n2901 ,n11[46]);
    nor g3313(n1011 ,n2913 ,n11[36]);
    nor g3314(n1010 ,n2845 ,n11[34]);
    nor g3315(n1009 ,n2905 ,n11[32]);
    nor g3316(n1008 ,n2919 ,n11[39]);
    nor g3317(n1007 ,n2821 ,n11[38]);
    nor g3318(n1006 ,n2863 ,n11[43]);
    nor g3319(n1005 ,n2865 ,n11[44]);
    nor g3320(n1004 ,n2925 ,n11[42]);
    nor g3321(n1003 ,n2833 ,n11[44]);
    nor g3322(n1002 ,n2861 ,n11[42]);
    nor g3323(n1001 ,n2883 ,n11[37]);
    nor g3324(n1000 ,n2931 ,n11[45]);
    nor g3325(n999 ,n2837 ,n11[46]);
    not g3326(n998 ,n2817);
    not g3327(n997 ,n2809);
    not g3328(n996 ,n2815);
    not g3329(n995 ,n11[42]);
    not g3330(n994 ,n11[40]);
    not g3331(n993 ,n2819);
    not g3332(n992 ,n2829);
    not g3333(n991 ,n2825);
    not g3334(n990 ,n10[49]);
    not g3335(n989 ,n11[36]);
    not g3336(n988 ,n11[35]);
    not g3337(n987 ,n11[37]);
    xor g3338(n2935 ,n12[2] ,n1255);
    nor g3339(n2936 ,n1255 ,n1254);
    nor g3340(n1255 ,n1253 ,n1252);
    nor g3341(n1254 ,n12[1] ,n12[0]);
    not g3342(n1253 ,n12[1]);
    not g3343(n1252 ,n12[0]);
    not g3344(n2940 ,n1);
    dff g3345(.RN(1'b1), .SN(n2940), .CK(n0), .D(n2939), .Q(n14[0]));
    xor g3346(n2939 ,n2938 ,n2937);
    xnor g3347(n2938 ,n10[60] ,n14[15]);
    xnor g3348(n2937 ,n14[10] ,n14[12]);
    dff g3349(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[9]), .Q(n10[57]));
    dff g3350(.RN(1'b1), .SN(n2940), .CK(n0), .D(n10[51]), .Q(n14[5]));
    dff g3351(.RN(n2940), .SN(1'b1), .CK(n0), .D(n10[48]), .Q(n10[49]));
    dff g3352(.RN(n2940), .SN(1'b1), .CK(n0), .D(n10[55]), .Q(n10[56]));
    dff g3353(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[11]), .Q(n10[59]));
    dff g3354(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[10]), .Q(n10[58]));
    dff g3355(.RN(n2940), .SN(1'b1), .CK(n0), .D(n10[60]), .Q(n10[61]));
    dff g3356(.RN(1'b1), .SN(n2940), .CK(n0), .D(n10[55]), .Q(n14[9]));
    dff g3357(.RN(1'b1), .SN(n2940), .CK(n0), .D(n10[60]), .Q(n14[14]));
    dff g3358(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[7]), .Q(n10[55]));
    dff g3359(.RN(1'b1), .SN(n2940), .CK(n0), .D(n14[11]), .Q(n14[12]));
    dff g3360(.RN(1'b1), .SN(n2940), .CK(n0), .D(n14[14]), .Q(n14[15]));
    dff g3361(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[0]), .Q(n10[48]));
    dff g3362(.RN(1'b1), .SN(n2940), .CK(n0), .D(n10[53]), .Q(n14[7]));
    dff g3363(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[15]), .Q(n10[47]));
    dff g3364(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[2]), .Q(n10[50]));
    dff g3365(.RN(n2940), .SN(1'b1), .CK(n0), .D(n10[51]), .Q(n10[52]));
    dff g3366(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[14]), .Q(n10[62]));
    dff g3367(.RN(n2940), .SN(1'b1), .CK(n0), .D(n10[53]), .Q(n10[54]));
    dff g3368(.RN(1'b1), .SN(n2940), .CK(n0), .D(n14[2]), .Q(n14[3]));
    dff g3369(.RN(1'b1), .SN(n2940), .CK(n0), .D(n10[48]), .Q(n14[2]));
    dff g3370(.RN(1'b1), .SN(n2940), .CK(n0), .D(n14[10]), .Q(n14[11]));
    dff g3371(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[5]), .Q(n10[53]));
    dff g3372(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[3]), .Q(n10[51]));
    dff g3373(.RN(1'b1), .SN(n2940), .CK(n0), .D(n14[9]), .Q(n14[10]));
    dff g3374(.RN(n2940), .SN(1'b1), .CK(n0), .D(n14[12]), .Q(n10[60]));
endmodule
