module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12);
    input n0, n1, n2, n3;
    input [1:0] n4, n5;
    output n6, n7;
    output [6:0] n8, n9;
    output [3:0] n10, n11, n12;
    wire n0, n1, n2, n3;
    wire [1:0] n4, n5;
    wire n6, n7;
    wire [6:0] n8, n9;
    wire [3:0] n10, n11, n12;
    wire [2:0] n13;
    wire [15:0] n14;
    wire n15, n16, n17, n18, n19, n20, n21, n22;
    wire n23, n24, n25, n26, n27, n28, n29, n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77;
    buf g0(n12[0], 1'b0);
    buf g1(n12[1], 1'b0);
    buf g2(n12[2], 1'b0);
    buf g3(n12[3], 1'b0);
    buf g4(n11[2], 1'b0);
    buf g5(n11[3], 1'b0);
    buf g6(n9[0], n8[6]);
    buf g7(n9[1], n8[6]);
    buf g8(n9[2], n8[6]);
    buf g9(n9[3], 1'b0);
    buf g10(n9[4], n8[6]);
    buf g11(n9[5], n8[6]);
    buf g12(n9[6], 1'b0);
    buf g13(n8[0], n8[6]);
    buf g14(n8[1], 1'b0);
    buf g15(n8[2], 1'b0);
    buf g16(n8[3], n8[6]);
    buf g17(n8[4], n8[6]);
    buf g18(n8[5], n8[6]);
    buf g19(n7, 1'b0);
    not g20(n28 ,n29);
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n27), .Q(n13[0]));
    nor g22(n27 ,n1 ,n26);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n24), .Q(n6));
    nor g24(n26 ,n13[0] ,n25);
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n13[0]), .Q(n8[6]));
    nor g26(n25 ,n22 ,n28);
    nor g27(n24 ,n23 ,n6);
    not g28(n23 ,n13[0]);
    not g29(n22 ,n2);
    nor g30(n11[1] ,n17 ,n21);
    nor g31(n11[0] ,n18 ,n21);
    nor g32(n21 ,n20 ,n19);
    or g33(n20 ,n10[3] ,n10[2]);
    or g34(n19 ,n10[1] ,n10[0]);
    not g35(n18 ,n14[4]);
    not g36(n17 ,n14[5]);
    or g37(n29 ,n16 ,n15);
    or g38(n16 ,n10[3] ,n10[2]);
    or g39(n15 ,n10[1] ,n10[0]);
    or g40(n14[5] ,n53 ,n77);
    xnor g41(n14[4] ,n59 ,n76);
    nor g42(n77 ,n52 ,n76);
    nor g43(n76 ,n64 ,n75);
    xnor g44(n10[3] ,n72 ,n74);
    nor g45(n75 ,n67 ,n74);
    xor g46(n10[2] ,n71 ,n69);
    nor g47(n74 ,n66 ,n73);
    nor g48(n73 ,n68 ,n70);
    nor g49(n72 ,n64 ,n67);
    nor g50(n71 ,n66 ,n68);
    nor g51(n10[1] ,n69 ,n65);
    not g52(n70 ,n69);
    nor g53(n69 ,n40 ,n60);
    nor g54(n68 ,n44 ,n58);
    nor g55(n67 ,n37 ,n63);
    nor g56(n66 ,n45 ,n57);
    nor g57(n65 ,n39 ,n61);
    nor g58(n64 ,n38 ,n62);
    not g59(n63 ,n62);
    nor g60(n62 ,n49 ,n56);
    not g61(n61 ,n60);
    nor g62(n60 ,n51 ,n55);
    nor g63(n59 ,n52 ,n53);
    not g64(n58 ,n57);
    nor g65(n57 ,n50 ,n54);
    nor g66(n56 ,n31 ,n46);
    nor g67(n55 ,n30 ,n46);
    nor g68(n10[0] ,n35 ,n46);
    nor g69(n54 ,n36 ,n46);
    nor g70(n53 ,n42 ,n48);
    nor g71(n52 ,n41 ,n47);
    nor g72(n51 ,n35 ,n43);
    nor g73(n50 ,n30 ,n43);
    nor g74(n49 ,n36 ,n43);
    not g75(n48 ,n47);
    nor g76(n47 ,n31 ,n43);
    xnor g77(n46 ,n13[0] ,n3);
    not g78(n45 ,n44);
    nor g79(n44 ,n30 ,n32);
    or g80(n43 ,n34 ,n33);
    not g81(n42 ,n41);
    nor g82(n41 ,n31 ,n32);
    not g83(n40 ,n39);
    nor g84(n39 ,n35 ,n32);
    not g85(n38 ,n37);
    nor g86(n37 ,n36 ,n32);
    not g87(n36 ,n4[0]);
    not g88(n35 ,n5[0]);
    not g89(n34 ,n3);
    not g90(n33 ,n13[0]);
    not g91(n32 ,n2);
    not g92(n31 ,n4[1]);
    not g93(n30 ,n5[1]);
endmodule
