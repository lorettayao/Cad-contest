module top(n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [3:0] n6;
    wire [2:0] n7;
    wire [3:0] n8;
    wire [31:0] n9;
    wire [31:0] n10;
    wire [31:0] n11;
    wire n12, n13, n14, n15, n16, n17, n18, n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
    wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
    wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627;
    wire n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635;
    wire n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643;
    wire n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
    wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
    wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
    wire n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675;
    wire n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683;
    wire n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
    wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
    wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707;
    wire n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715;
    wire n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723;
    wire n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
    wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
    wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
    wire n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755;
    wire n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763;
    wire n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
    wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
    wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787;
    wire n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795;
    wire n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803;
    wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
    wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
    wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
    wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
    wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
    wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
    wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
    wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
    wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
    wire n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883;
    wire n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
    wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
    wire n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907;
    wire n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915;
    wire n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923;
    wire n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931;
    wire n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939;
    wire n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947;
    wire n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955;
    wire n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963;
    wire n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
    wire n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979;
    wire n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987;
    wire n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995;
    wire n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;
    wire n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
    wire n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019;
    wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027;
    wire n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035;
    wire n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043;
    wire n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
    wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
    wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067;
    wire n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075;
    wire n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083;
    wire n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
    wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099;
    wire n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107;
    wire n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115;
    wire n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123;
    wire n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131;
    wire n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139;
    wire n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147;
    wire n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155;
    wire n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163;
    wire n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
    wire n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179;
    wire n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187;
    wire n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195;
    wire n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203;
    wire n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211;
    wire n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219;
    wire n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227;
    wire n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235;
    wire n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243;
    wire n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
    wire n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259;
    wire n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;
    wire n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275;
    wire n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283;
    wire n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291;
    wire n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299;
    wire n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307;
    wire n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315;
    wire n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323;
    wire n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331;
    wire n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339;
    wire n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347;
    wire n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355;
    wire n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363;
    wire n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371;
    wire n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379;
    wire n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387;
    wire n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395;
    wire n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403;
    wire n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411;
    wire n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419;
    wire n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427;
    wire n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435;
    wire n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443;
    wire n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451;
    wire n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459;
    wire n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467;
    wire n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475;
    wire n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483;
    wire n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491;
    wire n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499;
    wire n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507;
    wire n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515;
    wire n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523;
    wire n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531;
    wire n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539;
    wire n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547;
    wire n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555;
    wire n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563;
    wire n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571;
    wire n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579;
    wire n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587;
    wire n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595;
    wire n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603;
    wire n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;
    wire n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619;
    wire n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627;
    wire n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635;
    wire n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643;
    wire n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651;
    wire n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659;
    wire n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667;
    wire n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675;
    wire n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683;
    wire n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691;
    wire n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699;
    wire n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707;
    wire n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715;
    wire n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723;
    wire n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731;
    wire n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739;
    wire n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747;
    wire n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755;
    wire n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763;
    wire n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771;
    wire n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779;
    wire n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787;
    wire n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795;
    wire n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803;
    wire n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811;
    wire n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819;
    wire n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827;
    wire n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835;
    wire n2836, n2837, n2838, n2839, n2840, n2841, n2842;
    not g0(n2346 ,n1);
    or g1(n2482 ,n2260 ,n2345);
    or g2(n2481 ,n2256 ,n2344);
    or g3(n2480 ,n2252 ,n2343);
    or g4(n2479 ,n2268 ,n2342);
    nor g5(n2345 ,n2150 ,n2341);
    nor g6(n2344 ,n2150 ,n2340);
    nor g7(n2343 ,n2150 ,n2339);
    nor g8(n2342 ,n2150 ,n2338);
    or g9(n2483 ,n2234 ,n2320);
    or g10(n2517 ,n2276 ,n2334);
    or g11(n2491 ,n2275 ,n2335);
    or g12(n2490 ,n2274 ,n2332);
    or g13(n2516 ,n2245 ,n2329);
    or g14(n2489 ,n2272 ,n2331);
    or g15(n2529 ,n2269 ,n2326);
    or g16(n2515 ,n2225 ,n2327);
    or g17(n2488 ,n2270 ,n2330);
    or g18(n2487 ,n2217 ,n2328);
    or g19(n2514 ,n2266 ,n2322);
    or g20(n2486 ,n2267 ,n2325);
    or g21(n2535 ,n2257 ,n2313);
    or g22(n2485 ,n2265 ,n2323);
    or g23(n2484 ,n2263 ,n2321);
    or g24(n2528 ,n2262 ,n2318);
    or g25(n2536 ,n2271 ,n2324);
    or g26(n2513 ,n2261 ,n2319);
    or g27(n2542 ,n2241 ,n2316);
    or g28(n2527 ,n2255 ,n2314);
    or g29(n2512 ,n2258 ,n2317);
    or g30(n2541 ,n2264 ,n2308);
    or g31(n2539 ,n2259 ,n2311);
    or g32(n2511 ,n2254 ,n2315);
    or g33(n2534 ,n2273 ,n2304);
    or g34(n2510 ,n2251 ,n2312);
    or g35(n2526 ,n2249 ,n2309);
    or g36(n2538 ,n2230 ,n2301);
    or g37(n2509 ,n2248 ,n2310);
    or g38(n2508 ,n2247 ,n2307);
    or g39(n2525 ,n2244 ,n2337);
    or g40(n2507 ,n2243 ,n2306);
    or g41(n2537 ,n2220 ,n2280);
    or g42(n2524 ,n2240 ,n2299);
    or g43(n2505 ,n2239 ,n2302);
    or g44(n2540 ,n2223 ,n2305);
    or g45(n2533 ,n2238 ,n2296);
    or g46(n2523 ,n2236 ,n2297);
    or g47(n2504 ,n2237 ,n2300);
    or g48(n2503 ,n2235 ,n2298);
    or g49(n2522 ,n2232 ,n2294);
    or g50(n2502 ,n2233 ,n2295);
    or g51(n2532 ,n2228 ,n2285);
    or g52(n2501 ,n2231 ,n2293);
    or g53(n2500 ,n2229 ,n2292);
    or g54(n2521 ,n2227 ,n2290);
    or g55(n2499 ,n2226 ,n2291);
    or g56(n2498 ,n2224 ,n2289);
    or g57(n2506 ,n2242 ,n2303);
    or g58(n2531 ,n2218 ,n2282);
    or g59(n2520 ,n2222 ,n2287);
    or g60(n2497 ,n2221 ,n2288);
    or g61(n2519 ,n2253 ,n2283);
    or g62(n2496 ,n2219 ,n2286);
    or g63(n2495 ,n2246 ,n2284);
    or g64(n2530 ,n2277 ,n2333);
    or g65(n2518 ,n2215 ,n2278);
    or g66(n2494 ,n2216 ,n2281);
    or g67(n2493 ,n2250 ,n2279);
    or g68(n2492 ,n2214 ,n2336);
    xnor g69(n2341 ,n6[3] ,n2603);
    xnor g70(n2340 ,n6[2] ,n2604);
    xnor g71(n2339 ,n6[1] ,n2605);
    xnor g72(n2338 ,n6[0] ,n2606);
    nor g73(n2337 ,n2163 ,n2146);
    nor g74(n2336 ,n2185 ,n2150);
    nor g75(n2335 ,n2138 ,n2145);
    nor g76(n2334 ,n2192 ,n2146);
    nor g77(n2333 ,n2137 ,n2144);
    nor g78(n2332 ,n2209 ,n2147);
    nor g79(n2331 ,n2210 ,n2149);
    nor g80(n2330 ,n2175 ,n2148);
    nor g81(n2329 ,n2124 ,n2144);
    nor g82(n2328 ,n2199 ,n2145);
    nor g83(n2327 ,n2129 ,n2147);
    nor g84(n2326 ,n2190 ,n2144);
    nor g85(n2325 ,n2179 ,n2148);
    nor g86(n2324 ,n2184 ,n2143);
    nor g87(n2323 ,n2186 ,n2143);
    nor g88(n2322 ,n2202 ,n2146);
    nor g89(n2321 ,n2092 ,n2143);
    nor g90(n2320 ,n2188 ,n2143);
    nor g91(n2319 ,n2166 ,n2146);
    nor g92(n2318 ,n2168 ,n2143);
    nor g93(n2317 ,n2099 ,n2148);
    nor g94(n2316 ,n2123 ,n2144);
    nor g95(n2315 ,n2104 ,n2148);
    nor g96(n2314 ,n2094 ,n2147);
    nor g97(n2313 ,n2125 ,n2144);
    nor g98(n2312 ,n2206 ,n2150);
    nor g99(n2311 ,n2120 ,n2146);
    nor g100(n2310 ,n2085 ,n2147);
    nor g101(n2309 ,n2121 ,n2149);
    nor g102(n2308 ,n2157 ,n2147);
    nor g103(n2307 ,n2096 ,n2147);
    nor g104(n2306 ,n2117 ,n2146);
    nor g105(n2305 ,n2153 ,n2145);
    nor g106(n2304 ,n2160 ,n2150);
    nor g107(n2303 ,n2159 ,n2144);
    nor g108(n2302 ,n2113 ,n2148);
    nor g109(n2301 ,n2136 ,n2148);
    nor g110(n2300 ,n2132 ,n2148);
    nor g111(n2299 ,n2087 ,n2143);
    nor g112(n2298 ,n2177 ,n2143);
    nor g113(n2297 ,n2082 ,n2144);
    nor g114(n2296 ,n2212 ,n2149);
    nor g115(n2295 ,n2108 ,n2146);
    nor g116(n2294 ,n2130 ,n2147);
    nor g117(n2293 ,n2141 ,n2149);
    nor g118(n2292 ,n2205 ,n2146);
    nor g119(n2291 ,n2191 ,n2145);
    nor g120(n2290 ,n2196 ,n2144);
    nor g121(n2289 ,n2126 ,n2145);
    nor g122(n2288 ,n2122 ,n2143);
    nor g123(n2287 ,n2213 ,n2147);
    nor g124(n2286 ,n2211 ,n2145);
    nor g125(n2285 ,n2134 ,n2149);
    nor g126(n2284 ,n2170 ,n2150);
    nor g127(n2283 ,n2119 ,n2145);
    nor g128(n2282 ,n2165 ,n2145);
    nor g129(n2281 ,n2098 ,n2149);
    nor g130(n2280 ,n2086 ,n2148);
    nor g131(n2279 ,n2106 ,n2149);
    nor g132(n2278 ,n2103 ,n2149);
    nor g133(n2277 ,n2109 ,n2075);
    nor g134(n2276 ,n2083 ,n2077);
    nor g135(n2275 ,n2088 ,n2071);
    nor g136(n2274 ,n2115 ,n2074);
    nor g137(n2273 ,n2116 ,n2077);
    nor g138(n2272 ,n2140 ,n2074);
    nor g139(n2271 ,n2178 ,n2075);
    nor g140(n2270 ,n2101 ,n2077);
    nor g141(n2269 ,n2198 ,n2071);
    nor g142(n2268 ,n2139 ,n2074);
    nor g143(n2267 ,n2194 ,n2072);
    nor g144(n2266 ,n2128 ,n2077);
    nor g145(n2265 ,n2111 ,n2076);
    nor g146(n2476 ,n2079 ,n2072);
    nor g147(n2264 ,n2097 ,n2075);
    nor g148(n2263 ,n2183 ,n2076);
    nor g149(n2262 ,n2187 ,n2073);
    nor g150(n2261 ,n2176 ,n2070);
    nor g151(n2260 ,n2162 ,n2071);
    nor g152(n2259 ,n2180 ,n2070);
    nor g153(n2258 ,n2164 ,n2070);
    nor g154(n2257 ,n2093 ,n2073);
    nor g155(n2256 ,n2133 ,n2077);
    nor g156(n2255 ,n2193 ,n2070);
    nor g157(n2254 ,n2173 ,n2073);
    nor g158(n2253 ,n2112 ,n2073);
    nor g159(n2252 ,n2105 ,n2070);
    nor g160(n2478 ,n2078 ,n2073);
    nor g161(n2251 ,n2084 ,n2070);
    nor g162(n2250 ,n2100 ,n2073);
    nor g163(n2249 ,n2118 ,n2076);
    nor g164(n2248 ,n2208 ,n2072);
    nor g165(n2477 ,n2151 ,n2076);
    nor g166(n2475 ,n2080 ,n2074);
    nor g167(n2247 ,n2172 ,n2071);
    nor g168(n2246 ,n2171 ,n2075);
    nor g169(n2245 ,n2207 ,n2077);
    nor g170(n2244 ,n2095 ,n2076);
    nor g171(n2243 ,n2114 ,n2076);
    nor g172(n2242 ,n2161 ,n2077);
    nor g173(n2241 ,n2154 ,n2071);
    nor g174(n2240 ,n2102 ,n2075);
    nor g175(n2239 ,n2155 ,n2074);
    nor g176(n2238 ,n2089 ,n2072);
    nor g177(n2237 ,n2156 ,n2072);
    nor g178(n2236 ,n2110 ,n2072);
    nor g179(n2235 ,n2152 ,n2073);
    nor g180(n2234 ,n2174 ,n2077);
    nor g181(n2233 ,n2091 ,n2070);
    nor g182(n2232 ,n2107 ,n2075);
    nor g183(n2231 ,n2090 ,n2077);
    nor g184(n2230 ,n2142 ,n2077);
    nor g185(n2229 ,n2135 ,n2076);
    nor g186(n2228 ,n2195 ,n2077);
    nor g187(n2227 ,n2201 ,n2071);
    nor g188(n2226 ,n2200 ,n2074);
    nor g189(n2225 ,n2204 ,n2074);
    nor g190(n2224 ,n2197 ,n2073);
    nor g191(n2223 ,n2081 ,n2071);
    nor g192(n2222 ,n2182 ,n2072);
    nor g193(n2221 ,n2189 ,n2076);
    nor g194(n2220 ,n2158 ,n2075);
    nor g195(n2219 ,n2181 ,n2074);
    nor g196(n2218 ,n2167 ,n2070);
    nor g197(n2217 ,n2203 ,n2071);
    nor g198(n2216 ,n2169 ,n2072);
    nor g199(n2215 ,n2127 ,n2075);
    nor g200(n2214 ,n2131 ,n2077);
    not g201(n2213 ,n2580);
    not g202(n2212 ,n2593);
    not g203(n2211 ,n2556);
    not g204(n2210 ,n2549);
    not g205(n2209 ,n2550);
    not g206(n2208 ,n3[30]);
    not g207(n2207 ,n3[37]);
    not g208(n2206 ,n2570);
    not g209(n2205 ,n2560);
    not g210(n2204 ,n3[36]);
    not g211(n2203 ,n3[8]);
    not g212(n2202 ,n2574);
    not g213(n2201 ,n3[42]);
    not g214(n2200 ,n3[20]);
    not g215(n2199 ,n2547);
    not g216(n2198 ,n3[50]);
    not g217(n2197 ,n3[19]);
    not g218(n2196 ,n2581);
    not g219(n2195 ,n3[53]);
    not g220(n2194 ,n3[7]);
    not g221(n2193 ,n3[48]);
    not g222(n2192 ,n2577);
    not g223(n2191 ,n2559);
    not g224(n2190 ,n2589);
    not g225(n2189 ,n3[18]);
    not g226(n2188 ,n2543);
    not g227(n2187 ,n3[49]);
    not g228(n2186 ,n2545);
    not g229(n2185 ,n2552);
    not g230(n2184 ,n2596);
    not g231(n2183 ,n3[5]);
    not g232(n2182 ,n3[41]);
    not g233(n2181 ,n3[17]);
    not g234(n2180 ,n3[60]);
    not g235(n2179 ,n2546);
    not g236(n2178 ,n3[57]);
    not g237(n2177 ,n2563);
    not g238(n2176 ,n3[34]);
    not g239(n2175 ,n2548);
    not g240(n2174 ,n3[4]);
    not g241(n2173 ,n3[32]);
    not g242(n2172 ,n3[29]);
    not g243(n2171 ,n3[16]);
    not g244(n2170 ,n2555);
    not g245(n2169 ,n3[15]);
    not g246(n2168 ,n2588);
    not g247(n2167 ,n3[52]);
    not g248(n2166 ,n2573);
    not g249(n2165 ,n2591);
    not g250(n2164 ,n3[33]);
    not g251(n2163 ,n2585);
    not g252(n2162 ,n3[3]);
    not g253(n2161 ,n3[27]);
    not g254(n2160 ,n2594);
    not g255(n2159 ,n2566);
    not g256(n2158 ,n3[58]);
    not g257(n2157 ,n2601);
    not g258(n2156 ,n3[25]);
    not g259(n2155 ,n3[26]);
    not g260(n2154 ,n3[63]);
    not g261(n2153 ,n2600);
    not g262(n2152 ,n3[24]);
    not g263(n2151 ,n6[2]);
    not g264(n2150 ,n7[1]);
    not g265(n2149 ,n7[1]);
    not g266(n2148 ,n7[1]);
    not g267(n2147 ,n7[1]);
    not g268(n2146 ,n7[1]);
    not g269(n2145 ,n7[1]);
    not g270(n2144 ,n7[1]);
    not g271(n2143 ,n7[1]);
    not g272(n2142 ,n3[59]);
    not g273(n2141 ,n2561);
    not g274(n2140 ,n3[10]);
    not g275(n2139 ,n3[0]);
    not g276(n2138 ,n2551);
    not g277(n2137 ,n2590);
    not g278(n2136 ,n2598);
    not g279(n2135 ,n3[21]);
    not g280(n2134 ,n2592);
    not g281(n2133 ,n3[2]);
    not g282(n2132 ,n2564);
    not g283(n2131 ,n3[13]);
    not g284(n2130 ,n2582);
    not g285(n2129 ,n2575);
    not g286(n2128 ,n3[35]);
    not g287(n2127 ,n3[39]);
    not g288(n2126 ,n2558);
    not g289(n2125 ,n2595);
    not g290(n2124 ,n2576);
    not g291(n2123 ,n2602);
    not g292(n2122 ,n2557);
    not g293(n2121 ,n2586);
    not g294(n2120 ,n2599);
    not g295(n2119 ,n2579);
    not g296(n2118 ,n3[47]);
    not g297(n2117 ,n2567);
    not g298(n2116 ,n3[55]);
    not g299(n2115 ,n3[11]);
    not g300(n2114 ,n3[28]);
    not g301(n2113 ,n2565);
    not g302(n2112 ,n3[40]);
    not g303(n2111 ,n3[6]);
    not g304(n2110 ,n3[44]);
    not g305(n2109 ,n3[51]);
    not g306(n2108 ,n2562);
    not g307(n2107 ,n3[43]);
    not g308(n2106 ,n2553);
    not g309(n2105 ,n3[1]);
    not g310(n2104 ,n2571);
    not g311(n2103 ,n2578);
    not g312(n2102 ,n3[45]);
    not g313(n2101 ,n3[9]);
    not g314(n2100 ,n3[14]);
    not g315(n2099 ,n2572);
    not g316(n2098 ,n2554);
    not g317(n2097 ,n3[62]);
    not g318(n2096 ,n2568);
    not g319(n2095 ,n3[46]);
    not g320(n2094 ,n2587);
    not g321(n2093 ,n3[56]);
    not g322(n2092 ,n2544);
    not g323(n2091 ,n3[23]);
    not g324(n2090 ,n3[22]);
    not g325(n2089 ,n3[54]);
    not g326(n2088 ,n3[12]);
    not g327(n2087 ,n2584);
    not g328(n2086 ,n2597);
    not g329(n2085 ,n2569);
    not g330(n2084 ,n3[31]);
    not g331(n2083 ,n3[38]);
    not g332(n2082 ,n2583);
    not g333(n2081 ,n3[61]);
    not g334(n2080 ,n6[0]);
    not g335(n2079 ,n6[1]);
    not g336(n2078 ,n6[3]);
    not g337(n2077 ,n7[2]);
    not g338(n2076 ,n7[2]);
    not g339(n2075 ,n7[2]);
    not g340(n2074 ,n7[2]);
    not g341(n2073 ,n7[2]);
    not g342(n2072 ,n7[2]);
    not g343(n2071 ,n7[2]);
    not g344(n2070 ,n7[2]);
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2065), .Q(n5[0]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n5[1]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2064), .Q(n5[2]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2066), .Q(n5[3]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1891), .Q(n5[4]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n5[5]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1890), .Q(n5[6]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1888), .Q(n5[7]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n5[8]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n5[9]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1885), .Q(n5[10]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n5[11]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n5[12]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n5[13]));
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n5[14]));
    dff g360(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n5[15]));
    dff g361(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n5[16]));
    dff g362(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n5[17]));
    dff g363(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n5[18]));
    dff g364(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n5[19]));
    dff g365(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n5[20]));
    dff g366(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n5[21]));
    dff g367(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n5[22]));
    dff g368(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n5[23]));
    dff g369(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n5[24]));
    dff g370(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n5[25]));
    dff g371(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n5[26]));
    dff g372(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n5[27]));
    dff g373(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n5[28]));
    dff g374(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n5[29]));
    dff g375(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n5[30]));
    dff g376(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n5[31]));
    dff g377(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n5[32]));
    dff g378(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n5[33]));
    dff g379(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n5[34]));
    dff g380(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n5[35]));
    dff g381(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n5[36]));
    dff g382(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n5[37]));
    dff g383(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1852), .Q(n5[38]));
    dff g384(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1851), .Q(n5[39]));
    dff g385(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n5[40]));
    dff g386(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n5[41]));
    dff g387(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n5[42]));
    dff g388(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n5[43]));
    dff g389(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n5[44]));
    dff g390(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n5[45]));
    dff g391(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n5[46]));
    dff g392(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n5[47]));
    dff g393(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n5[48]));
    dff g394(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n5[49]));
    dff g395(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n5[50]));
    dff g396(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n5[51]));
    dff g397(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n5[52]));
    dff g398(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n5[53]));
    dff g399(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1837), .Q(n5[54]));
    dff g400(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1835), .Q(n5[55]));
    dff g401(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1834), .Q(n5[56]));
    dff g402(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n5[57]));
    dff g403(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n5[58]));
    dff g404(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n5[59]));
    dff g405(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n5[60]));
    dff g406(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n5[61]));
    dff g407(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n5[62]));
    dff g408(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n5[63]));
    dff g409(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1036), .Q(n8[0]));
    dff g410(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1039), .Q(n8[1]));
    dff g411(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1043), .Q(n8[2]));
    dff g412(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1040), .Q(n8[3]));
    dff g413(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2059), .Q(n3[0]));
    dff g414(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2063), .Q(n3[1]));
    dff g415(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2058), .Q(n3[2]));
    dff g416(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2052), .Q(n3[3]));
    dff g417(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n3[4]));
    dff g418(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n3[5]));
    dff g419(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n3[6]));
    dff g420(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n3[7]));
    dff g421(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1908), .Q(n3[8]));
    dff g422(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n3[9]));
    dff g423(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n3[10]));
    dff g424(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n3[11]));
    dff g425(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1904), .Q(n3[12]));
    dff g426(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n3[13]));
    dff g427(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1902), .Q(n3[14]));
    dff g428(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1901), .Q(n3[15]));
    dff g429(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1900), .Q(n3[16]));
    dff g430(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1899), .Q(n3[17]));
    dff g431(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n3[18]));
    dff g432(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n3[19]));
    dff g433(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n3[20]));
    dff g434(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n3[21]));
    dff g435(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n3[22]));
    dff g436(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n3[23]));
    dff g437(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n3[24]));
    dff g438(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n3[25]));
    dff g439(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n3[26]));
    dff g440(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n3[27]));
    dff g441(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n3[28]));
    dff g442(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n3[29]));
    dff g443(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n3[30]));
    dff g444(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n3[31]));
    dff g445(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n3[32]));
    dff g446(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n3[33]));
    dff g447(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n3[34]));
    dff g448(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n3[35]));
    dff g449(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n3[36]));
    dff g450(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n3[37]));
    dff g451(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n3[38]));
    dff g452(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n3[39]));
    dff g453(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n3[40]));
    dff g454(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n3[41]));
    dff g455(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n3[42]));
    dff g456(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n3[43]));
    dff g457(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n3[44]));
    dff g458(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n3[45]));
    dff g459(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n3[46]));
    dff g460(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n3[47]));
    dff g461(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n3[48]));
    dff g462(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n3[49]));
    dff g463(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n3[50]));
    dff g464(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n3[51]));
    dff g465(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n3[52]));
    dff g466(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n3[53]));
    dff g467(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n3[54]));
    dff g468(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n3[55]));
    dff g469(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n3[56]));
    dff g470(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n3[57]));
    dff g471(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n3[58]));
    dff g472(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n3[59]));
    dff g473(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n3[60]));
    dff g474(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n3[61]));
    dff g475(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n3[62]));
    dff g476(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n3[63]));
    dff g477(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1088), .Q(n9[0]));
    dff g478(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1087), .Q(n9[1]));
    dff g479(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1086), .Q(n9[2]));
    dff g480(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1085), .Q(n9[3]));
    dff g481(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1105), .Q(n9[4]));
    dff g482(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1084), .Q(n9[5]));
    dff g483(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1083), .Q(n9[6]));
    dff g484(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1082), .Q(n9[7]));
    dff g485(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1108), .Q(n9[8]));
    dff g486(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1081), .Q(n9[9]));
    dff g487(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1080), .Q(n9[10]));
    dff g488(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1079), .Q(n9[11]));
    dff g489(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1044), .Q(n9[12]));
    dff g490(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1078), .Q(n9[13]));
    dff g491(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1077), .Q(n9[14]));
    dff g492(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1076), .Q(n9[15]));
    dff g493(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1045), .Q(n9[16]));
    dff g494(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1075), .Q(n9[17]));
    dff g495(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1074), .Q(n9[18]));
    dff g496(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1071), .Q(n9[19]));
    dff g497(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1047), .Q(n9[20]));
    dff g498(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1070), .Q(n9[21]));
    dff g499(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1069), .Q(n9[22]));
    dff g500(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1068), .Q(n9[23]));
    dff g501(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1049), .Q(n9[24]));
    dff g502(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1067), .Q(n9[25]));
    dff g503(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1066), .Q(n9[26]));
    dff g504(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1065), .Q(n9[27]));
    dff g505(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1052), .Q(n9[28]));
    dff g506(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1064), .Q(n9[29]));
    dff g507(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1058), .Q(n9[30]));
    dff g508(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1063), .Q(n9[31]));
    dff g509(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2050), .Q(n7[0]));
    dff g510(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2051), .Q(n2068));
    dff g511(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n2069));
    dff g512(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2057), .Q(n4[0]));
    dff g513(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n4[1]));
    dff g514(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2061), .Q(n4[2]));
    dff g515(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2060), .Q(n4[3]));
    dff g516(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n4[4]));
    dff g517(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n4[5]));
    dff g518(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n4[6]));
    dff g519(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n4[7]));
    dff g520(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n4[8]));
    dff g521(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n4[9]));
    dff g522(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n4[10]));
    dff g523(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n4[11]));
    dff g524(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n4[12]));
    dff g525(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n4[13]));
    dff g526(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n4[14]));
    dff g527(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n4[15]));
    dff g528(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n4[16]));
    dff g529(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n4[17]));
    dff g530(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n4[18]));
    dff g531(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n4[19]));
    dff g532(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n4[20]));
    dff g533(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n4[21]));
    dff g534(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n4[22]));
    dff g535(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n4[23]));
    dff g536(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n4[24]));
    dff g537(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n4[25]));
    dff g538(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1950), .Q(n4[26]));
    dff g539(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n4[27]));
    dff g540(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n4[28]));
    dff g541(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1946), .Q(n4[29]));
    dff g542(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1945), .Q(n4[30]));
    dff g543(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n4[31]));
    dff g544(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1943), .Q(n4[32]));
    dff g545(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1942), .Q(n4[33]));
    dff g546(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1941), .Q(n4[34]));
    dff g547(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1940), .Q(n4[35]));
    dff g548(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1939), .Q(n4[36]));
    dff g549(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1938), .Q(n4[37]));
    dff g550(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1937), .Q(n4[38]));
    dff g551(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1936), .Q(n4[39]));
    dff g552(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n4[40]));
    dff g553(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n4[41]));
    dff g554(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n4[42]));
    dff g555(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n4[43]));
    dff g556(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n4[44]));
    dff g557(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n4[45]));
    dff g558(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2033), .Q(n4[46]));
    dff g559(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n4[47]));
    dff g560(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n4[48]));
    dff g561(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n4[49]));
    dff g562(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n4[50]));
    dff g563(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1924), .Q(n4[51]));
    dff g564(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1923), .Q(n4[52]));
    dff g565(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1922), .Q(n4[53]));
    dff g566(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1921), .Q(n4[54]));
    dff g567(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n4[55]));
    dff g568(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n4[56]));
    dff g569(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1919), .Q(n4[57]));
    dff g570(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n4[58]));
    dff g571(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1917), .Q(n4[59]));
    dff g572(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n4[60]));
    dff g573(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1915), .Q(n4[61]));
    dff g574(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1914), .Q(n4[62]));
    dff g575(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n4[63]));
    dff g576(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1090), .Q(n10[28]));
    dff g577(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1091), .Q(n10[29]));
    dff g578(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1048), .Q(n10[30]));
    dff g579(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1099), .Q(n10[31]));
    dff g580(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1094), .Q(n11[0]));
    dff g581(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1057), .Q(n11[1]));
    dff g582(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1042), .Q(n11[2]));
    dff g583(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1095), .Q(n11[3]));
    dff g584(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1096), .Q(n11[4]));
    dff g585(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1092), .Q(n11[5]));
    dff g586(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1051), .Q(n11[6]));
    dff g587(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1102), .Q(n11[7]));
    dff g588(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1053), .Q(n11[8]));
    dff g589(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1103), .Q(n11[9]));
    dff g590(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1055), .Q(n11[10]));
    dff g591(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1104), .Q(n11[11]));
    dff g592(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1110), .Q(n11[12]));
    dff g593(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1107), .Q(n11[13]));
    dff g594(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1059), .Q(n11[14]));
    dff g595(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1109), .Q(n11[15]));
    dff g596(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1062), .Q(n11[16]));
    dff g597(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1061), .Q(n11[17]));
    dff g598(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1041), .Q(n11[18]));
    dff g599(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1046), .Q(n11[19]));
    dff g600(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1038), .Q(n11[20]));
    dff g601(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1106), .Q(n11[21]));
    dff g602(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1089), .Q(n11[22]));
    dff g603(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1054), .Q(n11[23]));
    dff g604(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1097), .Q(n11[24]));
    dff g605(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1101), .Q(n11[25]));
    dff g606(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1060), .Q(n11[26]));
    dff g607(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1093), .Q(n11[27]));
    dff g608(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1050), .Q(n11[28]));
    dff g609(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1056), .Q(n11[29]));
    dff g610(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1098), .Q(n11[30]));
    dff g611(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1100), .Q(n11[31]));
    or g612(n2067 ,n1761 ,n2054);
    or g613(n2066 ,n1759 ,n2056);
    or g614(n2065 ,n1762 ,n2055);
    or g615(n2064 ,n2023 ,n2053);
    or g616(n2063 ,n2046 ,n1825);
    or g617(n2062 ,n2042 ,n1864);
    or g618(n2061 ,n2043 ,n1861);
    or g619(n2060 ,n2044 ,n1859);
    or g620(n2059 ,n2045 ,n1826);
    or g621(n2058 ,n2047 ,n1870);
    or g622(n2057 ,n2041 ,n1867);
    or g623(n2056 ,n2022 ,n2037);
    or g624(n2055 ,n2025 ,n2035);
    or g625(n2054 ,n2024 ,n2034);
    or g626(n2053 ,n1760 ,n2036);
    or g627(n2052 ,n2048 ,n1928);
    nor g628(n2051 ,n552 ,n2039);
    nor g629(n2050 ,n550 ,n2038);
    nor g630(n2049 ,n550 ,n2040);
    or g631(n2048 ,n1586 ,n2026);
    or g632(n2047 ,n1591 ,n2027);
    or g633(n2046 ,n1596 ,n2028);
    or g634(n2045 ,n1603 ,n2029);
    or g635(n2044 ,n1652 ,n2030);
    or g636(n2043 ,n1653 ,n2031);
    or g637(n2042 ,n1654 ,n2032);
    or g638(n2041 ,n1655 ,n1929);
    nor g639(n2040 ,n2020 ,n1973);
    nor g640(n2039 ,n2021 ,n1974);
    nor g641(n2038 ,n2019 ,n1975);
    nor g642(n2037 ,n1127 ,n1991);
    nor g643(n2036 ,n1128 ,n1993);
    nor g644(n2035 ,n1129 ,n2002);
    nor g645(n2034 ,n1130 ,n1999);
    or g646(n2033 ,n1607 ,n1461);
    nor g647(n2032 ,n820 ,n1625);
    nor g648(n2031 ,n823 ,n1625);
    nor g649(n2030 ,n826 ,n1625);
    nor g650(n2029 ,n828 ,n1624);
    nor g651(n2028 ,n827 ,n1624);
    nor g652(n2027 ,n829 ,n1624);
    nor g653(n2026 ,n818 ,n1624);
    nor g654(n2025 ,n822 ,n1627);
    nor g655(n2024 ,n825 ,n1627);
    nor g656(n2023 ,n824 ,n1627);
    nor g657(n2022 ,n821 ,n1627);
    nor g658(n2021 ,n528 ,n1622);
    nor g659(n2020 ,n817 ,n1622);
    nor g660(n2019 ,n816 ,n1622);
    or g661(n2018 ,n1699 ,n1546);
    or g662(n2017 ,n1697 ,n1545);
    or g663(n2016 ,n1696 ,n1544);
    or g664(n2015 ,n1695 ,n1543);
    or g665(n2014 ,n1694 ,n1542);
    or g666(n2013 ,n1692 ,n1539);
    or g667(n2012 ,n1693 ,n1541);
    or g668(n2011 ,n1691 ,n1538);
    or g669(n2010 ,n1690 ,n1537);
    or g670(n2009 ,n1689 ,n1536);
    or g671(n2008 ,n1687 ,n1535);
    or g672(n2007 ,n1686 ,n1534);
    or g673(n2006 ,n1685 ,n1532);
    or g674(n2005 ,n1684 ,n1529);
    or g675(n2004 ,n1683 ,n1528);
    or g676(n2003 ,n1682 ,n1527);
    or g677(n2002 ,n1033 ,n1626);
    or g678(n2001 ,n1681 ,n1525);
    or g679(n2000 ,n1680 ,n1621);
    or g680(n1999 ,n1037 ,n1626);
    or g681(n1998 ,n1679 ,n1522);
    or g682(n1997 ,n1678 ,n1520);
    or g683(n1996 ,n1677 ,n1519);
    or g684(n1995 ,n1676 ,n1518);
    or g685(n1994 ,n1675 ,n1517);
    or g686(n1993 ,n1032 ,n1626);
    or g687(n1992 ,n1673 ,n1516);
    or g688(n1991 ,n1025 ,n1626);
    or g689(n1990 ,n1672 ,n1515);
    or g690(n1989 ,n1671 ,n1513);
    or g691(n1988 ,n1670 ,n1512);
    or g692(n1987 ,n1669 ,n1511);
    or g693(n1986 ,n1668 ,n1510);
    or g694(n1985 ,n1666 ,n1509);
    or g695(n1984 ,n1665 ,n1507);
    or g696(n1983 ,n1664 ,n1505);
    or g697(n1982 ,n1663 ,n1504);
    or g698(n1981 ,n1662 ,n1502);
    or g699(n1980 ,n1661 ,n1501);
    or g700(n1979 ,n1660 ,n1500);
    or g701(n1978 ,n1659 ,n1499);
    or g702(n1977 ,n1658 ,n1497);
    or g703(n1976 ,n1657 ,n1496);
    nor g704(n1975 ,n1016 ,n1623);
    nor g705(n1974 ,n1134 ,n1623);
    nor g706(n1973 ,n1014 ,n1623);
    or g707(n1972 ,n1651 ,n1487);
    or g708(n1971 ,n1650 ,n1486);
    or g709(n1970 ,n1649 ,n1485);
    or g710(n1969 ,n1648 ,n1484);
    or g711(n1968 ,n1647 ,n1481);
    or g712(n1967 ,n1646 ,n1488);
    or g713(n1966 ,n1645 ,n1483);
    or g714(n1965 ,n1644 ,n1482);
    or g715(n1964 ,n1643 ,n1506);
    or g716(n1963 ,n1642 ,n1498);
    or g717(n1962 ,n1641 ,n1479);
    or g718(n1961 ,n1640 ,n1477);
    or g719(n1960 ,n1639 ,n1436);
    or g720(n1959 ,n1637 ,n1444);
    or g721(n1958 ,n1638 ,n1478);
    or g722(n1957 ,n1636 ,n1476);
    or g723(n1956 ,n1635 ,n1475);
    or g724(n1955 ,n1634 ,n1459);
    or g725(n1954 ,n1633 ,n1465);
    or g726(n1953 ,n1632 ,n1474);
    or g727(n1952 ,n1631 ,n1473);
    or g728(n1951 ,n1667 ,n1495);
    or g729(n1950 ,n1629 ,n1470);
    or g730(n1949 ,n1630 ,n1471);
    or g731(n1948 ,n1823 ,n1469);
    or g732(n1947 ,n1656 ,n1492);
    or g733(n1946 ,n1523 ,n1503);
    or g734(n1945 ,n1620 ,n1508);
    or g735(n1944 ,n1619 ,n1514);
    or g736(n1943 ,n1688 ,n1526);
    or g737(n1942 ,n1618 ,n1524);
    or g738(n1941 ,n1617 ,n1540);
    or g739(n1940 ,n1616 ,n1467);
    or g740(n1939 ,n1615 ,n1466);
    or g741(n1938 ,n1614 ,n1533);
    or g742(n1937 ,n1613 ,n1456);
    or g743(n1936 ,n1612 ,n1489);
    or g744(n1935 ,n1674 ,n1521);
    or g745(n1934 ,n1611 ,n1553);
    or g746(n1933 ,n1610 ,n1432);
    or g747(n1932 ,n1609 ,n1464);
    or g748(n1931 ,n1597 ,n1452);
    or g749(n1930 ,n1608 ,n1462);
    nor g750(n1929 ,n819 ,n1625);
    or g751(n1928 ,n1549 ,n1548);
    or g752(n1927 ,n1605 ,n1463);
    or g753(n1926 ,n1604 ,n1458);
    or g754(n1925 ,n1602 ,n1493);
    or g755(n1924 ,n1601 ,n1457);
    or g756(n1923 ,n1600 ,n1468);
    or g757(n1922 ,n1599 ,n1455);
    or g758(n1921 ,n1598 ,n1472);
    or g759(n1920 ,n1595 ,n1480);
    or g760(n1919 ,n1594 ,n1454);
    or g761(n1918 ,n1593 ,n1453);
    or g762(n1917 ,n1592 ,n1451);
    or g763(n1916 ,n1590 ,n1490);
    or g764(n1915 ,n1589 ,n1494);
    or g765(n1914 ,n1588 ,n1450);
    or g766(n1913 ,n1587 ,n1449);
    or g767(n1912 ,n1584 ,n1447);
    or g768(n1911 ,n1583 ,n1446);
    or g769(n1910 ,n1582 ,n1445);
    or g770(n1909 ,n1585 ,n1448);
    or g771(n1908 ,n1581 ,n1443);
    or g772(n1907 ,n1580 ,n1442);
    or g773(n1906 ,n1579 ,n1441);
    or g774(n1905 ,n1578 ,n1440);
    or g775(n1904 ,n1577 ,n1439);
    or g776(n1903 ,n1576 ,n1438);
    or g777(n1902 ,n1575 ,n1437);
    or g778(n1901 ,n1574 ,n1435);
    or g779(n1900 ,n1573 ,n1434);
    or g780(n1899 ,n1572 ,n1433);
    or g781(n1898 ,n1571 ,n1431);
    or g782(n1897 ,n1570 ,n1430);
    or g783(n1896 ,n1569 ,n1491);
    or g784(n1895 ,n1568 ,n1530);
    or g785(n1894 ,n1567 ,n1531);
    or g786(n1893 ,n1566 ,n1565);
    or g787(n1892 ,n1698 ,n1547);
    or g788(n1891 ,n1628 ,n1758);
    or g789(n1890 ,n1821 ,n1756);
    or g790(n1889 ,n1822 ,n1757);
    or g791(n1888 ,n1820 ,n1755);
    or g792(n1887 ,n1819 ,n1754);
    or g793(n1886 ,n1818 ,n1753);
    or g794(n1885 ,n1817 ,n1752);
    or g795(n1884 ,n1816 ,n1751);
    or g796(n1883 ,n1815 ,n1750);
    or g797(n1882 ,n1814 ,n1749);
    or g798(n1881 ,n1813 ,n1748);
    or g799(n1880 ,n1812 ,n1747);
    or g800(n1879 ,n1811 ,n1746);
    or g801(n1878 ,n1810 ,n1745);
    or g802(n1877 ,n1808 ,n1743);
    or g803(n1876 ,n1809 ,n1744);
    or g804(n1875 ,n1807 ,n1742);
    or g805(n1874 ,n1805 ,n1740);
    or g806(n1873 ,n1806 ,n1741);
    or g807(n1872 ,n1804 ,n1739);
    or g808(n1871 ,n1803 ,n1738);
    or g809(n1870 ,n1551 ,n1550);
    or g810(n1869 ,n1802 ,n1737);
    or g811(n1868 ,n1801 ,n1736);
    or g812(n1867 ,n1564 ,n1563);
    or g813(n1866 ,n1800 ,n1735);
    or g814(n1865 ,n1799 ,n1734);
    or g815(n1864 ,n1562 ,n1561);
    or g816(n1863 ,n1798 ,n1733);
    or g817(n1862 ,n1797 ,n1732);
    or g818(n1861 ,n1560 ,n1559);
    or g819(n1860 ,n1796 ,n1731);
    or g820(n1859 ,n1556 ,n1555);
    or g821(n1858 ,n1795 ,n1730);
    or g822(n1857 ,n1793 ,n1728);
    or g823(n1856 ,n1792 ,n1727);
    or g824(n1855 ,n1791 ,n1726);
    or g825(n1854 ,n1794 ,n1729);
    or g826(n1853 ,n1790 ,n1725);
    or g827(n1852 ,n1789 ,n1724);
    or g828(n1851 ,n1788 ,n1723);
    or g829(n1850 ,n1787 ,n1722);
    or g830(n1849 ,n1786 ,n1721);
    or g831(n1848 ,n1785 ,n1720);
    or g832(n1847 ,n1784 ,n1719);
    or g833(n1846 ,n1783 ,n1718);
    or g834(n1845 ,n1782 ,n1717);
    or g835(n1844 ,n1781 ,n1716);
    or g836(n1843 ,n1780 ,n1715);
    or g837(n1842 ,n1779 ,n1714);
    or g838(n1841 ,n1777 ,n1713);
    or g839(n1840 ,n1778 ,n1712);
    or g840(n1839 ,n1776 ,n1711);
    or g841(n1838 ,n1775 ,n1710);
    or g842(n1837 ,n1773 ,n1708);
    or g843(n1836 ,n1774 ,n1709);
    or g844(n1835 ,n1772 ,n1707);
    or g845(n1834 ,n1771 ,n1763);
    or g846(n1833 ,n1770 ,n1706);
    or g847(n1832 ,n1769 ,n1705);
    or g848(n1831 ,n1768 ,n1704);
    or g849(n1830 ,n1767 ,n1703);
    or g850(n1829 ,n1766 ,n1702);
    or g851(n1828 ,n1765 ,n1701);
    or g852(n1827 ,n1764 ,n1700);
    or g853(n1826 ,n1554 ,n1552);
    or g854(n1825 ,n1558 ,n1557);
    or g855(n1824 ,n1606 ,n1460);
    nor g856(n1823 ,n798 ,n536);
    nor g857(n1822 ,n878 ,n540);
    nor g858(n1821 ,n850 ,n541);
    nor g859(n1820 ,n916 ,n540);
    nor g860(n1819 ,n911 ,n541);
    nor g861(n1818 ,n1012 ,n541);
    nor g862(n1817 ,n972 ,n541);
    nor g863(n1816 ,n903 ,n540);
    nor g864(n1815 ,n926 ,n540);
    nor g865(n1814 ,n887 ,n541);
    nor g866(n1813 ,n919 ,n541);
    nor g867(n1812 ,n948 ,n540);
    nor g868(n1811 ,n867 ,n541);
    nor g869(n1810 ,n939 ,n540);
    nor g870(n1809 ,n894 ,n540);
    nor g871(n1808 ,n996 ,n541);
    nor g872(n1807 ,n922 ,n540);
    nor g873(n1806 ,n866 ,n540);
    nor g874(n1805 ,n930 ,n541);
    nor g875(n1804 ,n950 ,n541);
    nor g876(n1803 ,n862 ,n540);
    nor g877(n1802 ,n994 ,n541);
    nor g878(n1801 ,n833 ,n540);
    nor g879(n1800 ,n963 ,n540);
    nor g880(n1799 ,n1011 ,n540);
    nor g881(n1798 ,n1000 ,n540);
    nor g882(n1797 ,n966 ,n541);
    nor g883(n1796 ,n899 ,n541);
    nor g884(n1795 ,n844 ,n540);
    nor g885(n1794 ,n1007 ,n541);
    nor g886(n1793 ,n965 ,n541);
    nor g887(n1792 ,n988 ,n541);
    nor g888(n1791 ,n990 ,n541);
    nor g889(n1790 ,n979 ,n540);
    nor g890(n1789 ,n947 ,n541);
    nor g891(n1788 ,n923 ,n540);
    nor g892(n1787 ,n918 ,n540);
    nor g893(n1786 ,n863 ,n540);
    nor g894(n1785 ,n888 ,n540);
    nor g895(n1784 ,n974 ,n540);
    nor g896(n1783 ,n1008 ,n540);
    nor g897(n1782 ,n875 ,n541);
    nor g898(n1781 ,n845 ,n541);
    nor g899(n1780 ,n949 ,n541);
    nor g900(n1779 ,n959 ,n540);
    nor g901(n1778 ,n978 ,n541);
    nor g902(n1777 ,n968 ,n541);
    nor g903(n1776 ,n882 ,n540);
    nor g904(n1775 ,n914 ,n540);
    nor g905(n1774 ,n924 ,n540);
    nor g906(n1773 ,n1004 ,n540);
    nor g907(n1772 ,n910 ,n541);
    nor g908(n1771 ,n989 ,n540);
    nor g909(n1770 ,n889 ,n541);
    nor g910(n1769 ,n951 ,n541);
    nor g911(n1768 ,n995 ,n540);
    nor g912(n1767 ,n855 ,n541);
    nor g913(n1766 ,n851 ,n540);
    nor g914(n1765 ,n836 ,n540);
    nor g915(n1764 ,n946 ,n540);
    nor g916(n1763 ,n581 ,n539);
    nor g917(n1762 ,n641 ,n539);
    nor g918(n1761 ,n615 ,n1295);
    nor g919(n1760 ,n666 ,n1295);
    nor g920(n1759 ,n631 ,n539);
    nor g921(n1758 ,n630 ,n1295);
    nor g922(n1757 ,n681 ,n1295);
    nor g923(n1756 ,n668 ,n1295);
    nor g924(n1755 ,n671 ,n539);
    nor g925(n1754 ,n590 ,n539);
    nor g926(n1753 ,n684 ,n1295);
    nor g927(n1752 ,n617 ,n539);
    nor g928(n1751 ,n587 ,n539);
    nor g929(n1750 ,n645 ,n1295);
    nor g930(n1749 ,n680 ,n1295);
    nor g931(n1748 ,n683 ,n1295);
    nor g932(n1747 ,n626 ,n1295);
    nor g933(n1746 ,n672 ,n1295);
    nor g934(n1745 ,n583 ,n539);
    nor g935(n1744 ,n596 ,n1295);
    nor g936(n1743 ,n648 ,n539);
    nor g937(n1742 ,n640 ,n539);
    nor g938(n1741 ,n690 ,n539);
    nor g939(n1740 ,n673 ,n539);
    nor g940(n1739 ,n625 ,n539);
    nor g941(n1738 ,n678 ,n1295);
    nor g942(n1737 ,n675 ,n1295);
    nor g943(n1736 ,n566 ,n1295);
    nor g944(n1735 ,n692 ,n539);
    nor g945(n1734 ,n567 ,n539);
    nor g946(n1733 ,n674 ,n539);
    nor g947(n1732 ,n568 ,n1295);
    nor g948(n1731 ,n650 ,n1295);
    nor g949(n1730 ,n579 ,n539);
    nor g950(n1729 ,n609 ,n539);
    nor g951(n1728 ,n600 ,n1295);
    nor g952(n1727 ,n594 ,n539);
    nor g953(n1726 ,n571 ,n1295);
    nor g954(n1725 ,n679 ,n1295);
    nor g955(n1724 ,n638 ,n539);
    nor g956(n1723 ,n577 ,n539);
    nor g957(n1722 ,n620 ,n539);
    nor g958(n1721 ,n621 ,n539);
    nor g959(n1720 ,n598 ,n539);
    nor g960(n1719 ,n669 ,n1295);
    nor g961(n1718 ,n607 ,n1295);
    nor g962(n1717 ,n601 ,n539);
    nor g963(n1716 ,n614 ,n1295);
    nor g964(n1715 ,n605 ,n539);
    nor g965(n1714 ,n649 ,n1295);
    nor g966(n1713 ,n688 ,n539);
    nor g967(n1712 ,n685 ,n1295);
    nor g968(n1711 ,n656 ,n1295);
    nor g969(n1710 ,n623 ,n539);
    nor g970(n1709 ,n644 ,n539);
    nor g971(n1708 ,n667 ,n1295);
    nor g972(n1707 ,n686 ,n1295);
    nor g973(n1706 ,n661 ,n1295);
    nor g974(n1705 ,n660 ,n1295);
    nor g975(n1704 ,n642 ,n1295);
    nor g976(n1703 ,n646 ,n1295);
    nor g977(n1702 ,n565 ,n539);
    nor g978(n1701 ,n664 ,n539);
    nor g979(n1700 ,n632 ,n539);
    nor g980(n1699 ,n675 ,n538);
    nor g981(n1698 ,n678 ,n538);
    nor g982(n1697 ,n566 ,n538);
    nor g983(n1696 ,n692 ,n535);
    nor g984(n1695 ,n567 ,n535);
    nor g985(n1694 ,n674 ,n538);
    nor g986(n1693 ,n568 ,n538);
    nor g987(n1692 ,n650 ,n538);
    nor g988(n1691 ,n579 ,n535);
    nor g989(n1690 ,n609 ,n538);
    nor g990(n1689 ,n600 ,n538);
    nor g991(n1688 ,n772 ,n536);
    nor g992(n1687 ,n594 ,n535);
    nor g993(n1686 ,n571 ,n538);
    nor g994(n1685 ,n679 ,n535);
    nor g995(n1684 ,n638 ,n535);
    nor g996(n1683 ,n577 ,n535);
    nor g997(n1682 ,n620 ,n536);
    nor g998(n1681 ,n621 ,n535);
    nor g999(n1680 ,n598 ,n536);
    nor g1000(n1679 ,n669 ,n536);
    nor g1001(n1678 ,n607 ,n535);
    nor g1002(n1677 ,n601 ,n535);
    nor g1003(n1676 ,n614 ,n538);
    nor g1004(n1675 ,n605 ,n536);
    nor g1005(n1674 ,n796 ,n538);
    nor g1006(n1673 ,n649 ,n538);
    nor g1007(n1672 ,n688 ,n536);
    nor g1008(n1671 ,n685 ,n536);
    nor g1009(n1670 ,n656 ,n535);
    nor g1010(n1669 ,n623 ,n535);
    nor g1011(n1668 ,n644 ,n535);
    nor g1012(n1667 ,n786 ,n535);
    nor g1013(n1666 ,n667 ,n538);
    nor g1014(n1665 ,n686 ,n535);
    nor g1015(n1664 ,n581 ,n536);
    nor g1016(n1663 ,n661 ,n538);
    nor g1017(n1662 ,n660 ,n535);
    nor g1018(n1661 ,n642 ,n536);
    nor g1019(n1660 ,n646 ,n536);
    nor g1020(n1659 ,n565 ,n536);
    nor g1021(n1658 ,n664 ,n535);
    nor g1022(n1657 ,n632 ,n535);
    nor g1023(n1656 ,n757 ,n538);
    nor g1024(n1655 ,n776 ,n536);
    nor g1025(n1654 ,n789 ,n536);
    nor g1026(n1653 ,n732 ,n535);
    nor g1027(n1652 ,n814 ,n538);
    nor g1028(n1651 ,n769 ,n535);
    nor g1029(n1650 ,n755 ,n535);
    nor g1030(n1649 ,n695 ,n536);
    nor g1031(n1648 ,n698 ,n536);
    nor g1032(n1647 ,n718 ,n536);
    nor g1033(n1646 ,n749 ,n538);
    nor g1034(n1645 ,n735 ,n535);
    nor g1035(n1644 ,n693 ,n536);
    nor g1036(n1643 ,n779 ,n535);
    nor g1037(n1642 ,n697 ,n535);
    nor g1038(n1641 ,n799 ,n538);
    nor g1039(n1640 ,n700 ,n535);
    nor g1040(n1639 ,n791 ,n538);
    nor g1041(n1638 ,n725 ,n535);
    nor g1042(n1637 ,n743 ,n538);
    nor g1043(n1636 ,n777 ,n538);
    nor g1044(n1635 ,n794 ,n538);
    nor g1045(n1634 ,n803 ,n538);
    nor g1046(n1633 ,n738 ,n535);
    nor g1047(n1632 ,n767 ,n538);
    nor g1048(n1631 ,n788 ,n535);
    nor g1049(n1630 ,n809 ,n538);
    nor g1050(n1629 ,n797 ,n538);
    nor g1051(n1628 ,n883 ,n541);
    not g1052(n1622 ,n1623);
    or g1053(n1621 ,n1243 ,n1349);
    nor g1054(n1620 ,n739 ,n538);
    nor g1055(n1619 ,n775 ,n535);
    nor g1056(n1618 ,n750 ,n535);
    nor g1057(n1617 ,n726 ,n538);
    nor g1058(n1616 ,n806 ,n538);
    nor g1059(n1615 ,n704 ,n536);
    nor g1060(n1614 ,n751 ,n536);
    nor g1061(n1613 ,n746 ,n536);
    nor g1062(n1612 ,n696 ,n538);
    nor g1063(n1611 ,n707 ,n535);
    nor g1064(n1610 ,n810 ,n538);
    nor g1065(n1609 ,n761 ,n538);
    nor g1066(n1608 ,n787 ,n538);
    nor g1067(n1607 ,n694 ,n535);
    nor g1068(n1606 ,n699 ,n538);
    nor g1069(n1605 ,n719 ,n536);
    nor g1070(n1604 ,n805 ,n536);
    nor g1071(n1603 ,n641 ,n535);
    nor g1072(n1602 ,n752 ,n538);
    nor g1073(n1601 ,n705 ,n535);
    nor g1074(n1600 ,n747 ,n536);
    nor g1075(n1599 ,n784 ,n535);
    nor g1076(n1598 ,n714 ,n536);
    nor g1077(n1597 ,n728 ,n538);
    nor g1078(n1596 ,n615 ,n535);
    nor g1079(n1595 ,n763 ,n535);
    nor g1080(n1594 ,n742 ,n538);
    nor g1081(n1593 ,n808 ,n538);
    nor g1082(n1592 ,n733 ,n538);
    nor g1083(n1591 ,n666 ,n535);
    nor g1084(n1590 ,n711 ,n536);
    nor g1085(n1589 ,n731 ,n536);
    nor g1086(n1588 ,n745 ,n538);
    nor g1087(n1587 ,n795 ,n538);
    nor g1088(n1586 ,n631 ,n535);
    nor g1089(n1585 ,n630 ,n535);
    nor g1090(n1584 ,n681 ,n535);
    nor g1091(n1583 ,n668 ,n538);
    nor g1092(n1582 ,n671 ,n535);
    nor g1093(n1581 ,n590 ,n538);
    nor g1094(n1580 ,n684 ,n535);
    nor g1095(n1579 ,n617 ,n535);
    nor g1096(n1578 ,n587 ,n538);
    nor g1097(n1577 ,n645 ,n536);
    nor g1098(n1576 ,n680 ,n536);
    nor g1099(n1575 ,n683 ,n535);
    nor g1100(n1574 ,n626 ,n538);
    nor g1101(n1573 ,n672 ,n536);
    nor g1102(n1572 ,n583 ,n538);
    nor g1103(n1571 ,n596 ,n535);
    nor g1104(n1570 ,n648 ,n536);
    nor g1105(n1569 ,n640 ,n535);
    nor g1106(n1568 ,n690 ,n538);
    nor g1107(n1567 ,n673 ,n535);
    nor g1108(n1566 ,n625 ,n536);
    or g1109(n1565 ,n1186 ,n1246);
    nor g1110(n1564 ,n1122 ,n1182);
    nor g1111(n1563 ,n1121 ,n1173);
    nor g1112(n1562 ,n1119 ,n1179);
    nor g1113(n1561 ,n1118 ,n1172);
    nor g1114(n1560 ,n1120 ,n1181);
    nor g1115(n1559 ,n1124 ,n1171);
    nor g1116(n1558 ,n1116 ,n1178);
    nor g1117(n1557 ,n1115 ,n1169);
    nor g1118(n1556 ,n1125 ,n1180);
    nor g1119(n1555 ,n1126 ,n1174);
    nor g1120(n1554 ,n1112 ,n1177);
    or g1121(n1553 ,n1253 ,n1391);
    nor g1122(n1552 ,n1113 ,n1170);
    nor g1123(n1551 ,n1123 ,n1176);
    nor g1124(n1550 ,n1111 ,n1168);
    nor g1125(n1549 ,n1114 ,n1175);
    nor g1126(n1548 ,n1117 ,n1167);
    or g1127(n1547 ,n1245 ,n1369);
    or g1128(n1546 ,n1244 ,n1368);
    or g1129(n1545 ,n1242 ,n1367);
    or g1130(n1544 ,n1241 ,n1366);
    or g1131(n1543 ,n1240 ,n1365);
    or g1132(n1542 ,n1239 ,n1364);
    or g1133(n1541 ,n1238 ,n1363);
    or g1134(n1540 ,n1359 ,n1397);
    or g1135(n1539 ,n1237 ,n1362);
    or g1136(n1538 ,n1236 ,n1361);
    or g1137(n1537 ,n1235 ,n1360);
    or g1138(n1536 ,n1215 ,n1358);
    or g1139(n1535 ,n1234 ,n1356);
    or g1140(n1534 ,n1233 ,n1355);
    or g1141(n1533 ,n1317 ,n1426);
    or g1142(n1532 ,n1232 ,n1354);
    or g1143(n1531 ,n1187 ,n1248);
    or g1144(n1530 ,n1188 ,n1249);
    or g1145(n1529 ,n1231 ,n1353);
    or g1146(n1528 ,n1230 ,n1352);
    or g1147(n1527 ,n1229 ,n1351);
    or g1148(n1526 ,n1290 ,n1398);
    or g1149(n1525 ,n1228 ,n1350);
    or g1150(n1524 ,n1357 ,n1429);
    nor g1151(n1523 ,n703 ,n538);
    or g1152(n1522 ,n1227 ,n1348);
    or g1153(n1521 ,n1284 ,n1392);
    or g1154(n1520 ,n1226 ,n1347);
    or g1155(n1519 ,n1225 ,n1346);
    or g1156(n1518 ,n1224 ,n1345);
    or g1157(n1517 ,n1223 ,n1344);
    or g1158(n1516 ,n1222 ,n1342);
    or g1159(n1515 ,n1221 ,n1341);
    or g1160(n1514 ,n1343 ,n1399);
    or g1161(n1513 ,n1206 ,n1340);
    or g1162(n1512 ,n1220 ,n1338);
    or g1163(n1511 ,n1219 ,n1337);
    or g1164(n1510 ,n1218 ,n1336);
    or g1165(n1509 ,n1217 ,n1335);
    or g1166(n1508 ,n1333 ,n1400);
    or g1167(n1507 ,n1208 ,n1334);
    or g1168(n1506 ,n1306 ,n1417);
    or g1169(n1505 ,n1216 ,n1332);
    or g1170(n1504 ,n1214 ,n1331);
    or g1171(n1503 ,n1326 ,n1427);
    or g1172(n1502 ,n1209 ,n1328);
    or g1173(n1501 ,n1212 ,n1327);
    or g1174(n1500 ,n1213 ,n1325);
    or g1175(n1499 ,n1211 ,n1324);
    or g1176(n1498 ,n1329 ,n1428);
    or g1177(n1497 ,n1207 ,n1323);
    or g1178(n1496 ,n1210 ,n1322);
    or g1179(n1495 ,n1299 ,n1405);
    or g1180(n1494 ,n1320 ,n1373);
    or g1181(n1493 ,n1287 ,n1383);
    or g1182(n1492 ,n1339 ,n1401);
    or g1183(n1491 ,n1189 ,n1251);
    or g1184(n1490 ,n1316 ,n1374);
    or g1185(n1489 ,n1318 ,n1393);
    or g1186(n1488 ,n1312 ,n1420);
    or g1187(n1487 ,n1311 ,n1425);
    or g1188(n1486 ,n1289 ,n1424);
    or g1189(n1485 ,n1310 ,n1423);
    or g1190(n1484 ,n1301 ,n1422);
    or g1191(n1483 ,n1315 ,n1419);
    or g1192(n1482 ,n1319 ,n1418);
    or g1193(n1481 ,n1308 ,n1421);
    or g1194(n1480 ,n1302 ,n1379);
    or g1195(n1479 ,n1305 ,n1416);
    or g1196(n1478 ,n1275 ,n1378);
    or g1197(n1477 ,n1250 ,n1415);
    or g1198(n1476 ,n1273 ,n1412);
    or g1199(n1475 ,n1278 ,n1411);
    or g1200(n1474 ,n1285 ,n1407);
    or g1201(n1473 ,n1291 ,n1406);
    or g1202(n1472 ,n1277 ,n1409);
    or g1203(n1471 ,n1247 ,n1404);
    or g1204(n1470 ,n1309 ,n1403);
    or g1205(n1469 ,n1288 ,n1402);
    or g1206(n1468 ,n1292 ,n1381);
    or g1207(n1467 ,n1321 ,n1396);
    or g1208(n1466 ,n1293 ,n1395);
    or g1209(n1465 ,n1283 ,n1408);
    or g1210(n1464 ,n1269 ,n1389);
    or g1211(n1463 ,n1280 ,n1370);
    or g1212(n1462 ,n1276 ,n1387);
    or g1213(n1461 ,n1281 ,n1386);
    or g1214(n1460 ,n1298 ,n1385);
    or g1215(n1459 ,n1300 ,n1410);
    or g1216(n1458 ,n1313 ,n1384);
    or g1217(n1457 ,n1279 ,n1382);
    or g1218(n1456 ,n1314 ,n1394);
    or g1219(n1455 ,n1304 ,n1380);
    or g1220(n1454 ,n1307 ,n1377);
    or g1221(n1453 ,n1274 ,n1376);
    or g1222(n1452 ,n1282 ,n1388);
    or g1223(n1451 ,n1286 ,n1375);
    or g1224(n1450 ,n1272 ,n1372);
    or g1225(n1449 ,n1330 ,n1371);
    or g1226(n1448 ,n1205 ,n1271);
    or g1227(n1447 ,n1204 ,n1268);
    or g1228(n1446 ,n1203 ,n1267);
    or g1229(n1445 ,n1202 ,n1265);
    or g1230(n1444 ,n1270 ,n1413);
    or g1231(n1443 ,n1201 ,n1264);
    or g1232(n1442 ,n1200 ,n1263);
    or g1233(n1441 ,n1199 ,n1262);
    or g1234(n1440 ,n1198 ,n1261);
    or g1235(n1439 ,n1197 ,n1260);
    or g1236(n1438 ,n1196 ,n1259);
    or g1237(n1437 ,n1195 ,n1258);
    or g1238(n1436 ,n1303 ,n1414);
    or g1239(n1435 ,n1194 ,n1257);
    or g1240(n1434 ,n1193 ,n1256);
    or g1241(n1433 ,n1192 ,n1255);
    or g1242(n1432 ,n1266 ,n1390);
    or g1243(n1431 ,n1191 ,n1254);
    or g1244(n1430 ,n1190 ,n1252);
    nor g1245(n1627 ,n1133 ,n1184);
    or g1246(n1626 ,n548 ,n1166);
    or g1247(n1625 ,n548 ,n1297);
    or g1248(n1624 ,n1144 ,n1185);
    nor g1249(n1623 ,n1297 ,n1183);
    nor g1250(n1429 ,n864 ,n532);
    nor g1251(n1428 ,n956 ,n533);
    nor g1252(n1427 ,n945 ,n532);
    nor g1253(n1426 ,n973 ,n533);
    nor g1254(n1425 ,n940 ,n533);
    nor g1255(n1424 ,n831 ,n533);
    nor g1256(n1423 ,n835 ,n532);
    nor g1257(n1422 ,n838 ,n532);
    nor g1258(n1421 ,n842 ,n533);
    nor g1259(n1420 ,n846 ,n533);
    nor g1260(n1419 ,n849 ,n532);
    nor g1261(n1418 ,n852 ,n533);
    nor g1262(n1417 ,n856 ,n532);
    nor g1263(n1416 ,n915 ,n532);
    nor g1264(n1415 ,n929 ,n533);
    nor g1265(n1414 ,n913 ,n532);
    nor g1266(n1413 ,n997 ,n532);
    nor g1267(n1412 ,n859 ,n533);
    nor g1268(n1411 ,n884 ,n533);
    nor g1269(n1410 ,n879 ,n532);
    nor g1270(n1409 ,n1009 ,n533);
    nor g1271(n1408 ,n908 ,n532);
    nor g1272(n1407 ,n953 ,n532);
    nor g1273(n1406 ,n834 ,n532);
    nor g1274(n1405 ,n876 ,n532);
    nor g1275(n1404 ,n987 ,n533);
    nor g1276(n1403 ,n857 ,n533);
    nor g1277(n1402 ,n901 ,n532);
    nor g1278(n1401 ,n832 ,n533);
    nor g1279(n1400 ,n976 ,n533);
    nor g1280(n1399 ,n870 ,n533);
    nor g1281(n1398 ,n872 ,n533);
    nor g1282(n1397 ,n880 ,n532);
    nor g1283(n1396 ,n1013 ,n533);
    nor g1284(n1395 ,n970 ,n532);
    nor g1285(n1394 ,n999 ,n532);
    nor g1286(n1393 ,n1003 ,n532);
    nor g1287(n1392 ,n885 ,n532);
    nor g1288(n1391 ,n971 ,n532);
    nor g1289(n1390 ,n955 ,n532);
    nor g1290(n1389 ,n906 ,n533);
    nor g1291(n1388 ,n967 ,n533);
    nor g1292(n1387 ,n941 ,n533);
    nor g1293(n1386 ,n935 ,n532);
    nor g1294(n1385 ,n853 ,n533);
    nor g1295(n1384 ,n986 ,n533);
    nor g1296(n1383 ,n992 ,n532);
    nor g1297(n1382 ,n936 ,n532);
    nor g1298(n1381 ,n998 ,n532);
    nor g1299(n1380 ,n891 ,n532);
    nor g1300(n1379 ,n847 ,n533);
    nor g1301(n1378 ,n961 ,n532);
    nor g1302(n1377 ,n942 ,n533);
    nor g1303(n1376 ,n931 ,n533);
    nor g1304(n1375 ,n1006 ,n532);
    nor g1305(n1374 ,n991 ,n533);
    nor g1306(n1373 ,n964 ,n532);
    nor g1307(n1372 ,n917 ,n532);
    nor g1308(n1371 ,n837 ,n532);
    nor g1309(n1370 ,n962 ,n533);
    nor g1310(n1369 ,n778 ,n534);
    nor g1311(n1368 ,n804 ,n1159);
    nor g1312(n1367 ,n702 ,n534);
    nor g1313(n1366 ,n774 ,n534);
    nor g1314(n1365 ,n628 ,n534);
    nor g1315(n1364 ,n662 ,n534);
    nor g1316(n1363 ,n603 ,n1159);
    nor g1317(n1362 ,n602 ,n534);
    nor g1318(n1361 ,n658 ,n534);
    nor g1319(n1360 ,n592 ,n534);
    nor g1320(n1359 ,n790 ,n529);
    nor g1321(n1358 ,n657 ,n1159);
    nor g1322(n1357 ,n760 ,n1155);
    nor g1323(n1356 ,n595 ,n534);
    nor g1324(n1355 ,n569 ,n534);
    nor g1325(n1354 ,n573 ,n1159);
    nor g1326(n1353 ,n636 ,n534);
    nor g1327(n1352 ,n653 ,n1159);
    nor g1328(n1351 ,n585 ,n1159);
    nor g1329(n1350 ,n564 ,n1159);
    nor g1330(n1349 ,n639 ,n1159);
    nor g1331(n1348 ,n588 ,n1159);
    nor g1332(n1347 ,n643 ,n1159);
    nor g1333(n1346 ,n619 ,n1159);
    nor g1334(n1345 ,n652 ,n534);
    nor g1335(n1344 ,n591 ,n534);
    nor g1336(n1343 ,n608 ,n529);
    nor g1337(n1342 ,n582 ,n534);
    nor g1338(n1341 ,n634 ,n1159);
    nor g1339(n1340 ,n663 ,n1159);
    nor g1340(n1339 ,n599 ,n529);
    nor g1341(n1338 ,n574 ,n1159);
    nor g1342(n1337 ,n570 ,n534);
    nor g1343(n1336 ,n593 ,n534);
    nor g1344(n1335 ,n659 ,n1159);
    nor g1345(n1334 ,n562 ,n1159);
    nor g1346(n1333 ,n647 ,n529);
    nor g1347(n1332 ,n589 ,n534);
    nor g1348(n1331 ,n610 ,n1159);
    nor g1349(n1330 ,n759 ,n529);
    nor g1350(n1329 ,n622 ,n1155);
    nor g1351(n1328 ,n670 ,n1159);
    nor g1352(n1327 ,n689 ,n1159);
    nor g1353(n1326 ,n616 ,n529);
    nor g1354(n1325 ,n665 ,n1159);
    nor g1355(n1324 ,n612 ,n1159);
    nor g1356(n1323 ,n576 ,n1159);
    nor g1357(n1322 ,n627 ,n534);
    nor g1358(n1321 ,n807 ,n529);
    nor g1359(n1320 ,n765 ,n529);
    nor g1360(n1319 ,n572 ,n1155);
    nor g1361(n1318 ,n712 ,n529);
    nor g1362(n1317 ,n783 ,n529);
    nor g1363(n1316 ,n713 ,n1155);
    nor g1364(n1315 ,n687 ,n529);
    nor g1365(n1314 ,n800 ,n1155);
    nor g1366(n1313 ,n734 ,n1155);
    nor g1367(n1312 ,n654 ,n1155);
    nor g1368(n1311 ,n676 ,n1155);
    nor g1369(n1310 ,n655 ,n1155);
    nor g1370(n1309 ,n637 ,n1155);
    nor g1371(n1308 ,n575 ,n1155);
    nor g1372(n1307 ,n710 ,n529);
    nor g1373(n1306 ,n618 ,n529);
    nor g1374(n1305 ,n651 ,n529);
    nor g1375(n1304 ,n812 ,n1155);
    nor g1376(n1303 ,n606 ,n1155);
    nor g1377(n1302 ,n748 ,n1155);
    nor g1378(n1301 ,n635 ,n529);
    nor g1379(n1300 ,n580 ,n529);
    nor g1380(n1299 ,n677 ,n1155);
    nor g1381(n1298 ,n744 ,n1155);
    not g1382(n540 ,n1296);
    not g1383(n541 ,n1296);
    not g1384(n1295 ,n1294);
    not g1385(n539 ,n1294);
    not g1386(n535 ,n537);
    not g1387(n536 ,n537);
    not g1388(n537 ,n538);
    nor g1389(n1293 ,n730 ,n529);
    nor g1390(n1292 ,n741 ,n1155);
    nor g1391(n1291 ,n633 ,n1155);
    nor g1392(n1290 ,n811 ,n1155);
    nor g1393(n1289 ,n604 ,n1155);
    nor g1394(n1288 ,n613 ,n1155);
    nor g1395(n1287 ,n715 ,n1155);
    nor g1396(n1286 ,n782 ,n529);
    nor g1397(n1285 ,n611 ,n529);
    nor g1398(n1284 ,n813 ,n529);
    nor g1399(n1283 ,n561 ,n529);
    nor g1400(n1282 ,n780 ,n529);
    nor g1401(n1281 ,n766 ,n1155);
    nor g1402(n1280 ,n723 ,n1155);
    nor g1403(n1279 ,n724 ,n1155);
    nor g1404(n1278 ,n691 ,n529);
    nor g1405(n1277 ,n722 ,n529);
    nor g1406(n1276 ,n758 ,n1155);
    nor g1407(n1275 ,n768 ,n1155);
    nor g1408(n1274 ,n717 ,n1155);
    nor g1409(n1273 ,n624 ,n529);
    nor g1410(n1272 ,n708 ,n529);
    nor g1411(n1271 ,n771 ,n534);
    nor g1412(n1270 ,n586 ,n1155);
    nor g1413(n1269 ,n764 ,n529);
    nor g1414(n1268 ,n720 ,n534);
    nor g1415(n1267 ,n773 ,n534);
    nor g1416(n1266 ,n792 ,n1155);
    nor g1417(n1265 ,n716 ,n534);
    nor g1418(n1264 ,n762 ,n1159);
    nor g1419(n1263 ,n740 ,n1159);
    nor g1420(n1262 ,n781 ,n1159);
    nor g1421(n1261 ,n793 ,n534);
    nor g1422(n1260 ,n729 ,n534);
    nor g1423(n1259 ,n801 ,n1159);
    nor g1424(n1258 ,n815 ,n1159);
    nor g1425(n1257 ,n721 ,n1159);
    nor g1426(n1256 ,n756 ,n534);
    nor g1427(n1255 ,n785 ,n534);
    nor g1428(n1254 ,n754 ,n1159);
    nor g1429(n1253 ,n753 ,n1155);
    nor g1430(n1252 ,n701 ,n534);
    nor g1431(n1251 ,n727 ,n1159);
    nor g1432(n1250 ,n578 ,n529);
    nor g1433(n1249 ,n770 ,n1159);
    nor g1434(n1248 ,n709 ,n534);
    nor g1435(n1247 ,n563 ,n1155);
    nor g1436(n1246 ,n736 ,n1159);
    nor g1437(n1245 ,n993 ,n530);
    nor g1438(n1244 ,n1002 ,n531);
    nor g1439(n1243 ,n900 ,n530);
    nor g1440(n1242 ,n925 ,n531);
    nor g1441(n1241 ,n977 ,n531);
    nor g1442(n1240 ,n890 ,n531);
    nor g1443(n1239 ,n938 ,n530);
    nor g1444(n1238 ,n905 ,n530);
    nor g1445(n1237 ,n921 ,n531);
    nor g1446(n1236 ,n981 ,n531);
    nor g1447(n1235 ,n944 ,n530);
    nor g1448(n1234 ,n854 ,n531);
    nor g1449(n1233 ,n975 ,n530);
    nor g1450(n1232 ,n933 ,n530);
    nor g1451(n1231 ,n877 ,n531);
    nor g1452(n1230 ,n898 ,n530);
    nor g1453(n1229 ,n952 ,n530);
    nor g1454(n1228 ,n839 ,n531);
    nor g1455(n1227 ,n907 ,n531);
    nor g1456(n1226 ,n893 ,n530);
    nor g1457(n1225 ,n984 ,n531);
    nor g1458(n1224 ,n937 ,n530);
    nor g1459(n1223 ,n904 ,n530);
    nor g1460(n1222 ,n927 ,n530);
    nor g1461(n1221 ,n843 ,n530);
    nor g1462(n1220 ,n886 ,n531);
    nor g1463(n1219 ,n912 ,n531);
    nor g1464(n1218 ,n954 ,n530);
    nor g1465(n1217 ,n983 ,n531);
    nor g1466(n1216 ,n868 ,n531);
    nor g1467(n1215 ,n841 ,n531);
    nor g1468(n1214 ,n980 ,n531);
    nor g1469(n1213 ,n896 ,n530);
    nor g1470(n1212 ,n892 ,n531);
    nor g1471(n1211 ,n920 ,n530);
    nor g1472(n1210 ,n873 ,n530);
    nor g1473(n1209 ,n865 ,n530);
    nor g1474(n1208 ,n1001 ,n530);
    nor g1475(n1207 ,n874 ,n530);
    nor g1476(n1206 ,n932 ,n530);
    nor g1477(n1205 ,n869 ,n531);
    nor g1478(n1204 ,n848 ,n531);
    nor g1479(n1203 ,n1010 ,n531);
    nor g1480(n1202 ,n982 ,n530);
    nor g1481(n1201 ,n969 ,n531);
    nor g1482(n1200 ,n902 ,n531);
    nor g1483(n1199 ,n943 ,n530);
    nor g1484(n1198 ,n909 ,n530);
    nor g1485(n1197 ,n858 ,n530);
    nor g1486(n1196 ,n840 ,n530);
    nor g1487(n1195 ,n928 ,n531);
    nor g1488(n1194 ,n1005 ,n530);
    nor g1489(n1193 ,n881 ,n531);
    nor g1490(n1192 ,n860 ,n531);
    nor g1491(n1191 ,n934 ,n530);
    nor g1492(n1190 ,n985 ,n531);
    nor g1493(n1189 ,n958 ,n530);
    nor g1494(n1188 ,n960 ,n530);
    nor g1495(n1187 ,n897 ,n530);
    nor g1496(n1186 ,n957 ,n531);
    or g1497(n1185 ,n548 ,n1163);
    nor g1498(n1184 ,n547 ,n1152);
    or g1499(n1183 ,n1161 ,n1150);
    or g1500(n1182 ,n1027 ,n1160);
    or g1501(n1181 ,n1017 ,n1160);
    or g1502(n1180 ,n1028 ,n1160);
    or g1503(n1179 ,n1021 ,n1160);
    or g1504(n1178 ,n1029 ,n1160);
    or g1505(n1177 ,n1019 ,n1160);
    or g1506(n1176 ,n1030 ,n1160);
    or g1507(n1175 ,n1031 ,n1160);
    or g1508(n1174 ,n1018 ,n529);
    or g1509(n1173 ,n1020 ,n529);
    or g1510(n1172 ,n1024 ,n529);
    or g1511(n1171 ,n1026 ,n529);
    or g1512(n1170 ,n1023 ,n534);
    or g1513(n1169 ,n1022 ,n534);
    or g1514(n1168 ,n1035 ,n534);
    or g1515(n1167 ,n1034 ,n534);
    nor g1516(n1166 ,n1163 ,n1164);
    nor g1517(n1297 ,n1142 ,n1153);
    nor g1518(n1296 ,n551 ,n1161);
    nor g1519(n1294 ,n552 ,n1162);
    or g1520(n538 ,n548 ,n1165);
    not g1521(n1165 ,n1164);
    not g1522(n1162 ,n1161);
    not g1523(n1159 ,n1158);
    not g1524(n534 ,n1158);
    nor g1525(n1164 ,n7[0] ,n1149);
    nor g1526(n1163 ,n816 ,n1147);
    nor g1527(n1161 ,n7[0] ,n1147);
    or g1528(n1160 ,n1073 ,n1147);
    nor g1529(n1158 ,n551 ,n1151);
    not g1530(n532 ,n1157);
    not g1531(n533 ,n1157);
    not g1532(n530 ,n1156);
    not g1533(n531 ,n1156);
    not g1534(n1155 ,n1154);
    not g1535(n529 ,n1154);
    nor g1536(n1153 ,n7[0] ,n1148);
    or g1537(n1152 ,n1148 ,n1146);
    nor g1538(n1157 ,n542 ,n1143);
    or g1539(n1156 ,n1072 ,n1141);
    nor g1540(n1154 ,n2068 ,n1145);
    not g1541(n1151 ,n1150);
    not g1542(n1149 ,n1148);
    not g1543(n1147 ,n1146);
    or g1544(n1145 ,n1073 ,n1140);
    nor g1545(n1150 ,n1015 ,n1140);
    nor g1546(n1148 ,n817 ,n1138);
    nor g1547(n1146 ,n528 ,n1140);
    nor g1548(n1144 ,n7[0] ,n1138);
    nor g1549(n1143 ,n1135 ,n1138);
    nor g1550(n1142 ,n816 ,n1139);
    nor g1551(n1141 ,n550 ,n1137);
    not g1552(n1140 ,n1139);
    nor g1553(n1139 ,n2069 ,n1136);
    not g1554(n1138 ,n1137);
    nor g1555(n1137 ,n2068 ,n1136);
    xnor g1556(n1135 ,n817 ,n816);
    xnor g1557(n1134 ,n7[0] ,n2068);
    nor g1558(n1133 ,n817 ,n1073);
    or g1559(n1136 ,n1132 ,n1131);
    or g1560(n1132 ,n830 ,n895);
    or g1561(n1131 ,n861 ,n871);
    nor g1562(n1130 ,n825 ,n556);
    nor g1563(n1129 ,n822 ,n554);
    nor g1564(n1128 ,n824 ,n555);
    nor g1565(n1127 ,n821 ,n553);
    nor g1566(n1126 ,n559 ,n553);
    nor g1567(n1125 ,n826 ,n553);
    nor g1568(n1124 ,n558 ,n555);
    nor g1569(n1123 ,n829 ,n555);
    nor g1570(n1122 ,n819 ,n554);
    nor g1571(n1121 ,n557 ,n554);
    nor g1572(n1120 ,n823 ,n555);
    nor g1573(n1119 ,n820 ,n556);
    nor g1574(n1118 ,n560 ,n556);
    nor g1575(n1117 ,n597 ,n553);
    nor g1576(n1116 ,n827 ,n556);
    nor g1577(n1115 ,n584 ,n556);
    nor g1578(n1114 ,n818 ,n553);
    nor g1579(n1113 ,n682 ,n554);
    nor g1580(n1112 ,n828 ,n554);
    nor g1581(n1111 ,n629 ,n555);
    nor g1582(n1110 ,n643 ,n542);
    nor g1583(n1109 ,n591 ,n551);
    nor g1584(n1108 ,n575 ,n552);
    nor g1585(n1107 ,n619 ,n546);
    nor g1586(n1106 ,n593 ,n551);
    nor g1587(n1105 ,n676 ,n551);
    nor g1588(n1104 ,n588 ,n550);
    nor g1589(n1103 ,n564 ,n542);
    nor g1590(n1102 ,n653 ,n551);
    nor g1591(n1101 ,n610 ,n547);
    nor g1592(n1100 ,n627 ,n544);
    nor g1593(n1099 ,n602 ,n544);
    nor g1594(n1098 ,n576 ,n549);
    nor g1595(n1097 ,n589 ,n546);
    nor g1596(n1096 ,n569 ,n547);
    nor g1597(n1095 ,n595 ,n543);
    nor g1598(n1094 ,n658 ,n547);
    nor g1599(n1093 ,n689 ,n545);
    nor g1600(n1092 ,n573 ,n547);
    nor g1601(n1091 ,n662 ,n542);
    nor g1602(n1090 ,n628 ,n543);
    nor g1603(n1089 ,n659 ,n543);
    nor g1604(n1088 ,n557 ,n545);
    nor g1605(n1087 ,n560 ,n545);
    nor g1606(n1086 ,n558 ,n543);
    nor g1607(n1085 ,n559 ,n548);
    nor g1608(n1084 ,n604 ,n543);
    nor g1609(n1083 ,n655 ,n542);
    nor g1610(n1082 ,n635 ,n545);
    nor g1611(n1081 ,n654 ,n547);
    nor g1612(n1080 ,n687 ,n546);
    nor g1613(n1079 ,n572 ,n549);
    nor g1614(n1078 ,n622 ,n544);
    nor g1615(n1077 ,n651 ,n544);
    nor g1616(n1076 ,n578 ,n544);
    nor g1617(n1075 ,n586 ,n544);
    nor g1618(n1074 ,n624 ,n550);
    not g1619(n1073 ,n1072);
    nor g1620(n1071 ,n691 ,n546);
    nor g1621(n1070 ,n561 ,n546);
    nor g1622(n1069 ,n611 ,n551);
    nor g1623(n1068 ,n633 ,n551);
    nor g1624(n1067 ,n563 ,n552);
    nor g1625(n1066 ,n637 ,n542);
    nor g1626(n1065 ,n613 ,n542);
    nor g1627(n1064 ,n616 ,n548);
    nor g1628(n1063 ,n608 ,n549);
    nor g1629(n1062 ,n582 ,n545);
    nor g1630(n1061 ,n634 ,n546);
    nor g1631(n1060 ,n670 ,n543);
    nor g1632(n1059 ,n652 ,n548);
    nor g1633(n1058 ,n647 ,n547);
    nor g1634(n1057 ,n592 ,n543);
    nor g1635(n1056 ,n612 ,n544);
    nor g1636(n1055 ,n639 ,n544);
    nor g1637(n1054 ,n562 ,n550);
    nor g1638(n1053 ,n585 ,n546);
    nor g1639(n1052 ,n599 ,n542);
    nor g1640(n1051 ,n636 ,n550);
    nor g1641(n1050 ,n665 ,n548);
    nor g1642(n1049 ,n677 ,n549);
    nor g1643(n1048 ,n603 ,n546);
    nor g1644(n1047 ,n580 ,n545);
    nor g1645(n1046 ,n574 ,n547);
    nor g1646(n1045 ,n606 ,n549);
    nor g1647(n1044 ,n618 ,n552);
    nor g1648(n1043 ,n802 ,n552);
    nor g1649(n1042 ,n657 ,n545);
    nor g1650(n1041 ,n663 ,n545);
    nor g1651(n1040 ,n706 ,n549);
    nor g1652(n1039 ,n737 ,n552);
    nor g1653(n1038 ,n570 ,n543);
    nor g1654(n1037 ,n5[1] ,n6[1]);
    nor g1655(n1036 ,n8[0] ,n552);
    nor g1656(n1035 ,n2[2] ,n6[2]);
    nor g1657(n1034 ,n2[3] ,n6[3]);
    nor g1658(n1033 ,n5[0] ,n6[0]);
    nor g1659(n1032 ,n5[2] ,n6[2]);
    nor g1660(n1031 ,n3[3] ,n6[3]);
    nor g1661(n1030 ,n3[2] ,n6[2]);
    nor g1662(n1029 ,n3[1] ,n6[1]);
    nor g1663(n1028 ,n4[3] ,n6[3]);
    nor g1664(n1027 ,n4[0] ,n6[0]);
    nor g1665(n1026 ,n2[66] ,n6[2]);
    nor g1666(n1025 ,n5[3] ,n6[3]);
    nor g1667(n1024 ,n2[65] ,n6[1]);
    nor g1668(n1023 ,n2[0] ,n6[0]);
    nor g1669(n1022 ,n2[1] ,n6[1]);
    nor g1670(n1021 ,n4[1] ,n6[1]);
    nor g1671(n1020 ,n2[64] ,n6[0]);
    nor g1672(n1019 ,n3[0] ,n6[0]);
    nor g1673(n1018 ,n2[67] ,n6[3]);
    nor g1674(n1017 ,n4[2] ,n6[2]);
    or g1675(n1016 ,n7[0] ,n2069);
    or g1676(n1015 ,n7[0] ,n2068);
    or g1677(n1014 ,n816 ,n528);
    nor g1678(n1072 ,n816 ,n550);
    not g1679(n1013 ,n4[35]);
    not g1680(n1012 ,n5[9]);
    not g1681(n1011 ,n5[28]);
    not g1682(n1010 ,n3[6]);
    not g1683(n1009 ,n4[54]);
    not g1684(n1008 ,n5[44]);
    not g1685(n1007 ,n5[33]);
    not g1686(n1006 ,n4[59]);
    not g1687(n1005 ,n3[15]);
    not g1688(n1004 ,n5[54]);
    not g1689(n1003 ,n4[39]);
    not g1690(n1002 ,n3[25]);
    not g1691(n1001 ,n3[55]);
    not g1692(n1000 ,n5[29]);
    not g1693(n999 ,n4[38]);
    not g1694(n998 ,n4[52]);
    not g1695(n997 ,n4[17]);
    not g1696(n996 ,n5[19]);
    not g1697(n995 ,n5[59]);
    not g1698(n994 ,n5[25]);
    not g1699(n993 ,n3[24]);
    not g1700(n992 ,n4[50]);
    not g1701(n991 ,n4[60]);
    not g1702(n990 ,n5[36]);
    not g1703(n989 ,n5[56]);
    not g1704(n988 ,n5[35]);
    not g1705(n987 ,n4[25]);
    not g1706(n986 ,n4[49]);
    not g1707(n985 ,n3[19]);
    not g1708(n984 ,n3[45]);
    not g1709(n983 ,n3[54]);
    not g1710(n982 ,n3[7]);
    not g1711(n981 ,n3[32]);
    not g1712(n980 ,n3[57]);
    not g1713(n979 ,n5[37]);
    not g1714(n978 ,n5[50]);
    not g1715(n977 ,n3[27]);
    not g1716(n976 ,n4[30]);
    not g1717(n975 ,n3[36]);
    not g1718(n974 ,n5[43]);
    not g1719(n973 ,n4[37]);
    not g1720(n972 ,n5[10]);
    not g1721(n971 ,n4[41]);
    not g1722(n970 ,n4[36]);
    not g1723(n969 ,n3[8]);
    not g1724(n968 ,n5[49]);
    not g1725(n967 ,n4[44]);
    not g1726(n966 ,n5[30]);
    not g1727(n965 ,n5[34]);
    not g1728(n964 ,n4[61]);
    not g1729(n963 ,n5[27]);
    not g1730(n962 ,n4[48]);
    not g1731(n961 ,n4[56]);
    not g1732(n960 ,n3[21]);
    not g1733(n959 ,n5[48]);
    not g1734(n958 ,n3[20]);
    not g1735(n957 ,n3[23]);
    not g1736(n956 ,n4[13]);
    not g1737(n955 ,n4[42]);
    not g1738(n954 ,n3[53]);
    not g1739(n953 ,n4[22]);
    not g1740(n952 ,n3[40]);
    not g1741(n951 ,n5[58]);
    not g1742(n950 ,n5[23]);
    not g1743(n949 ,n5[47]);
    not g1744(n948 ,n5[15]);
    not g1745(n947 ,n5[38]);
    not g1746(n946 ,n5[63]);
    not g1747(n945 ,n4[29]);
    not g1748(n944 ,n3[33]);
    not g1749(n943 ,n3[10]);
    not g1750(n942 ,n4[57]);
    not g1751(n941 ,n4[45]);
    not g1752(n940 ,n4[4]);
    not g1753(n939 ,n5[17]);
    not g1754(n938 ,n3[29]);
    not g1755(n937 ,n3[46]);
    not g1756(n936 ,n4[51]);
    not g1757(n935 ,n4[46]);
    not g1758(n934 ,n3[18]);
    not g1759(n933 ,n3[37]);
    not g1760(n932 ,n3[50]);
    not g1761(n931 ,n4[58]);
    not g1762(n930 ,n5[22]);
    not g1763(n929 ,n4[15]);
    not g1764(n928 ,n3[14]);
    not g1765(n927 ,n3[48]);
    not g1766(n926 ,n5[12]);
    not g1767(n925 ,n3[26]);
    not g1768(n924 ,n5[53]);
    not g1769(n923 ,n5[39]);
    not g1770(n922 ,n5[20]);
    not g1771(n921 ,n3[31]);
    not g1772(n920 ,n3[61]);
    not g1773(n919 ,n5[14]);
    not g1774(n918 ,n5[40]);
    not g1775(n917 ,n4[62]);
    not g1776(n916 ,n5[7]);
    not g1777(n915 ,n4[14]);
    not g1778(n914 ,n5[52]);
    not g1779(n913 ,n4[16]);
    not g1780(n912 ,n3[52]);
    not g1781(n911 ,n5[8]);
    not g1782(n910 ,n5[55]);
    not g1783(n909 ,n3[11]);
    not g1784(n908 ,n4[21]);
    not g1785(n907 ,n3[43]);
    not g1786(n906 ,n4[43]);
    not g1787(n905 ,n3[30]);
    not g1788(n904 ,n3[47]);
    not g1789(n903 ,n5[11]);
    not g1790(n902 ,n3[9]);
    not g1791(n901 ,n4[27]);
    not g1792(n900 ,n3[42]);
    not g1793(n899 ,n5[31]);
    not g1794(n898 ,n3[39]);
    not g1795(n897 ,n3[22]);
    not g1796(n896 ,n3[60]);
    not g1797(n895 ,n8[1]);
    not g1798(n894 ,n5[18]);
    not g1799(n893 ,n3[44]);
    not g1800(n892 ,n3[59]);
    not g1801(n891 ,n4[53]);
    not g1802(n890 ,n3[28]);
    not g1803(n889 ,n5[57]);
    not g1804(n888 ,n5[42]);
    not g1805(n887 ,n5[13]);
    not g1806(n886 ,n3[51]);
    not g1807(n885 ,n4[40]);
    not g1808(n884 ,n4[19]);
    not g1809(n883 ,n5[4]);
    not g1810(n882 ,n5[51]);
    not g1811(n881 ,n3[16]);
    not g1812(n880 ,n4[34]);
    not g1813(n879 ,n4[20]);
    not g1814(n878 ,n5[5]);
    not g1815(n877 ,n3[38]);
    not g1816(n876 ,n4[24]);
    not g1817(n875 ,n5[45]);
    not g1818(n874 ,n3[62]);
    not g1819(n873 ,n3[63]);
    not g1820(n872 ,n4[32]);
    not g1821(n871 ,n8[3]);
    not g1822(n870 ,n4[31]);
    not g1823(n869 ,n3[4]);
    not g1824(n868 ,n3[56]);
    not g1825(n867 ,n5[16]);
    not g1826(n866 ,n5[21]);
    not g1827(n865 ,n3[58]);
    not g1828(n864 ,n4[33]);
    not g1829(n863 ,n5[41]);
    not g1830(n862 ,n5[24]);
    not g1831(n861 ,n8[2]);
    not g1832(n860 ,n3[17]);
    not g1833(n859 ,n4[18]);
    not g1834(n858 ,n3[12]);
    not g1835(n857 ,n4[26]);
    not g1836(n856 ,n4[12]);
    not g1837(n855 ,n5[60]);
    not g1838(n854 ,n3[35]);
    not g1839(n853 ,n4[47]);
    not g1840(n852 ,n4[11]);
    not g1841(n851 ,n5[61]);
    not g1842(n850 ,n5[6]);
    not g1843(n849 ,n4[10]);
    not g1844(n848 ,n3[5]);
    not g1845(n847 ,n4[55]);
    not g1846(n846 ,n4[9]);
    not g1847(n845 ,n5[46]);
    not g1848(n844 ,n5[32]);
    not g1849(n843 ,n3[49]);
    not g1850(n842 ,n4[8]);
    not g1851(n841 ,n3[34]);
    not g1852(n840 ,n3[13]);
    not g1853(n839 ,n3[41]);
    not g1854(n838 ,n4[7]);
    not g1855(n837 ,n4[63]);
    not g1856(n836 ,n5[62]);
    not g1857(n835 ,n4[6]);
    not g1858(n834 ,n4[23]);
    not g1859(n833 ,n5[26]);
    not g1860(n832 ,n4[28]);
    not g1861(n831 ,n4[5]);
    not g1862(n830 ,n8[0]);
    not g1863(n829 ,n3[2]);
    not g1864(n828 ,n3[0]);
    not g1865(n827 ,n3[1]);
    not g1866(n826 ,n4[3]);
    not g1867(n825 ,n5[1]);
    not g1868(n824 ,n5[2]);
    not g1869(n823 ,n4[2]);
    not g1870(n822 ,n5[0]);
    not g1871(n821 ,n5[3]);
    not g1872(n820 ,n4[1]);
    not g1873(n819 ,n4[0]);
    not g1874(n818 ,n3[3]);
    not g1875(n528 ,n2068);
    buf g1876(n7[1] ,n2068);
    not g1877(n817 ,n2069);
    buf g1878(n7[2] ,n2069);
    not g1879(n816 ,n7[0]);
    not g1880(n815 ,n2[14]);
    not g1881(n814 ,n2350);
    not g1882(n813 ,n2[104]);
    not g1883(n812 ,n2[117]);
    not g1884(n811 ,n2[96]);
    not g1885(n810 ,n2389);
    not g1886(n809 ,n2372);
    not g1887(n808 ,n2405);
    not g1888(n807 ,n2[99]);
    not g1889(n806 ,n2382);
    not g1890(n805 ,n2396);
    not g1891(n804 ,n2[25]);
    not g1892(n803 ,n2367);
    not g1893(n802 ,n2608);
    not g1894(n801 ,n2[13]);
    not g1895(n800 ,n2[102]);
    not g1896(n799 ,n2361);
    not g1897(n798 ,n2374);
    not g1898(n797 ,n2373);
    not g1899(n796 ,n2387);
    not g1900(n795 ,n2410);
    not g1901(n794 ,n2366);
    not g1902(n793 ,n2[11]);
    not g1903(n792 ,n2[106]);
    not g1904(n791 ,n2363);
    not g1905(n790 ,n2[98]);
    not g1906(n789 ,n2348);
    not g1907(n788 ,n2370);
    not g1908(n787 ,n2392);
    not g1909(n786 ,n2371);
    not g1910(n785 ,n2[17]);
    not g1911(n784 ,n2400);
    not g1912(n783 ,n2[101]);
    not g1913(n782 ,n2[123]);
    not g1914(n781 ,n2[10]);
    not g1915(n780 ,n2[108]);
    not g1916(n779 ,n2359);
    not g1917(n778 ,n2[24]);
    not g1918(n777 ,n2365);
    not g1919(n776 ,n2347);
    not g1920(n775 ,n2378);
    not g1921(n774 ,n2[27]);
    not g1922(n773 ,n2[6]);
    not g1923(n772 ,n2379);
    not g1924(n771 ,n2[4]);
    not g1925(n770 ,n2[21]);
    not g1926(n769 ,n2351);
    not g1927(n768 ,n2[120]);
    not g1928(n767 ,n2369);
    not g1929(n766 ,n2[110]);
    not g1930(n765 ,n2[125]);
    not g1931(n764 ,n2[107]);
    not g1932(n763 ,n2402);
    not g1933(n762 ,n2[8]);
    not g1934(n761 ,n2390);
    not g1935(n760 ,n2[97]);
    not g1936(n759 ,n2[127]);
    not g1937(n758 ,n2[109]);
    not g1938(n757 ,n2375);
    not g1939(n756 ,n2[16]);
    not g1940(n755 ,n2352);
    not g1941(n754 ,n2[18]);
    not g1942(n753 ,n2[105]);
    not g1943(n752 ,n2397);
    not g1944(n751 ,n2384);
    not g1945(n750 ,n2380);
    not g1946(n749 ,n2356);
    not g1947(n748 ,n2[119]);
    not g1948(n747 ,n2399);
    not g1949(n746 ,n2385);
    not g1950(n745 ,n2409);
    not g1951(n744 ,n2[111]);
    not g1952(n743 ,n2364);
    not g1953(n742 ,n2404);
    not g1954(n741 ,n2[116]);
    not g1955(n740 ,n2[9]);
    not g1956(n739 ,n2377);
    not g1957(n738 ,n2368);
    not g1958(n737 ,n2609);
    not g1959(n736 ,n2[23]);
    not g1960(n735 ,n2357);
    not g1961(n734 ,n2[113]);
    not g1962(n733 ,n2406);
    not g1963(n732 ,n2349);
    not g1964(n731 ,n2408);
    not g1965(n730 ,n2[100]);
    not g1966(n729 ,n2[12]);
    not g1967(n728 ,n2391);
    not g1968(n727 ,n2[20]);
    not g1969(n726 ,n2381);
    not g1970(n725 ,n2403);
    not g1971(n724 ,n2[115]);
    not g1972(n723 ,n2[112]);
    not g1973(n722 ,n2[118]);
    not g1974(n721 ,n2[15]);
    not g1975(n720 ,n2[5]);
    not g1976(n719 ,n2395);
    not g1977(n718 ,n2355);
    not g1978(n717 ,n2[122]);
    not g1979(n716 ,n2[7]);
    not g1980(n715 ,n2[114]);
    not g1981(n714 ,n2401);
    not g1982(n713 ,n2[124]);
    not g1983(n712 ,n2[103]);
    not g1984(n711 ,n2407);
    not g1985(n710 ,n2[121]);
    not g1986(n709 ,n2[22]);
    not g1987(n708 ,n2[126]);
    not g1988(n707 ,n2388);
    not g1989(n706 ,n2607);
    not g1990(n705 ,n2398);
    not g1991(n704 ,n2383);
    not g1992(n703 ,n2376);
    not g1993(n702 ,n2[26]);
    not g1994(n701 ,n2[19]);
    not g1995(n700 ,n2362);
    not g1996(n699 ,n2394);
    not g1997(n698 ,n2354);
    not g1998(n697 ,n2360);
    not g1999(n696 ,n2386);
    not g2000(n695 ,n2353);
    not g2001(n694 ,n2393);
    not g2002(n693 ,n2358);
    not g2003(n692 ,n2438);
    not g2004(n691 ,n2[83]);
    not g2005(n690 ,n2432);
    not g2006(n689 ,n2[59]);
    not g2007(n688 ,n2460);
    not g2008(n687 ,n2[74]);
    not g2009(n686 ,n2466);
    not g2010(n685 ,n2461);
    not g2011(n684 ,n2420);
    not g2012(n683 ,n2425);
    not g2013(n682 ,n2[0]);
    not g2014(n681 ,n2416);
    not g2015(n680 ,n2424);
    not g2016(n679 ,n2448);
    not g2017(n678 ,n2435);
    not g2018(n677 ,n2[88]);
    not g2019(n676 ,n2[68]);
    not g2020(n675 ,n2436);
    not g2021(n674 ,n2440);
    not g2022(n673 ,n2433);
    not g2023(n672 ,n2427);
    not g2024(n671 ,n2418);
    not g2025(n670 ,n2[58]);
    not g2026(n669 ,n2454);
    not g2027(n668 ,n2417);
    not g2028(n667 ,n2465);
    not g2029(n666 ,n2413);
    not g2030(n665 ,n2[60]);
    not g2031(n664 ,n2473);
    not g2032(n663 ,n2[50]);
    not g2033(n662 ,n2[29]);
    not g2034(n661 ,n2468);
    not g2035(n660 ,n2469);
    not g2036(n659 ,n2[54]);
    not g2037(n658 ,n2[32]);
    not g2038(n657 ,n2[34]);
    not g2039(n656 ,n2462);
    not g2040(n655 ,n2[70]);
    not g2041(n654 ,n2[73]);
    not g2042(n653 ,n2[39]);
    not g2043(n652 ,n2[46]);
    not g2044(n651 ,n2[78]);
    not g2045(n650 ,n2442);
    not g2046(n649 ,n2459);
    not g2047(n648 ,n2430);
    not g2048(n647 ,n2[94]);
    not g2049(n646 ,n2471);
    not g2050(n645 ,n2423);
    not g2051(n644 ,n2464);
    not g2052(n643 ,n2[44]);
    not g2053(n642 ,n2470);
    not g2054(n641 ,n2411);
    not g2055(n640 ,n2431);
    not g2056(n639 ,n2[42]);
    not g2057(n638 ,n2449);
    not g2058(n637 ,n2[90]);
    not g2059(n636 ,n2[38]);
    not g2060(n635 ,n2[71]);
    not g2061(n634 ,n2[49]);
    not g2062(n633 ,n2[87]);
    not g2063(n632 ,n2474);
    not g2064(n631 ,n2414);
    not g2065(n630 ,n2415);
    not g2066(n629 ,n2[2]);
    not g2067(n628 ,n2[28]);
    not g2068(n627 ,n2[63]);
    not g2069(n626 ,n2426);
    not g2070(n625 ,n2434);
    not g2071(n624 ,n2[82]);
    not g2072(n623 ,n2463);
    not g2073(n622 ,n2[77]);
    not g2074(n621 ,n2452);
    not g2075(n620 ,n2451);
    not g2076(n619 ,n2[45]);
    not g2077(n618 ,n2[76]);
    not g2078(n617 ,n2421);
    not g2079(n616 ,n2[93]);
    not g2080(n615 ,n2412);
    not g2081(n614 ,n2457);
    not g2082(n613 ,n2[91]);
    not g2083(n612 ,n2[61]);
    not g2084(n611 ,n2[86]);
    not g2085(n610 ,n2[57]);
    not g2086(n609 ,n2444);
    not g2087(n608 ,n2[95]);
    not g2088(n607 ,n2455);
    not g2089(n606 ,n2[80]);
    not g2090(n605 ,n2458);
    not g2091(n604 ,n2[69]);
    not g2092(n603 ,n2[30]);
    not g2093(n602 ,n2[31]);
    not g2094(n601 ,n2456);
    not g2095(n600 ,n2445);
    not g2096(n599 ,n2[92]);
    not g2097(n598 ,n2453);
    not g2098(n597 ,n2[3]);
    not g2099(n596 ,n2429);
    not g2100(n595 ,n2[35]);
    not g2101(n594 ,n2446);
    not g2102(n593 ,n2[53]);
    not g2103(n592 ,n2[33]);
    not g2104(n591 ,n2[47]);
    not g2105(n590 ,n2419);
    not g2106(n589 ,n2[56]);
    not g2107(n588 ,n2[43]);
    not g2108(n587 ,n2422);
    not g2109(n586 ,n2[81]);
    not g2110(n585 ,n2[40]);
    not g2111(n584 ,n2[1]);
    not g2112(n583 ,n2428);
    not g2113(n582 ,n2[48]);
    not g2114(n581 ,n2467);
    not g2115(n580 ,n2[84]);
    not g2116(n579 ,n2443);
    not g2117(n578 ,n2[79]);
    not g2118(n577 ,n2450);
    not g2119(n576 ,n2[62]);
    not g2120(n575 ,n2[72]);
    not g2121(n574 ,n2[51]);
    not g2122(n573 ,n2[37]);
    not g2123(n572 ,n2[75]);
    not g2124(n571 ,n2447);
    not g2125(n570 ,n2[52]);
    not g2126(n569 ,n2[36]);
    not g2127(n568 ,n2441);
    not g2128(n567 ,n2439);
    not g2129(n566 ,n2437);
    not g2130(n565 ,n2472);
    not g2131(n564 ,n2[41]);
    not g2132(n563 ,n2[89]);
    not g2133(n562 ,n2[55]);
    not g2134(n561 ,n2[85]);
    not g2135(n560 ,n2[65]);
    not g2136(n559 ,n2[67]);
    not g2137(n558 ,n2[66]);
    not g2138(n557 ,n2[64]);
    not g2139(n556 ,n6[1]);
    not g2140(n555 ,n6[2]);
    not g2141(n554 ,n6[0]);
    not g2142(n553 ,n6[3]);
    not g2143(n552 ,n2346);
    not g2144(n551 ,n2346);
    not g2145(n550 ,n2346);
    not g2146(n549 ,n2346);
    not g2147(n548 ,n2346);
    not g2148(n547 ,n2346);
    not g2149(n546 ,n2346);
    not g2150(n545 ,n2346);
    not g2151(n544 ,n2346);
    not g2152(n543 ,n2346);
    not g2153(n542 ,n2346);
    xnor g2154(n2602 ,n80 ,n268);
    nor g2155(n268 ,n53 ,n267);
    xnor g2156(n2601 ,n96 ,n266);
    nor g2157(n267 ,n96 ,n266);
    nor g2158(n266 ,n42 ,n265);
    xnor g2159(n2600 ,n117 ,n264);
    nor g2160(n265 ,n117 ,n264);
    nor g2161(n264 ,n71 ,n263);
    xnor g2162(n2599 ,n99 ,n262);
    nor g2163(n263 ,n99 ,n262);
    nor g2164(n262 ,n45 ,n261);
    xnor g2165(n2598 ,n104 ,n260);
    nor g2166(n261 ,n104 ,n260);
    nor g2167(n260 ,n57 ,n259);
    xnor g2168(n2597 ,n126 ,n258);
    nor g2169(n259 ,n126 ,n258);
    nor g2170(n258 ,n38 ,n257);
    xnor g2171(n2596 ,n109 ,n256);
    nor g2172(n257 ,n109 ,n256);
    nor g2173(n256 ,n72 ,n255);
    xnor g2174(n2595 ,n98 ,n254);
    nor g2175(n255 ,n98 ,n254);
    nor g2176(n254 ,n18 ,n253);
    xnor g2177(n2594 ,n137 ,n252);
    nor g2178(n253 ,n137 ,n252);
    nor g2179(n252 ,n37 ,n251);
    xnor g2180(n2593 ,n91 ,n250);
    nor g2181(n251 ,n91 ,n250);
    nor g2182(n250 ,n64 ,n249);
    xnor g2183(n2592 ,n132 ,n248);
    nor g2184(n249 ,n132 ,n248);
    nor g2185(n248 ,n49 ,n247);
    xnor g2186(n2591 ,n127 ,n246);
    nor g2187(n247 ,n127 ,n246);
    nor g2188(n246 ,n41 ,n245);
    xnor g2189(n2590 ,n121 ,n244);
    nor g2190(n245 ,n121 ,n244);
    nor g2191(n244 ,n33 ,n243);
    xnor g2192(n2589 ,n113 ,n242);
    nor g2193(n243 ,n113 ,n242);
    nor g2194(n242 ,n29 ,n241);
    xnor g2195(n2588 ,n102 ,n240);
    nor g2196(n241 ,n102 ,n240);
    nor g2197(n240 ,n23 ,n239);
    xnor g2198(n2587 ,n111 ,n238);
    nor g2199(n239 ,n111 ,n238);
    nor g2200(n238 ,n16 ,n237);
    xnor g2201(n2586 ,n87 ,n236);
    nor g2202(n237 ,n87 ,n236);
    nor g2203(n236 ,n59 ,n235);
    xnor g2204(n2585 ,n82 ,n234);
    nor g2205(n235 ,n82 ,n234);
    nor g2206(n234 ,n77 ,n233);
    xnor g2207(n2584 ,n84 ,n232);
    nor g2208(n233 ,n84 ,n232);
    nor g2209(n232 ,n58 ,n231);
    xnor g2210(n2583 ,n90 ,n230);
    nor g2211(n231 ,n90 ,n230);
    nor g2212(n230 ,n65 ,n229);
    xnor g2213(n2582 ,n139 ,n228);
    nor g2214(n229 ,n139 ,n228);
    nor g2215(n228 ,n32 ,n227);
    xnor g2216(n2581 ,n135 ,n226);
    nor g2217(n227 ,n135 ,n226);
    nor g2218(n226 ,n51 ,n225);
    xnor g2219(n2580 ,n130 ,n224);
    nor g2220(n225 ,n130 ,n224);
    nor g2221(n224 ,n27 ,n223);
    xnor g2222(n2579 ,n100 ,n222);
    nor g2223(n223 ,n100 ,n222);
    nor g2224(n222 ,n43 ,n221);
    xnor g2225(n2578 ,n124 ,n220);
    nor g2226(n221 ,n124 ,n220);
    nor g2227(n220 ,n68 ,n219);
    xnor g2228(n2577 ,n120 ,n218);
    nor g2229(n219 ,n120 ,n218);
    nor g2230(n218 ,n35 ,n217);
    xnor g2231(n2576 ,n115 ,n216);
    nor g2232(n217 ,n115 ,n216);
    nor g2233(n216 ,n40 ,n215);
    xnor g2234(n2575 ,n112 ,n214);
    nor g2235(n215 ,n112 ,n214);
    nor g2236(n214 ,n55 ,n213);
    xnor g2237(n2574 ,n110 ,n212);
    nor g2238(n213 ,n110 ,n212);
    nor g2239(n212 ,n19 ,n211);
    xnor g2240(n2573 ,n106 ,n210);
    nor g2241(n211 ,n106 ,n210);
    nor g2242(n210 ,n25 ,n209);
    xnor g2243(n2572 ,n101 ,n208);
    nor g2244(n209 ,n101 ,n208);
    nor g2245(n208 ,n48 ,n207);
    xnor g2246(n2571 ,n94 ,n206);
    nor g2247(n207 ,n94 ,n206);
    nor g2248(n206 ,n74 ,n205);
    xnor g2249(n2570 ,n89 ,n204);
    nor g2250(n205 ,n89 ,n204);
    nor g2251(n204 ,n75 ,n203);
    xnor g2252(n2569 ,n86 ,n202);
    nor g2253(n203 ,n86 ,n202);
    nor g2254(n202 ,n17 ,n201);
    xnor g2255(n2568 ,n81 ,n200);
    nor g2256(n201 ,n81 ,n200);
    nor g2257(n200 ,n54 ,n199);
    xnor g2258(n2567 ,n83 ,n198);
    nor g2259(n199 ,n83 ,n198);
    nor g2260(n198 ,n69 ,n197);
    xnor g2261(n2566 ,n85 ,n196);
    nor g2262(n197 ,n85 ,n196);
    nor g2263(n196 ,n66 ,n195);
    xnor g2264(n2565 ,n88 ,n194);
    nor g2265(n195 ,n88 ,n194);
    nor g2266(n194 ,n46 ,n193);
    xnor g2267(n2564 ,n93 ,n192);
    nor g2268(n193 ,n93 ,n192);
    nor g2269(n192 ,n44 ,n191);
    xnor g2270(n2563 ,n92 ,n190);
    nor g2271(n191 ,n92 ,n190);
    nor g2272(n190 ,n20 ,n189);
    xnor g2273(n2562 ,n141 ,n188);
    nor g2274(n189 ,n141 ,n188);
    nor g2275(n188 ,n63 ,n187);
    xnor g2276(n2561 ,n138 ,n186);
    nor g2277(n187 ,n138 ,n186);
    nor g2278(n186 ,n60 ,n185);
    xnor g2279(n2560 ,n136 ,n184);
    nor g2280(n185 ,n136 ,n184);
    nor g2281(n184 ,n56 ,n183);
    xnor g2282(n2559 ,n134 ,n182);
    nor g2283(n183 ,n134 ,n182);
    nor g2284(n182 ,n52 ,n181);
    xnor g2285(n2558 ,n133 ,n180);
    nor g2286(n181 ,n133 ,n180);
    nor g2287(n180 ,n50 ,n179);
    xnor g2288(n2557 ,n131 ,n178);
    nor g2289(n179 ,n131 ,n178);
    nor g2290(n178 ,n31 ,n177);
    xnor g2291(n2556 ,n128 ,n176);
    nor g2292(n177 ,n128 ,n176);
    nor g2293(n176 ,n22 ,n175);
    xnor g2294(n2555 ,n107 ,n174);
    nor g2295(n175 ,n107 ,n174);
    nor g2296(n174 ,n24 ,n173);
    xnor g2297(n2554 ,n125 ,n172);
    nor g2298(n173 ,n125 ,n172);
    nor g2299(n172 ,n67 ,n171);
    xnor g2300(n2553 ,n123 ,n170);
    nor g2301(n171 ,n123 ,n170);
    nor g2302(n170 ,n39 ,n169);
    xnor g2303(n2552 ,n122 ,n168);
    nor g2304(n169 ,n122 ,n168);
    nor g2305(n168 ,n36 ,n167);
    xnor g2306(n2551 ,n119 ,n166);
    nor g2307(n167 ,n119 ,n166);
    nor g2308(n166 ,n70 ,n165);
    xnor g2309(n2550 ,n118 ,n164);
    nor g2310(n165 ,n118 ,n164);
    nor g2311(n164 ,n34 ,n163);
    xnor g2312(n2549 ,n116 ,n162);
    nor g2313(n163 ,n116 ,n162);
    nor g2314(n162 ,n47 ,n161);
    xnor g2315(n2548 ,n114 ,n160);
    nor g2316(n161 ,n114 ,n160);
    nor g2317(n160 ,n30 ,n159);
    xnor g2318(n2547 ,n129 ,n158);
    nor g2319(n159 ,n129 ,n158);
    nor g2320(n158 ,n61 ,n157);
    xnor g2321(n2546 ,n95 ,n156);
    nor g2322(n157 ,n95 ,n156);
    nor g2323(n156 ,n28 ,n155);
    xnor g2324(n2545 ,n140 ,n154);
    nor g2325(n155 ,n140 ,n154);
    nor g2326(n154 ,n26 ,n153);
    xnor g2327(n2544 ,n108 ,n152);
    nor g2328(n153 ,n108 ,n152);
    nor g2329(n152 ,n76 ,n151);
    xnor g2330(n2543 ,n105 ,n150);
    nor g2331(n151 ,n105 ,n150);
    nor g2332(n150 ,n73 ,n149);
    xor g2333(n2603 ,n103 ,n147);
    nor g2334(n149 ,n103 ,n148);
    not g2335(n148 ,n147);
    nor g2336(n147 ,n62 ,n146);
    xnor g2337(n2604 ,n142 ,n144);
    nor g2338(n146 ,n142 ,n145);
    not g2339(n145 ,n144);
    nor g2340(n144 ,n21 ,n143);
    xnor g2341(n2605 ,n97 ,n79);
    nor g2342(n143 ,n79 ,n97);
    nor g2343(n2606 ,n79 ,n78);
    xnor g2344(n142 ,n2[2] ,n2[66]);
    xnor g2345(n141 ,n2[23] ,n2[87]);
    xnor g2346(n140 ,n2[6] ,n2[70]);
    xnor g2347(n139 ,n2[43] ,n2[107]);
    xnor g2348(n138 ,n2[22] ,n2[86]);
    xnor g2349(n137 ,n2[55] ,n2[119]);
    xnor g2350(n136 ,n2[21] ,n2[85]);
    xnor g2351(n135 ,n2[42] ,n2[106]);
    xnor g2352(n134 ,n2[20] ,n2[84]);
    xnor g2353(n133 ,n2[19] ,n2[83]);
    xnor g2354(n132 ,n2[53] ,n2[117]);
    xnor g2355(n131 ,n2[18] ,n2[82]);
    xnor g2356(n130 ,n2[41] ,n2[105]);
    xnor g2357(n129 ,n2[8] ,n2[72]);
    xnor g2358(n128 ,n2[17] ,n2[81]);
    xnor g2359(n127 ,n2[52] ,n2[116]);
    xnor g2360(n126 ,n2[58] ,n2[122]);
    xnor g2361(n125 ,n2[15] ,n2[79]);
    xnor g2362(n124 ,n2[39] ,n2[103]);
    xnor g2363(n123 ,n2[14] ,n2[78]);
    xnor g2364(n122 ,n2[13] ,n2[77]);
    xnor g2365(n121 ,n2[51] ,n2[115]);
    xnor g2366(n120 ,n2[38] ,n2[102]);
    xnor g2367(n119 ,n2[12] ,n2[76]);
    xnor g2368(n118 ,n2[11] ,n2[75]);
    xnor g2369(n117 ,n2[61] ,n2[125]);
    xnor g2370(n116 ,n2[10] ,n2[74]);
    xnor g2371(n115 ,n2[37] ,n2[101]);
    xnor g2372(n114 ,n2[9] ,n2[73]);
    xnor g2373(n113 ,n2[50] ,n2[114]);
    xnor g2374(n112 ,n2[36] ,n2[100]);
    xnor g2375(n111 ,n2[48] ,n2[112]);
    xnor g2376(n110 ,n2[35] ,n2[99]);
    xnor g2377(n109 ,n2[57] ,n2[121]);
    xnor g2378(n108 ,n2[5] ,n2[69]);
    xnor g2379(n107 ,n2[16] ,n2[80]);
    xnor g2380(n106 ,n2[34] ,n2[98]);
    xnor g2381(n105 ,n2[4] ,n2[68]);
    xnor g2382(n104 ,n2[59] ,n2[123]);
    xnor g2383(n103 ,n2[3] ,n2[67]);
    xnor g2384(n102 ,n2[49] ,n2[113]);
    xnor g2385(n101 ,n2[33] ,n2[97]);
    xnor g2386(n100 ,n2[40] ,n2[104]);
    xnor g2387(n99 ,n2[60] ,n2[124]);
    xnor g2388(n98 ,n2[56] ,n2[120]);
    xnor g2389(n97 ,n2[1] ,n2[65]);
    xnor g2390(n96 ,n2[62] ,n2[126]);
    xnor g2391(n95 ,n2[7] ,n2[71]);
    xnor g2392(n94 ,n2[32] ,n2[96]);
    xnor g2393(n93 ,n2[25] ,n2[89]);
    xnor g2394(n92 ,n2[24] ,n2[88]);
    xnor g2395(n91 ,n2[54] ,n2[118]);
    xnor g2396(n90 ,n2[44] ,n2[108]);
    xnor g2397(n89 ,n2[31] ,n2[95]);
    xnor g2398(n88 ,n2[26] ,n2[90]);
    xnor g2399(n87 ,n2[47] ,n2[111]);
    xnor g2400(n86 ,n2[30] ,n2[94]);
    xnor g2401(n85 ,n2[27] ,n2[91]);
    xnor g2402(n84 ,n2[45] ,n2[109]);
    xnor g2403(n83 ,n2[28] ,n2[92]);
    xnor g2404(n82 ,n2[46] ,n2[110]);
    xnor g2405(n81 ,n2[29] ,n2[93]);
    xnor g2406(n80 ,n2[63] ,n2[127]);
    nor g2407(n78 ,n2[0] ,n2[64]);
    nor g2408(n77 ,n2[45] ,n2[109]);
    nor g2409(n76 ,n2[4] ,n2[68]);
    nor g2410(n75 ,n2[30] ,n2[94]);
    nor g2411(n74 ,n2[31] ,n2[95]);
    nor g2412(n73 ,n2[3] ,n2[67]);
    nor g2413(n72 ,n2[56] ,n2[120]);
    nor g2414(n71 ,n2[60] ,n2[124]);
    nor g2415(n70 ,n2[11] ,n2[75]);
    nor g2416(n69 ,n2[27] ,n2[91]);
    nor g2417(n68 ,n2[38] ,n2[102]);
    nor g2418(n67 ,n2[14] ,n2[78]);
    nor g2419(n66 ,n2[26] ,n2[90]);
    nor g2420(n65 ,n2[43] ,n2[107]);
    nor g2421(n64 ,n2[53] ,n2[117]);
    nor g2422(n63 ,n2[22] ,n2[86]);
    nor g2423(n62 ,n14 ,n13);
    nor g2424(n61 ,n2[7] ,n2[71]);
    nor g2425(n60 ,n2[21] ,n2[85]);
    nor g2426(n59 ,n2[46] ,n2[110]);
    nor g2427(n58 ,n2[44] ,n2[108]);
    nor g2428(n57 ,n2[58] ,n2[122]);
    nor g2429(n56 ,n2[20] ,n2[84]);
    nor g2430(n55 ,n2[35] ,n2[99]);
    nor g2431(n54 ,n2[28] ,n2[92]);
    nor g2432(n53 ,n2[62] ,n2[126]);
    nor g2433(n52 ,n2[19] ,n2[83]);
    nor g2434(n51 ,n2[41] ,n2[105]);
    nor g2435(n50 ,n2[18] ,n2[82]);
    nor g2436(n49 ,n2[52] ,n2[116]);
    nor g2437(n48 ,n2[32] ,n2[96]);
    nor g2438(n79 ,n15 ,n12);
    nor g2439(n47 ,n2[9] ,n2[73]);
    nor g2440(n46 ,n2[25] ,n2[89]);
    nor g2441(n45 ,n2[59] ,n2[123]);
    nor g2442(n44 ,n2[24] ,n2[88]);
    nor g2443(n43 ,n2[39] ,n2[103]);
    nor g2444(n42 ,n2[61] ,n2[125]);
    nor g2445(n41 ,n2[51] ,n2[115]);
    nor g2446(n40 ,n2[36] ,n2[100]);
    nor g2447(n39 ,n2[13] ,n2[77]);
    nor g2448(n38 ,n2[57] ,n2[121]);
    nor g2449(n37 ,n2[54] ,n2[118]);
    nor g2450(n36 ,n2[12] ,n2[76]);
    nor g2451(n35 ,n2[37] ,n2[101]);
    nor g2452(n34 ,n2[10] ,n2[74]);
    nor g2453(n33 ,n2[50] ,n2[114]);
    nor g2454(n32 ,n2[42] ,n2[106]);
    nor g2455(n31 ,n2[17] ,n2[81]);
    nor g2456(n30 ,n2[8] ,n2[72]);
    nor g2457(n29 ,n2[49] ,n2[113]);
    nor g2458(n28 ,n2[6] ,n2[70]);
    nor g2459(n27 ,n2[40] ,n2[104]);
    nor g2460(n26 ,n2[5] ,n2[69]);
    nor g2461(n25 ,n2[33] ,n2[97]);
    nor g2462(n24 ,n2[15] ,n2[79]);
    nor g2463(n23 ,n2[48] ,n2[112]);
    nor g2464(n22 ,n2[16] ,n2[80]);
    nor g2465(n21 ,n2[1] ,n2[65]);
    nor g2466(n20 ,n2[23] ,n2[87]);
    nor g2467(n19 ,n2[34] ,n2[98]);
    nor g2468(n18 ,n2[55] ,n2[119]);
    nor g2469(n17 ,n2[29] ,n2[93]);
    nor g2470(n16 ,n2[47] ,n2[111]);
    not g2471(n15 ,n2[0]);
    not g2472(n14 ,n2[2]);
    not g2473(n13 ,n2[66]);
    not g2474(n12 ,n2[64]);
    xor g2475(n2474 ,n2542 ,n519);
    nor g2476(n2468 ,n504 ,n517);
    nor g2477(n2473 ,n518 ,n519);
    xor g2478(n2470 ,n2538 ,n516);
    nor g2479(n519 ,n279 ,n514);
    nor g2480(n518 ,n2541 ,n513);
    nor g2481(n517 ,n2536 ,n515);
    nor g2482(n2472 ,n512 ,n513);
    nor g2483(n2469 ,n511 ,n516);
    xor g2484(n2467 ,n2535 ,n509);
    xor g2485(n2466 ,n2534 ,n508);
    xor g2486(n2464 ,n2532 ,n503);
    nor g2487(n516 ,n299 ,n505);
    nor g2488(n515 ,n303 ,n510);
    not g2489(n514 ,n513);
    nor g2490(n513 ,n327 ,n507);
    nor g2491(n512 ,n2540 ,n506);
    nor g2492(n511 ,n2537 ,n504);
    nor g2493(n2462 ,n496 ,n499);
    nor g2494(n2471 ,n502 ,n506);
    nor g2495(n2465 ,n501 ,n508);
    nor g2496(n2463 ,n500 ,n503);
    not g2497(n510 ,n509);
    not g2498(n507 ,n506);
    not g2499(n505 ,n504);
    nor g2500(n509 ,n344 ,n497);
    nor g2501(n508 ,n300 ,n493);
    nor g2502(n506 ,n321 ,n495);
    nor g2503(n504 ,n348 ,n497);
    nor g2504(n503 ,n302 ,n497);
    nor g2505(n502 ,n2539 ,n494);
    nor g2506(n501 ,n2533 ,n492);
    nor g2507(n500 ,n2531 ,n496);
    nor g2508(n499 ,n2530 ,n498);
    xor g2509(n2461 ,n2529 ,n488);
    xor g2510(n2460 ,n2528 ,n490);
    nor g2511(n498 ,n270 ,n489);
    not g2512(n497 ,n496);
    nor g2513(n496 ,n337 ,n489);
    not g2514(n495 ,n494);
    nor g2515(n494 ,n352 ,n491);
    not g2516(n493 ,n492);
    nor g2517(n492 ,n334 ,n487);
    nor g2518(n2459 ,n486 ,n490);
    or g2519(n491 ,n273 ,n485);
    nor g2520(n490 ,n272 ,n485);
    not g2521(n489 ,n488);
    nor g2522(n488 ,n336 ,n485);
    or g2523(n487 ,n341 ,n485);
    nor g2524(n486 ,n2527 ,n484);
    xor g2525(n2458 ,n2526 ,n482);
    not g2526(n485 ,n484);
    nor g2527(n484 ,n269 ,n483);
    nor g2528(n2457 ,n481 ,n482);
    not g2529(n483 ,n482);
    nor g2530(n482 ,n297 ,n480);
    nor g2531(n481 ,n2525 ,n479);
    nor g2532(n2456 ,n478 ,n479);
    not g2533(n480 ,n479);
    nor g2534(n479 ,n290 ,n477);
    nor g2535(n478 ,n2524 ,n476);
    nor g2536(n2455 ,n475 ,n476);
    not g2537(n477 ,n476);
    nor g2538(n476 ,n320 ,n474);
    nor g2539(n475 ,n2523 ,n473);
    nor g2540(n2454 ,n472 ,n473);
    not g2541(n474 ,n473);
    nor g2542(n473 ,n326 ,n471);
    nor g2543(n472 ,n2522 ,n470);
    nor g2544(n2453 ,n469 ,n470);
    not g2545(n471 ,n470);
    nor g2546(n470 ,n295 ,n468);
    nor g2547(n469 ,n2521 ,n467);
    nor g2548(n2452 ,n466 ,n467);
    not g2549(n468 ,n467);
    nor g2550(n467 ,n310 ,n465);
    nor g2551(n466 ,n2520 ,n464);
    nor g2552(n2451 ,n463 ,n464);
    not g2553(n465 ,n464);
    nor g2554(n464 ,n313 ,n462);
    nor g2555(n463 ,n2519 ,n461);
    nor g2556(n2450 ,n460 ,n461);
    not g2557(n462 ,n461);
    nor g2558(n461 ,n311 ,n459);
    nor g2559(n460 ,n2518 ,n458);
    nor g2560(n2449 ,n457 ,n458);
    not g2561(n459 ,n458);
    nor g2562(n458 ,n308 ,n456);
    nor g2563(n457 ,n2517 ,n455);
    nor g2564(n2448 ,n454 ,n455);
    not g2565(n456 ,n455);
    nor g2566(n455 ,n325 ,n453);
    nor g2567(n454 ,n2516 ,n452);
    nor g2568(n2447 ,n451 ,n452);
    not g2569(n453 ,n452);
    nor g2570(n452 ,n275 ,n450);
    nor g2571(n451 ,n2515 ,n449);
    nor g2572(n2446 ,n448 ,n449);
    not g2573(n450 ,n449);
    nor g2574(n449 ,n278 ,n447);
    nor g2575(n448 ,n2514 ,n446);
    nor g2576(n2445 ,n445 ,n446);
    not g2577(n447 ,n446);
    nor g2578(n446 ,n329 ,n444);
    nor g2579(n445 ,n2513 ,n443);
    nor g2580(n2444 ,n442 ,n443);
    not g2581(n444 ,n443);
    nor g2582(n443 ,n285 ,n441);
    nor g2583(n442 ,n2512 ,n440);
    nor g2584(n2443 ,n439 ,n440);
    not g2585(n441 ,n440);
    nor g2586(n440 ,n277 ,n438);
    nor g2587(n439 ,n2511 ,n437);
    nor g2588(n2442 ,n436 ,n437);
    not g2589(n438 ,n437);
    nor g2590(n437 ,n322 ,n435);
    nor g2591(n436 ,n2510 ,n434);
    nor g2592(n2441 ,n433 ,n434);
    not g2593(n435 ,n434);
    nor g2594(n434 ,n283 ,n432);
    nor g2595(n433 ,n2509 ,n431);
    nor g2596(n2440 ,n430 ,n431);
    not g2597(n432 ,n431);
    nor g2598(n431 ,n280 ,n429);
    nor g2599(n430 ,n2508 ,n428);
    nor g2600(n2439 ,n427 ,n428);
    not g2601(n429 ,n428);
    nor g2602(n428 ,n284 ,n426);
    nor g2603(n427 ,n2507 ,n425);
    nor g2604(n2438 ,n424 ,n425);
    not g2605(n426 ,n425);
    nor g2606(n425 ,n307 ,n423);
    nor g2607(n424 ,n2506 ,n422);
    nor g2608(n2437 ,n421 ,n422);
    not g2609(n423 ,n422);
    nor g2610(n422 ,n312 ,n420);
    nor g2611(n421 ,n2505 ,n419);
    nor g2612(n2436 ,n418 ,n419);
    not g2613(n420 ,n419);
    nor g2614(n419 ,n328 ,n417);
    nor g2615(n418 ,n2504 ,n416);
    nor g2616(n2435 ,n415 ,n416);
    not g2617(n417 ,n416);
    nor g2618(n416 ,n276 ,n414);
    nor g2619(n415 ,n2503 ,n413);
    nor g2620(n2434 ,n412 ,n413);
    not g2621(n414 ,n413);
    nor g2622(n413 ,n305 ,n411);
    nor g2623(n412 ,n2502 ,n410);
    nor g2624(n2433 ,n409 ,n410);
    not g2625(n411 ,n410);
    nor g2626(n410 ,n287 ,n408);
    nor g2627(n409 ,n2501 ,n407);
    nor g2628(n2432 ,n406 ,n407);
    not g2629(n408 ,n407);
    nor g2630(n407 ,n318 ,n405);
    nor g2631(n406 ,n2500 ,n404);
    nor g2632(n2431 ,n403 ,n404);
    not g2633(n405 ,n404);
    nor g2634(n404 ,n323 ,n402);
    nor g2635(n403 ,n2499 ,n401);
    nor g2636(n2430 ,n400 ,n401);
    not g2637(n402 ,n401);
    nor g2638(n401 ,n289 ,n399);
    nor g2639(n400 ,n2498 ,n398);
    nor g2640(n2429 ,n397 ,n398);
    not g2641(n399 ,n398);
    nor g2642(n398 ,n316 ,n396);
    nor g2643(n397 ,n2497 ,n395);
    nor g2644(n2428 ,n394 ,n395);
    not g2645(n396 ,n395);
    nor g2646(n395 ,n291 ,n393);
    nor g2647(n394 ,n2496 ,n392);
    nor g2648(n2427 ,n391 ,n392);
    not g2649(n393 ,n392);
    nor g2650(n392 ,n288 ,n390);
    nor g2651(n391 ,n2495 ,n389);
    nor g2652(n2426 ,n388 ,n389);
    not g2653(n390 ,n389);
    nor g2654(n389 ,n292 ,n387);
    nor g2655(n388 ,n2494 ,n386);
    nor g2656(n2425 ,n385 ,n386);
    not g2657(n387 ,n386);
    nor g2658(n386 ,n306 ,n384);
    nor g2659(n385 ,n2493 ,n383);
    nor g2660(n2424 ,n382 ,n383);
    not g2661(n384 ,n383);
    nor g2662(n383 ,n294 ,n381);
    nor g2663(n382 ,n2492 ,n380);
    nor g2664(n2423 ,n379 ,n380);
    not g2665(n381 ,n380);
    nor g2666(n380 ,n309 ,n378);
    nor g2667(n379 ,n2491 ,n377);
    nor g2668(n2422 ,n376 ,n377);
    not g2669(n378 ,n377);
    nor g2670(n377 ,n324 ,n375);
    nor g2671(n376 ,n2490 ,n374);
    nor g2672(n2421 ,n373 ,n374);
    not g2673(n375 ,n374);
    nor g2674(n374 ,n282 ,n372);
    nor g2675(n373 ,n2489 ,n371);
    nor g2676(n2420 ,n370 ,n371);
    not g2677(n372 ,n371);
    nor g2678(n371 ,n314 ,n369);
    nor g2679(n370 ,n2488 ,n368);
    nor g2680(n2419 ,n367 ,n368);
    not g2681(n369 ,n368);
    nor g2682(n368 ,n317 ,n366);
    nor g2683(n367 ,n2487 ,n365);
    nor g2684(n2418 ,n364 ,n365);
    not g2685(n366 ,n365);
    nor g2686(n365 ,n298 ,n363);
    nor g2687(n364 ,n2486 ,n362);
    nor g2688(n2417 ,n361 ,n362);
    not g2689(n363 ,n362);
    nor g2690(n362 ,n315 ,n360);
    nor g2691(n361 ,n2485 ,n359);
    nor g2692(n2416 ,n358 ,n359);
    not g2693(n360 ,n359);
    nor g2694(n359 ,n281 ,n357);
    nor g2695(n358 ,n2484 ,n356);
    nor g2696(n2415 ,n355 ,n356);
    not g2697(n357 ,n356);
    nor g2698(n356 ,n296 ,n354);
    nor g2699(n355 ,n2483 ,n353);
    not g2700(n354 ,n353);
    nor g2701(n353 ,n331 ,n351);
    xnor g2702(n2414 ,n340 ,n349);
    or g2703(n352 ,n299 ,n350);
    nor g2704(n351 ,n340 ,n349);
    or g2705(n350 ,n341 ,n348);
    nor g2706(n349 ,n333 ,n347);
    xnor g2707(n2413 ,n338 ,n345);
    or g2708(n348 ,n303 ,n346);
    nor g2709(n347 ,n338 ,n345);
    or g2710(n346 ,n286 ,n344);
    nor g2711(n345 ,n332 ,n343);
    xnor g2712(n2412 ,n339 ,n335);
    or g2713(n344 ,n300 ,n342);
    nor g2714(n343 ,n335 ,n339);
    or g2715(n342 ,n271 ,n334);
    or g2716(n341 ,n337 ,n336);
    nor g2717(n2411 ,n335 ,n330);
    xnor g2718(n340 ,n2482 ,n2478);
    xnor g2719(n339 ,n2480 ,n2476);
    xnor g2720(n338 ,n2481 ,n2477);
    or g2721(n337 ,n319 ,n270);
    or g2722(n336 ,n301 ,n272);
    nor g2723(n335 ,n274 ,n293);
    or g2724(n334 ,n304 ,n302);
    nor g2725(n333 ,n2481 ,n2477);
    nor g2726(n332 ,n2480 ,n2476);
    nor g2727(n331 ,n2482 ,n2478);
    nor g2728(n330 ,n2479 ,n2475);
    not g2729(n329 ,n2513);
    not g2730(n328 ,n2504);
    not g2731(n327 ,n2540);
    not g2732(n326 ,n2522);
    not g2733(n325 ,n2516);
    not g2734(n324 ,n2490);
    not g2735(n323 ,n2499);
    not g2736(n322 ,n2510);
    not g2737(n321 ,n2539);
    not g2738(n320 ,n2523);
    not g2739(n319 ,n2530);
    not g2740(n318 ,n2500);
    not g2741(n317 ,n2487);
    not g2742(n316 ,n2497);
    not g2743(n315 ,n2485);
    not g2744(n314 ,n2488);
    not g2745(n313 ,n2519);
    not g2746(n312 ,n2505);
    not g2747(n311 ,n2518);
    not g2748(n310 ,n2520);
    not g2749(n309 ,n2491);
    not g2750(n308 ,n2517);
    not g2751(n307 ,n2506);
    not g2752(n306 ,n2493);
    not g2753(n305 ,n2502);
    not g2754(n304 ,n2532);
    not g2755(n303 ,n2535);
    not g2756(n302 ,n2531);
    not g2757(n301 ,n2528);
    not g2758(n300 ,n2533);
    not g2759(n299 ,n2537);
    not g2760(n298 ,n2486);
    not g2761(n297 ,n2525);
    not g2762(n296 ,n2483);
    not g2763(n295 ,n2521);
    not g2764(n294 ,n2492);
    not g2765(n293 ,n2475);
    not g2766(n292 ,n2494);
    not g2767(n291 ,n2496);
    not g2768(n290 ,n2524);
    not g2769(n289 ,n2498);
    not g2770(n288 ,n2495);
    not g2771(n287 ,n2501);
    not g2772(n286 ,n2536);
    not g2773(n285 ,n2512);
    not g2774(n284 ,n2507);
    not g2775(n283 ,n2509);
    not g2776(n282 ,n2489);
    not g2777(n281 ,n2484);
    not g2778(n280 ,n2508);
    not g2779(n279 ,n2541);
    not g2780(n278 ,n2514);
    not g2781(n277 ,n2511);
    not g2782(n276 ,n2503);
    not g2783(n275 ,n2515);
    not g2784(n274 ,n2479);
    not g2785(n273 ,n2538);
    not g2786(n272 ,n2527);
    not g2787(n271 ,n2534);
    not g2788(n270 ,n2529);
    not g2789(n269 ,n2526);
    xor g2790(n2607 ,n8[3] ,n527);
    nor g2791(n2608 ,n526 ,n527);
    nor g2792(n527 ,n522 ,n525);
    nor g2793(n526 ,n8[2] ,n524);
    nor g2794(n2609 ,n524 ,n523);
    not g2795(n525 ,n524);
    nor g2796(n524 ,n520 ,n521);
    nor g2797(n523 ,n8[1] ,n8[0]);
    not g2798(n522 ,n8[2]);
    not g2799(n521 ,n8[0]);
    not g2800(n520 ,n8[1]);
    xor g2801(n2410 ,n4[63] ,n2747);
    xor g2802(n2409 ,n4[62] ,n2745);
    nor g2803(n2747 ,n4[62] ,n2746);
    xor g2804(n2408 ,n4[61] ,n2743);
    not g2805(n2746 ,n2745);
    nor g2806(n2745 ,n4[61] ,n2744);
    xor g2807(n2407 ,n4[60] ,n2741);
    not g2808(n2744 ,n2743);
    nor g2809(n2743 ,n4[60] ,n2742);
    xor g2810(n2406 ,n4[59] ,n2739);
    not g2811(n2742 ,n2741);
    nor g2812(n2741 ,n4[59] ,n2740);
    xor g2813(n2405 ,n4[58] ,n2737);
    not g2814(n2740 ,n2739);
    nor g2815(n2739 ,n4[58] ,n2738);
    xor g2816(n2404 ,n4[57] ,n2735);
    not g2817(n2738 ,n2737);
    nor g2818(n2737 ,n4[57] ,n2736);
    xor g2819(n2403 ,n4[56] ,n2733);
    not g2820(n2736 ,n2735);
    nor g2821(n2735 ,n4[56] ,n2734);
    xor g2822(n2402 ,n4[55] ,n2731);
    not g2823(n2734 ,n2733);
    nor g2824(n2733 ,n4[55] ,n2732);
    xor g2825(n2401 ,n4[54] ,n2729);
    not g2826(n2732 ,n2731);
    nor g2827(n2731 ,n4[54] ,n2730);
    xor g2828(n2400 ,n4[53] ,n2727);
    not g2829(n2730 ,n2729);
    nor g2830(n2729 ,n4[53] ,n2728);
    xor g2831(n2399 ,n4[52] ,n2725);
    not g2832(n2728 ,n2727);
    nor g2833(n2727 ,n4[52] ,n2726);
    xor g2834(n2398 ,n4[51] ,n2723);
    not g2835(n2726 ,n2725);
    nor g2836(n2725 ,n4[51] ,n2724);
    xor g2837(n2397 ,n4[50] ,n2721);
    not g2838(n2724 ,n2723);
    nor g2839(n2723 ,n4[50] ,n2722);
    xor g2840(n2396 ,n4[49] ,n2719);
    not g2841(n2722 ,n2721);
    nor g2842(n2721 ,n4[49] ,n2720);
    xor g2843(n2395 ,n4[48] ,n2717);
    not g2844(n2720 ,n2719);
    nor g2845(n2719 ,n4[48] ,n2718);
    xor g2846(n2394 ,n4[47] ,n2715);
    not g2847(n2718 ,n2717);
    nor g2848(n2717 ,n4[47] ,n2716);
    xor g2849(n2393 ,n4[46] ,n2713);
    not g2850(n2716 ,n2715);
    nor g2851(n2715 ,n4[46] ,n2714);
    xor g2852(n2392 ,n4[45] ,n2711);
    not g2853(n2714 ,n2713);
    nor g2854(n2713 ,n4[45] ,n2712);
    xor g2855(n2391 ,n4[44] ,n2709);
    not g2856(n2712 ,n2711);
    nor g2857(n2711 ,n4[44] ,n2710);
    xor g2858(n2390 ,n4[43] ,n2707);
    not g2859(n2710 ,n2709);
    nor g2860(n2709 ,n4[43] ,n2708);
    xor g2861(n2389 ,n4[42] ,n2705);
    not g2862(n2708 ,n2707);
    nor g2863(n2707 ,n4[42] ,n2706);
    xor g2864(n2388 ,n4[41] ,n2703);
    not g2865(n2706 ,n2705);
    nor g2866(n2705 ,n4[41] ,n2704);
    xor g2867(n2387 ,n4[40] ,n2701);
    not g2868(n2704 ,n2703);
    nor g2869(n2703 ,n4[40] ,n2702);
    xor g2870(n2386 ,n4[39] ,n2699);
    not g2871(n2702 ,n2701);
    nor g2872(n2701 ,n4[39] ,n2700);
    xor g2873(n2385 ,n4[38] ,n2697);
    not g2874(n2700 ,n2699);
    nor g2875(n2699 ,n4[38] ,n2698);
    xor g2876(n2384 ,n4[37] ,n2695);
    not g2877(n2698 ,n2697);
    nor g2878(n2697 ,n4[37] ,n2696);
    xor g2879(n2383 ,n4[36] ,n2693);
    not g2880(n2696 ,n2695);
    nor g2881(n2695 ,n4[36] ,n2694);
    xor g2882(n2382 ,n4[35] ,n2691);
    not g2883(n2694 ,n2693);
    nor g2884(n2693 ,n4[35] ,n2692);
    xor g2885(n2381 ,n4[34] ,n2689);
    not g2886(n2692 ,n2691);
    nor g2887(n2691 ,n4[34] ,n2690);
    xor g2888(n2380 ,n4[33] ,n2687);
    not g2889(n2690 ,n2689);
    nor g2890(n2689 ,n4[33] ,n2688);
    xor g2891(n2379 ,n4[32] ,n2685);
    not g2892(n2688 ,n2687);
    nor g2893(n2687 ,n4[32] ,n2686);
    xor g2894(n2378 ,n4[31] ,n2683);
    not g2895(n2686 ,n2685);
    nor g2896(n2685 ,n4[31] ,n2684);
    xor g2897(n2377 ,n4[30] ,n2681);
    not g2898(n2684 ,n2683);
    nor g2899(n2683 ,n4[30] ,n2682);
    xor g2900(n2376 ,n4[29] ,n2679);
    not g2901(n2682 ,n2681);
    nor g2902(n2681 ,n4[29] ,n2680);
    xor g2903(n2375 ,n4[28] ,n2677);
    not g2904(n2680 ,n2679);
    nor g2905(n2679 ,n4[28] ,n2678);
    xor g2906(n2374 ,n4[27] ,n2675);
    not g2907(n2678 ,n2677);
    nor g2908(n2677 ,n4[27] ,n2676);
    xor g2909(n2373 ,n4[26] ,n2673);
    not g2910(n2676 ,n2675);
    nor g2911(n2675 ,n4[26] ,n2674);
    xor g2912(n2372 ,n4[25] ,n2671);
    not g2913(n2674 ,n2673);
    nor g2914(n2673 ,n4[25] ,n2672);
    xor g2915(n2371 ,n4[24] ,n2669);
    not g2916(n2672 ,n2671);
    nor g2917(n2671 ,n4[24] ,n2670);
    xor g2918(n2370 ,n4[23] ,n2667);
    not g2919(n2670 ,n2669);
    nor g2920(n2669 ,n4[23] ,n2668);
    xor g2921(n2369 ,n4[22] ,n2665);
    not g2922(n2668 ,n2667);
    nor g2923(n2667 ,n4[22] ,n2666);
    xor g2924(n2368 ,n4[21] ,n2663);
    not g2925(n2666 ,n2665);
    nor g2926(n2665 ,n4[21] ,n2664);
    xor g2927(n2367 ,n4[20] ,n2661);
    not g2928(n2664 ,n2663);
    nor g2929(n2663 ,n4[20] ,n2662);
    xor g2930(n2366 ,n4[19] ,n2659);
    not g2931(n2662 ,n2661);
    nor g2932(n2661 ,n4[19] ,n2660);
    xor g2933(n2365 ,n4[18] ,n2657);
    not g2934(n2660 ,n2659);
    nor g2935(n2659 ,n4[18] ,n2658);
    xor g2936(n2364 ,n4[17] ,n2655);
    not g2937(n2658 ,n2657);
    nor g2938(n2657 ,n4[17] ,n2656);
    xor g2939(n2363 ,n4[16] ,n2653);
    not g2940(n2656 ,n2655);
    nor g2941(n2655 ,n4[16] ,n2654);
    xor g2942(n2362 ,n4[15] ,n2651);
    not g2943(n2654 ,n2653);
    nor g2944(n2653 ,n4[15] ,n2652);
    xor g2945(n2361 ,n4[14] ,n2649);
    not g2946(n2652 ,n2651);
    nor g2947(n2651 ,n4[14] ,n2650);
    xor g2948(n2360 ,n4[13] ,n2647);
    not g2949(n2650 ,n2649);
    nor g2950(n2649 ,n4[13] ,n2648);
    xor g2951(n2359 ,n4[12] ,n2645);
    not g2952(n2648 ,n2647);
    nor g2953(n2647 ,n4[12] ,n2646);
    xor g2954(n2358 ,n4[11] ,n2643);
    not g2955(n2646 ,n2645);
    nor g2956(n2645 ,n4[11] ,n2644);
    xor g2957(n2357 ,n4[10] ,n2641);
    not g2958(n2644 ,n2643);
    nor g2959(n2643 ,n4[10] ,n2642);
    xor g2960(n2356 ,n4[9] ,n2639);
    not g2961(n2642 ,n2641);
    nor g2962(n2641 ,n4[9] ,n2640);
    xor g2963(n2355 ,n4[8] ,n2637);
    not g2964(n2640 ,n2639);
    nor g2965(n2639 ,n4[8] ,n2638);
    xor g2966(n2354 ,n4[7] ,n2635);
    not g2967(n2638 ,n2637);
    nor g2968(n2637 ,n4[7] ,n2636);
    xor g2969(n2353 ,n4[6] ,n2633);
    not g2970(n2636 ,n2635);
    nor g2971(n2635 ,n4[6] ,n2634);
    xor g2972(n2352 ,n4[5] ,n2631);
    not g2973(n2634 ,n2633);
    nor g2974(n2633 ,n4[5] ,n2632);
    xnor g2975(n2351 ,n4[4] ,n2630);
    not g2976(n2632 ,n2631);
    nor g2977(n2631 ,n4[4] ,n2630);
    nor g2978(n2630 ,n2614 ,n2629);
    xor g2979(n2350 ,n2628 ,n2619);
    nor g2980(n2629 ,n2620 ,n2628);
    nor g2981(n2628 ,n2615 ,n2627);
    xor g2982(n2349 ,n2626 ,n2621);
    nor g2983(n2627 ,n2622 ,n2626);
    nor g2984(n2626 ,n2618 ,n2625);
    xnor g2985(n2348 ,n2623 ,n2616);
    nor g2986(n2625 ,n2617 ,n2624);
    not g2987(n2624 ,n2623);
    xnor g2988(n2623 ,n6[1] ,n4[1]);
    not g2989(n2622 ,n2621);
    xnor g2990(n2621 ,n6[2] ,n4[2]);
    xor g2991(n2347 ,n6[0] ,n4[0]);
    not g2992(n2620 ,n2619);
    xnor g2993(n2619 ,n6[3] ,n4[3]);
    nor g2994(n2618 ,n2612 ,n4[1]);
    not g2995(n2617 ,n2616);
    nor g2996(n2616 ,n2613 ,n4[0]);
    nor g2997(n2615 ,n2611 ,n4[2]);
    nor g2998(n2614 ,n2610 ,n4[3]);
    not g2999(n2613 ,n6[0]);
    not g3000(n2612 ,n6[1]);
    not g3001(n2611 ,n6[2]);
    not g3002(n2610 ,n6[3]);
    xnor g3003(n6[3] ,n2842 ,n10[31]);
    xnor g3004(n6[2] ,n2842 ,n10[30]);
    xnor g3005(n6[1] ,n2842 ,n10[29]);
    xnor g3006(n6[0] ,n2842 ,n10[28]);
    or g3007(n2842 ,n2840 ,n2841);
    or g3008(n2841 ,n2839 ,n2836);
    or g3009(n2840 ,n2837 ,n2838);
    or g3010(n2839 ,n2833 ,n2835);
    or g3011(n2838 ,n2834 ,n2829);
    or g3012(n2837 ,n2831 ,n2832);
    or g3013(n2836 ,n2830 ,n2828);
    or g3014(n2835 ,n2827 ,n2820);
    or g3015(n2834 ,n2825 ,n2821);
    or g3016(n2833 ,n2826 ,n2824);
    or g3017(n2832 ,n2822 ,n2814);
    or g3018(n2831 ,n2823 ,n2819);
    or g3019(n2830 ,n2815 ,n2817);
    or g3020(n2829 ,n2818 ,n2813);
    or g3021(n2828 ,n2816 ,n2812);
    or g3022(n2827 ,n2798 ,n2797);
    or g3023(n2826 ,n2810 ,n2809);
    or g3024(n2825 ,n2808 ,n2799);
    or g3025(n2824 ,n2802 ,n2801);
    or g3026(n2823 ,n2796 ,n2794);
    or g3027(n2822 ,n2807 ,n2791);
    or g3028(n2821 ,n2780 ,n2793);
    or g3029(n2820 ,n2786 ,n2782);
    or g3030(n2819 ,n2804 ,n2803);
    or g3031(n2818 ,n2789 ,n2795);
    or g3032(n2817 ,n2806 ,n2781);
    or g3033(n2816 ,n2788 ,n2787);
    or g3034(n2815 ,n2792 ,n2790);
    or g3035(n2814 ,n2805 ,n2783);
    or g3036(n2813 ,n2800 ,n2784);
    or g3037(n2812 ,n2811 ,n2785);
    or g3038(n2811 ,n2757 ,n9[8]);
    or g3039(n2810 ,n2754 ,n2748);
    or g3040(n2809 ,n2750 ,n2756);
    or g3041(n2808 ,n2753 ,n2760);
    or g3042(n2807 ,n2769 ,n2777);
    or g3043(n2806 ,n2765 ,n2758);
    or g3044(n2805 ,n2749 ,n2779);
    or g3045(n2804 ,n2764 ,n9[23]);
    or g3046(n2803 ,n2767 ,n9[21]);
    or g3047(n2802 ,n2755 ,n11[26]);
    or g3048(n2801 ,n2761 ,n11[24]);
    or g3049(n2800 ,n2778 ,n9[29]);
    or g3050(n2799 ,n2770 ,n9[24]);
    or g3051(n2798 ,n2752 ,n11[18]);
    or g3052(n2797 ,n2751 ,n11[16]);
    or g3053(n2796 ,n2768 ,n2771);
    or g3054(n2795 ,n11[31] ,n11[30]);
    or g3055(n2794 ,n2774 ,n11[14]);
    or g3056(n2793 ,n2766 ,n9[17]);
    or g3057(n2792 ,n2763 ,n9[6]);
    or g3058(n2791 ,n2775 ,n11[4]);
    or g3059(n2790 ,n2776 ,n9[4]);
    or g3060(n2789 ,n2759 ,n11[28]);
    or g3061(n2788 ,n2773 ,n9[15]);
    or g3062(n2787 ,n2772 ,n9[13]);
    or g3063(n2786 ,n11[3] ,n11[2]);
    or g3064(n2785 ,n9[11] ,n9[10]);
    or g3065(n2784 ,n9[31] ,n9[30]);
    or g3066(n2783 ,n11[9] ,n11[8]);
    or g3067(n2782 ,n11[1] ,n11[0]);
    or g3068(n2781 ,n9[1] ,n9[0]);
    or g3069(n2780 ,n2762 ,n9[19]);
    not g3070(n2779 ,n11[10]);
    not g3071(n2778 ,n9[28]);
    not g3072(n2777 ,n11[6]);
    not g3073(n2776 ,n9[5]);
    not g3074(n2775 ,n11[5]);
    not g3075(n2774 ,n11[15]);
    not g3076(n2773 ,n9[14]);
    not g3077(n2772 ,n9[12]);
    not g3078(n2771 ,n11[12]);
    not g3079(n2770 ,n9[25]);
    not g3080(n2769 ,n11[7]);
    not g3081(n2768 ,n11[13]);
    not g3082(n2767 ,n9[20]);
    not g3083(n2766 ,n9[16]);
    not g3084(n2765 ,n9[3]);
    not g3085(n2764 ,n9[22]);
    not g3086(n2763 ,n9[7]);
    not g3087(n2762 ,n9[18]);
    not g3088(n2761 ,n11[25]);
    not g3089(n2760 ,n9[26]);
    not g3090(n2759 ,n11[29]);
    not g3091(n2758 ,n9[2]);
    not g3092(n2757 ,n9[9]);
    not g3093(n2756 ,n11[20]);
    not g3094(n2755 ,n11[27]);
    not g3095(n2754 ,n11[23]);
    not g3096(n2753 ,n9[27]);
    not g3097(n2752 ,n11[19]);
    not g3098(n2751 ,n11[17]);
    not g3099(n2750 ,n11[21]);
    not g3100(n2749 ,n11[11]);
    not g3101(n2748 ,n11[22]);
endmodule
