module top(n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [3:0] n6;
    wire [31:0] n7;
    wire [31:0] n8;
    wire [1:0] n9;
    wire [31:0] n10;
    wire n11, n12, n13, n14, n15, n16, n17, n18;
    wire n19, n20, n21, n22, n23, n24, n25, n26;
    wire n27, n28, n29, n30, n31, n32, n33, n34;
    wire n35, n36, n37, n38, n39, n40, n41, n42;
    wire n43, n44, n45, n46, n47, n48, n49, n50;
    wire n51, n52, n53, n54, n55, n56, n57, n58;
    wire n59, n60, n61, n62, n63, n64, n65, n66;
    wire n67, n68, n69, n70, n71, n72, n73, n74;
    wire n75, n76, n77, n78, n79, n80, n81, n82;
    wire n83, n84, n85, n86, n87, n88, n89, n90;
    wire n91, n92, n93, n94, n95, n96, n97, n98;
    wire n99, n100, n101, n102, n103, n104, n105, n106;
    wire n107, n108, n109, n110, n111, n112, n113, n114;
    wire n115, n116, n117, n118, n119, n120, n121, n122;
    wire n123, n124, n125, n126, n127, n128, n129, n130;
    wire n131, n132, n133, n134, n135, n136, n137, n138;
    wire n139, n140, n141, n142, n143, n144, n145, n146;
    wire n147, n148, n149, n150, n151, n152, n153, n154;
    wire n155, n156, n157, n158, n159, n160, n161, n162;
    wire n163, n164, n165, n166, n167, n168, n169, n170;
    wire n171, n172, n173, n174, n175, n176, n177, n178;
    wire n179, n180, n181, n182, n183, n184, n185, n186;
    wire n187, n188, n189, n190, n191, n192, n193, n194;
    wire n195, n196, n197, n198, n199, n200, n201, n202;
    wire n203, n204, n205, n206, n207, n208, n209, n210;
    wire n211, n212, n213, n214, n215, n216, n217, n218;
    wire n219, n220, n221, n222, n223, n224, n225, n226;
    wire n227, n228, n229, n230, n231, n232, n233, n234;
    wire n235, n236, n237, n238, n239, n240, n241, n242;
    wire n243, n244, n245, n246, n247, n248, n249, n250;
    wire n251, n252, n253, n254, n255, n256, n257, n258;
    wire n259, n260, n261, n262, n263, n264, n265, n266;
    wire n267, n268, n269, n270, n271, n272, n273, n274;
    wire n275, n276, n277, n278, n279, n280, n281, n282;
    wire n283, n284, n285, n286, n287, n288, n289, n290;
    wire n291, n292, n293, n294, n295, n296, n297, n298;
    wire n299, n300, n301, n302, n303, n304, n305, n306;
    wire n307, n308, n309, n310, n311, n312, n313, n314;
    wire n315, n316, n317, n318, n319, n320, n321, n322;
    wire n323, n324, n325, n326, n327, n328, n329, n330;
    wire n331, n332, n333, n334, n335, n336, n337, n338;
    wire n339, n340, n341, n342, n343, n344, n345, n346;
    wire n347, n348, n349, n350, n351, n352, n353, n354;
    wire n355, n356, n357, n358, n359, n360, n361, n362;
    wire n363, n364, n365, n366, n367, n368, n369, n370;
    wire n371, n372, n373, n374, n375, n376, n377, n378;
    wire n379, n380, n381, n382, n383, n384, n385, n386;
    wire n387, n388, n389, n390, n391, n392, n393, n394;
    wire n395, n396, n397, n398, n399, n400, n401, n402;
    wire n403, n404, n405, n406, n407, n408, n409, n410;
    wire n411, n412, n413, n414, n415, n416, n417, n418;
    wire n419, n420, n421, n422, n423, n424, n425, n426;
    wire n427, n428, n429, n430, n431, n432, n433, n434;
    wire n435, n436, n437, n438, n439, n440, n441, n442;
    wire n443, n444, n445, n446, n447, n448, n449, n450;
    wire n451, n452, n453, n454, n455, n456, n457, n458;
    wire n459, n460, n461, n462, n463, n464, n465, n466;
    wire n467, n468, n469, n470, n471, n472, n473, n474;
    wire n475, n476, n477, n478, n479, n480, n481, n482;
    wire n483, n484, n485, n486, n487, n488, n489, n490;
    wire n491, n492, n493, n494, n495, n496, n497, n498;
    wire n499, n500, n501, n502, n503, n504, n505, n506;
    wire n507, n508, n509, n510, n511, n512, n513, n514;
    wire n515, n516, n517, n518, n519, n520, n521, n522;
    wire n523, n524, n525, n526, n527, n528, n529, n530;
    wire n531, n532, n533, n534, n535, n536, n537, n538;
    wire n539, n540, n541, n542, n543, n544, n545, n546;
    wire n547, n548, n549, n550, n551, n552, n553, n554;
    wire n555, n556, n557, n558, n559, n560, n561, n562;
    wire n563, n564, n565, n566, n567, n568, n569, n570;
    wire n571, n572, n573, n574, n575, n576, n577, n578;
    wire n579, n580, n581, n582, n583, n584, n585, n586;
    wire n587, n588, n589, n590, n591, n592, n593, n594;
    wire n595, n596, n597, n598, n599, n600, n601, n602;
    wire n603, n604, n605, n606, n607, n608, n609, n610;
    wire n611, n612, n613, n614, n615, n616, n617, n618;
    wire n619, n620, n621, n622, n623, n624, n625, n626;
    wire n627, n628, n629, n630, n631, n632, n633, n634;
    wire n635, n636, n637, n638, n639, n640, n641, n642;
    wire n643, n644, n645, n646, n647, n648, n649, n650;
    wire n651, n652, n653, n654, n655, n656, n657, n658;
    wire n659, n660, n661, n662, n663, n664, n665, n666;
    wire n667, n668, n669, n670, n671, n672, n673, n674;
    wire n675, n676, n677, n678, n679, n680, n681, n682;
    wire n683, n684, n685, n686, n687, n688, n689, n690;
    wire n691, n692, n693, n694, n695, n696, n697, n698;
    wire n699, n700, n701, n702, n703, n704, n705, n706;
    wire n707, n708, n709, n710, n711, n712, n713, n714;
    wire n715, n716, n717, n718, n719, n720, n721, n722;
    wire n723, n724, n725, n726, n727, n728, n729, n730;
    wire n731, n732, n733, n734, n735, n736, n737, n738;
    wire n739, n740, n741, n742, n743, n744, n745, n746;
    wire n747, n748, n749, n750, n751, n752, n753, n754;
    wire n755, n756, n757, n758, n759, n760, n761, n762;
    wire n763, n764, n765, n766, n767, n768, n769, n770;
    wire n771, n772, n773, n774, n775, n776, n777, n778;
    wire n779, n780, n781, n782, n783, n784, n785, n786;
    wire n787, n788, n789, n790, n791, n792, n793, n794;
    wire n795, n796, n797, n798, n799, n800, n801, n802;
    wire n803, n804, n805, n806, n807, n808, n809, n810;
    wire n811, n812, n813, n814, n815, n816, n817, n818;
    wire n819, n820, n821, n822, n823, n824, n825, n826;
    wire n827, n828, n829, n830, n831, n832, n833, n834;
    wire n835, n836, n837, n838, n839, n840, n841, n842;
    wire n843, n844, n845, n846, n847, n848, n849, n850;
    wire n851, n852, n853, n854, n855, n856, n857, n858;
    wire n859, n860, n861, n862, n863, n864, n865, n866;
    wire n867, n868, n869, n870, n871, n872, n873, n874;
    wire n875, n876, n877, n878, n879, n880, n881, n882;
    wire n883, n884, n885, n886, n887, n888, n889, n890;
    wire n891, n892, n893, n894, n895, n896, n897, n898;
    wire n899, n900, n901, n902, n903, n904, n905, n906;
    wire n907, n908, n909, n910, n911, n912, n913, n914;
    wire n915, n916, n917, n918, n919, n920, n921, n922;
    wire n923, n924, n925, n926, n927, n928, n929, n930;
    wire n931, n932, n933, n934, n935, n936, n937, n938;
    wire n939, n940, n941, n942, n943, n944, n945, n946;
    wire n947, n948, n949, n950, n951, n952, n953, n954;
    wire n955, n956, n957, n958, n959, n960, n961, n962;
    wire n963, n964, n965, n966, n967, n968, n969, n970;
    wire n971, n972, n973, n974, n975, n976, n977, n978;
    wire n979, n980, n981, n982, n983, n984, n985, n986;
    wire n987, n988, n989, n990, n991, n992, n993, n994;
    wire n995, n996, n997, n998, n999, n1000, n1001, n1002;
    wire n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010;
    wire n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
    wire n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
    wire n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
    wire n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
    wire n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050;
    wire n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058;
    wire n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066;
    wire n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074;
    wire n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082;
    wire n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090;
    wire n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098;
    wire n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106;
    wire n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114;
    wire n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122;
    wire n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130;
    wire n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138;
    wire n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146;
    wire n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154;
    wire n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162;
    wire n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170;
    wire n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178;
    wire n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186;
    wire n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194;
    wire n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202;
    wire n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210;
    wire n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218;
    wire n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226;
    wire n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234;
    wire n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242;
    wire n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250;
    wire n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258;
    wire n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266;
    wire n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274;
    wire n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282;
    wire n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
    wire n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298;
    wire n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306;
    wire n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314;
    wire n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322;
    wire n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330;
    wire n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338;
    wire n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346;
    wire n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;
    wire n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;
    wire n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370;
    wire n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378;
    wire n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386;
    wire n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394;
    wire n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402;
    wire n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410;
    wire n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418;
    wire n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426;
    wire n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434;
    wire n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442;
    wire n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450;
    wire n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458;
    wire n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466;
    wire n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474;
    wire n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482;
    wire n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490;
    wire n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498;
    wire n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506;
    wire n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514;
    wire n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522;
    wire n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530;
    wire n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538;
    wire n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546;
    wire n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554;
    wire n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562;
    wire n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570;
    wire n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578;
    wire n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586;
    wire n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594;
    wire n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602;
    wire n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610;
    wire n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618;
    wire n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626;
    wire n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634;
    wire n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642;
    wire n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650;
    wire n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658;
    wire n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666;
    wire n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674;
    wire n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682;
    wire n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690;
    wire n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698;
    wire n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706;
    wire n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714;
    wire n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722;
    wire n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730;
    wire n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738;
    wire n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746;
    wire n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754;
    wire n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762;
    wire n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770;
    wire n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778;
    wire n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786;
    wire n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794;
    wire n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802;
    wire n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810;
    wire n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818;
    wire n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826;
    wire n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834;
    wire n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842;
    wire n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850;
    wire n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858;
    wire n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866;
    wire n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874;
    wire n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882;
    wire n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
    wire n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898;
    wire n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906;
    wire n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914;
    wire n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922;
    wire n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930;
    wire n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938;
    wire n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946;
    wire n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954;
    wire n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962;
    wire n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970;
    wire n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978;
    wire n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986;
    wire n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994;
    wire n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002;
    wire n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010;
    wire n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018;
    wire n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026;
    wire n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034;
    wire n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042;
    wire n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050;
    wire n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058;
    wire n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066;
    wire n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074;
    wire n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082;
    wire n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090;
    wire n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098;
    wire n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106;
    wire n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114;
    wire n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122;
    wire n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130;
    wire n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138;
    wire n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146;
    wire n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154;
    wire n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162;
    wire n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170;
    wire n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178;
    wire n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186;
    wire n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194;
    wire n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202;
    wire n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210;
    wire n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218;
    wire n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226;
    wire n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234;
    wire n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242;
    wire n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250;
    wire n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258;
    wire n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266;
    wire n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274;
    wire n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282;
    wire n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290;
    wire n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298;
    wire n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306;
    wire n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314;
    wire n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322;
    wire n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330;
    wire n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338;
    wire n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346;
    wire n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354;
    wire n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362;
    wire n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370;
    wire n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378;
    wire n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386;
    wire n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394;
    wire n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402;
    wire n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410;
    wire n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418;
    wire n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426;
    wire n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434;
    wire n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442;
    wire n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450;
    wire n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458;
    wire n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466;
    wire n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474;
    wire n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482;
    wire n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490;
    wire n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498;
    wire n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506;
    wire n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514;
    wire n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522;
    wire n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530;
    wire n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538;
    wire n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546;
    wire n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554;
    wire n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562;
    wire n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570;
    wire n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578;
    wire n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586;
    wire n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594;
    wire n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602;
    wire n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610;
    wire n2611, n2612, n2613, n2614, n2615, n2616;
    not g0(n2505 ,n1);
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2397), .Q(n5[0]));
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2420), .Q(n5[1]));
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2408), .Q(n5[2]));
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2393), .Q(n5[3]));
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2389), .Q(n5[4]));
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2382), .Q(n5[5]));
    dff g7(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2479), .Q(n5[6]));
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2488), .Q(n5[7]));
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2475), .Q(n5[8]));
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2471), .Q(n5[9]));
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2463), .Q(n5[10]));
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2449), .Q(n5[11]));
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2450), .Q(n5[12]));
    dff g14(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2448), .Q(n5[13]));
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2447), .Q(n5[14]));
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2446), .Q(n5[15]));
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2445), .Q(n5[16]));
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2444), .Q(n5[17]));
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2443), .Q(n5[18]));
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2442), .Q(n5[19]));
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2441), .Q(n5[20]));
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2440), .Q(n5[21]));
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2439), .Q(n5[22]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2438), .Q(n5[23]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2437), .Q(n5[24]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2436), .Q(n5[25]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2435), .Q(n5[26]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2434), .Q(n5[27]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2433), .Q(n5[28]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2432), .Q(n5[29]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2430), .Q(n5[30]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2431), .Q(n5[31]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2429), .Q(n5[32]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2428), .Q(n5[33]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2427), .Q(n5[34]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2426), .Q(n5[35]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2423), .Q(n5[36]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2418), .Q(n5[37]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2414), .Q(n5[38]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2413), .Q(n5[39]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2411), .Q(n5[40]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2407), .Q(n5[41]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2404), .Q(n5[42]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2401), .Q(n5[43]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2399), .Q(n5[44]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2395), .Q(n5[45]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2391), .Q(n5[46]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2387), .Q(n5[47]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2384), .Q(n5[48]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2381), .Q(n5[49]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2377), .Q(n5[50]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2501), .Q(n5[51]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2499), .Q(n5[52]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2497), .Q(n5[53]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2492), .Q(n5[54]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2490), .Q(n5[55]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2487), .Q(n5[56]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2485), .Q(n5[57]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2482), .Q(n5[58]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2477), .Q(n5[59]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2473), .Q(n5[60]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2469), .Q(n5[61]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2466), .Q(n5[62]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2462), .Q(n5[63]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n760), .Q(n6[0]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n960), .Q(n6[1]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n961), .Q(n6[2]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n965), .Q(n6[3]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2375), .Q(n3[0]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2328), .Q(n3[1]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2374), .Q(n3[2]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2373), .Q(n3[3]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2372), .Q(n3[4]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2371), .Q(n3[5]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2370), .Q(n3[6]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2369), .Q(n3[7]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2368), .Q(n3[8]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2367), .Q(n3[9]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2366), .Q(n3[10]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2365), .Q(n3[11]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2364), .Q(n3[12]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2363), .Q(n3[13]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2362), .Q(n3[14]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2361), .Q(n3[15]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2360), .Q(n3[16]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2359), .Q(n3[17]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2358), .Q(n3[18]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2357), .Q(n3[19]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2356), .Q(n3[20]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2355), .Q(n3[21]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2354), .Q(n3[22]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2353), .Q(n3[23]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2352), .Q(n3[24]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2351), .Q(n3[25]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2350), .Q(n3[26]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2349), .Q(n3[27]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2348), .Q(n3[28]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2347), .Q(n3[29]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2346), .Q(n3[30]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2345), .Q(n3[31]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2344), .Q(n3[32]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2343), .Q(n3[33]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2342), .Q(n3[34]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2341), .Q(n3[35]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2340), .Q(n3[36]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2339), .Q(n3[37]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2338), .Q(n3[38]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2337), .Q(n3[39]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2336), .Q(n3[40]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2335), .Q(n3[41]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2334), .Q(n3[42]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2333), .Q(n3[43]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2332), .Q(n3[44]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2331), .Q(n3[45]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2330), .Q(n3[46]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2329), .Q(n3[47]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2376), .Q(n3[48]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2327), .Q(n3[49]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2326), .Q(n3[50]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2325), .Q(n3[51]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2324), .Q(n3[52]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2323), .Q(n3[53]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2322), .Q(n3[54]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2321), .Q(n3[55]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2320), .Q(n3[56]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2319), .Q(n3[57]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2318), .Q(n3[58]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2317), .Q(n3[59]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2316), .Q(n3[60]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2315), .Q(n3[61]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2314), .Q(n3[62]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2313), .Q(n3[63]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2425), .Q(n4[0]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2472), .Q(n4[1]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2422), .Q(n4[2]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2421), .Q(n4[3]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2419), .Q(n4[4]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n4[5]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2416), .Q(n4[6]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2415), .Q(n4[7]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2412), .Q(n4[8]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2410), .Q(n4[9]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2409), .Q(n4[10]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2406), .Q(n4[11]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2405), .Q(n4[12]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2403), .Q(n4[13]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2402), .Q(n4[14]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2400), .Q(n4[15]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2398), .Q(n4[16]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2396), .Q(n4[17]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2394), .Q(n4[18]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2392), .Q(n4[19]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2390), .Q(n4[20]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2388), .Q(n4[21]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2386), .Q(n4[22]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2385), .Q(n4[23]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2383), .Q(n4[24]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2380), .Q(n4[25]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2379), .Q(n4[26]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2378), .Q(n4[27]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2503), .Q(n4[28]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2502), .Q(n4[29]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2500), .Q(n4[30]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2498), .Q(n4[31]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2496), .Q(n4[32]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2495), .Q(n4[33]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2494), .Q(n4[34]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2493), .Q(n4[35]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2491), .Q(n4[36]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2489), .Q(n4[37]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2504), .Q(n4[38]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2486), .Q(n4[39]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2484), .Q(n4[40]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2483), .Q(n4[41]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2481), .Q(n4[42]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2480), .Q(n4[43]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2478), .Q(n4[44]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2476), .Q(n4[45]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2474), .Q(n4[46]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2424), .Q(n4[47]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2470), .Q(n4[48]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2468), .Q(n4[49]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2467), .Q(n4[50]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2465), .Q(n4[51]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2464), .Q(n4[52]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2461), .Q(n4[53]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2460), .Q(n4[54]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2459), .Q(n4[55]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2458), .Q(n4[56]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2457), .Q(n4[57]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2456), .Q(n4[58]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2455), .Q(n4[59]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2454), .Q(n4[60]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2453), .Q(n4[61]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2452), .Q(n4[62]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2451), .Q(n4[63]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n934), .Q(n7[0]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n954), .Q(n7[1]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n923), .Q(n7[2]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n913), .Q(n7[3]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n926), .Q(n7[4]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n971), .Q(n7[5]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n943), .Q(n7[6]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n970), .Q(n7[7]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n908), .Q(n7[8]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n911), .Q(n7[9]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n949), .Q(n7[10]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n936), .Q(n7[11]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n969), .Q(n7[12]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n952), .Q(n7[13]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n953), .Q(n7[14]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n958), .Q(n7[15]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n920), .Q(n7[16]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n939), .Q(n7[17]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n973), .Q(n7[18]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n929), .Q(n7[19]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n937), .Q(n7[20]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n918), .Q(n7[21]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n917), .Q(n7[22]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n928), .Q(n7[23]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n916), .Q(n7[24]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n910), .Q(n7[25]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n921), .Q(n7[26]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n966), .Q(n7[27]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n946), .Q(n7[28]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n959), .Q(n7[29]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n962), .Q(n7[30]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n935), .Q(n7[31]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n933), .Q(n8[0]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n930), .Q(n8[1]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n827), .Q(n8[2]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n931), .Q(n8[3]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n957), .Q(n8[4]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n925), .Q(n8[5]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n938), .Q(n8[6]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n947), .Q(n8[7]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n948), .Q(n8[8]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n914), .Q(n8[9]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n951), .Q(n8[10]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n968), .Q(n8[11]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n912), .Q(n8[12]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n924), .Q(n8[13]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n972), .Q(n8[14]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n963), .Q(n8[15]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n945), .Q(n8[16]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n915), .Q(n8[17]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n955), .Q(n8[18]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1167), .Q(n8[19]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n922), .Q(n8[20]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n927), .Q(n8[21]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n919), .Q(n8[22]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n950), .Q(n8[23]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n974), .Q(n8[24]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n909), .Q(n8[25]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n944), .Q(n8[26]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n940), .Q(n8[27]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n964), .Q(n8[28]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n932), .Q(n8[29]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n956), .Q(n8[30]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n967), .Q(n8[31]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1232), .Q(n9[0]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1230), .Q(n9[1]));
    or g263(n2504 ,n2168 ,n2295);
    or g264(n2503 ,n2184 ,n2311);
    or g265(n2502 ,n2182 ,n2310);
    or g266(n2501 ,n2181 ,n2312);
    or g267(n2500 ,n2180 ,n2309);
    or g268(n2499 ,n2179 ,n2307);
    or g269(n2498 ,n2178 ,n2308);
    or g270(n2497 ,n2176 ,n2304);
    or g271(n2496 ,n2177 ,n2306);
    or g272(n2495 ,n2175 ,n2305);
    or g273(n2494 ,n2174 ,n2303);
    or g274(n2493 ,n2172 ,n2300);
    or g275(n2492 ,n2173 ,n2301);
    or g276(n2491 ,n2171 ,n2299);
    or g277(n2490 ,n2049 ,n2297);
    or g278(n2489 ,n2169 ,n2296);
    or g279(n2488 ,n2170 ,n2294);
    or g280(n2487 ,n2167 ,n2292);
    or g281(n2486 ,n2166 ,n2293);
    or g282(n2485 ,n2164 ,n2290);
    or g283(n2484 ,n2165 ,n2291);
    or g284(n2483 ,n2163 ,n2289);
    or g285(n2482 ,n2161 ,n2286);
    or g286(n2481 ,n2162 ,n2288);
    or g287(n2480 ,n2160 ,n2285);
    or g288(n2479 ,n2183 ,n2302);
    or g289(n2478 ,n2159 ,n2284);
    or g290(n2477 ,n1999 ,n2283);
    or g291(n2476 ,n2157 ,n2282);
    or g292(n2475 ,n2158 ,n2287);
    or g293(n2474 ,n2156 ,n2281);
    or g294(n2473 ,n2155 ,n2279);
    or g295(n2472 ,n2040 ,n2231);
    or g296(n2471 ,n2150 ,n2268);
    or g297(n2470 ,n2153 ,n2278);
    or g298(n2469 ,n2152 ,n2277);
    or g299(n2468 ,n2151 ,n2276);
    or g300(n2467 ,n2149 ,n2275);
    or g301(n2466 ,n2148 ,n2274);
    or g302(n2465 ,n2147 ,n2273);
    or g303(n2464 ,n2146 ,n2272);
    or g304(n2463 ,n2142 ,n2265);
    or g305(n2462 ,n2144 ,n2271);
    or g306(n2461 ,n2145 ,n2270);
    or g307(n2460 ,n2143 ,n2269);
    or g308(n2459 ,n2141 ,n2267);
    or g309(n2458 ,n2139 ,n2266);
    or g310(n2457 ,n2138 ,n2264);
    or g311(n2456 ,n2137 ,n2263);
    or g312(n2455 ,n2136 ,n2262);
    or g313(n2454 ,n2061 ,n2260);
    or g314(n2453 ,n2134 ,n2259);
    or g315(n2452 ,n2132 ,n2258);
    or g316(n2451 ,n2130 ,n2257);
    or g317(n2450 ,n2128 ,n2256);
    or g318(n2449 ,n2133 ,n2261);
    or g319(n2448 ,n2125 ,n2255);
    or g320(n2447 ,n2120 ,n2254);
    or g321(n2446 ,n2117 ,n2252);
    or g322(n2445 ,n2114 ,n2253);
    or g323(n2444 ,n2109 ,n2251);
    or g324(n2443 ,n2107 ,n2250);
    or g325(n2442 ,n2103 ,n2249);
    or g326(n2441 ,n2099 ,n2248);
    or g327(n2440 ,n2096 ,n2247);
    or g328(n2439 ,n2092 ,n2246);
    or g329(n2438 ,n2089 ,n2245);
    or g330(n2437 ,n2085 ,n2244);
    or g331(n2436 ,n2078 ,n2243);
    or g332(n2435 ,n2076 ,n2242);
    or g333(n2434 ,n2072 ,n2241);
    or g334(n2433 ,n2069 ,n2240);
    or g335(n2432 ,n2064 ,n2239);
    or g336(n2431 ,n2055 ,n2237);
    or g337(n2430 ,n2056 ,n2238);
    or g338(n2429 ,n2051 ,n2236);
    or g339(n2428 ,n2047 ,n2235);
    or g340(n2427 ,n2044 ,n2234);
    or g341(n2426 ,n2041 ,n2233);
    or g342(n2425 ,n2042 ,n2280);
    or g343(n2424 ,n2154 ,n2232);
    or g344(n2423 ,n2039 ,n2227);
    or g345(n2422 ,n2038 ,n2230);
    or g346(n2421 ,n2037 ,n2228);
    or g347(n2420 ,n2033 ,n2229);
    or g348(n2419 ,n2036 ,n2226);
    or g349(n2418 ,n2035 ,n2225);
    or g350(n2417 ,n2034 ,n2224);
    or g351(n2416 ,n2031 ,n2222);
    or g352(n2415 ,n2030 ,n2221);
    or g353(n2414 ,n2032 ,n2223);
    or g354(n2413 ,n2029 ,n2220);
    or g355(n2412 ,n2028 ,n2219);
    or g356(n2411 ,n2026 ,n2216);
    or g357(n2410 ,n2027 ,n2217);
    or g358(n2409 ,n2025 ,n2215);
    or g359(n2408 ,n2024 ,n2211);
    or g360(n2407 ,n2022 ,n2213);
    or g361(n2406 ,n2023 ,n2214);
    or g362(n2405 ,n2021 ,n2212);
    or g363(n2404 ,n2020 ,n2210);
    or g364(n2403 ,n2019 ,n2209);
    or g365(n2402 ,n2018 ,n2208);
    or g366(n2401 ,n2017 ,n2207);
    or g367(n2400 ,n2016 ,n2206);
    or g368(n2399 ,n2014 ,n2202);
    or g369(n2398 ,n2015 ,n2204);
    or g370(n2397 ,n2080 ,n2218);
    or g371(n2396 ,n2012 ,n2203);
    or g372(n2395 ,n2010 ,n2199);
    or g373(n2394 ,n2011 ,n2201);
    or g374(n2393 ,n2013 ,n2205);
    or g375(n2392 ,n2009 ,n2200);
    or g376(n2391 ,n2008 ,n2197);
    or g377(n2390 ,n2007 ,n2198);
    or g378(n2389 ,n2006 ,n2190);
    or g379(n2388 ,n2005 ,n2196);
    or g380(n2387 ,n2004 ,n2195);
    or g381(n2386 ,n2003 ,n2194);
    or g382(n2385 ,n2002 ,n2193);
    or g383(n2384 ,n2001 ,n2192);
    or g384(n2383 ,n2000 ,n2191);
    or g385(n2382 ,n1995 ,n2298);
    or g386(n2381 ,n1997 ,n2188);
    or g387(n2380 ,n1998 ,n2189);
    or g388(n2379 ,n1996 ,n2187);
    or g389(n2378 ,n1994 ,n2186);
    or g390(n2377 ,n1993 ,n2185);
    or g391(n2376 ,n2066 ,n1816);
    or g392(n2375 ,n2140 ,n1864);
    or g393(n2374 ,n2131 ,n1862);
    or g394(n2373 ,n2129 ,n1861);
    or g395(n2372 ,n2127 ,n1860);
    or g396(n2371 ,n2126 ,n1859);
    or g397(n2370 ,n2124 ,n1858);
    or g398(n2369 ,n2123 ,n1857);
    or g399(n2368 ,n2122 ,n1856);
    or g400(n2367 ,n2121 ,n1855);
    or g401(n2366 ,n2119 ,n1854);
    or g402(n2365 ,n2118 ,n1853);
    or g403(n2364 ,n2116 ,n1852);
    or g404(n2363 ,n2115 ,n1851);
    or g405(n2362 ,n2113 ,n1850);
    or g406(n2361 ,n2112 ,n1849);
    or g407(n2360 ,n2111 ,n1848);
    or g408(n2359 ,n2110 ,n1847);
    or g409(n2358 ,n2108 ,n1846);
    or g410(n2357 ,n2106 ,n1845);
    or g411(n2356 ,n2105 ,n1844);
    or g412(n2355 ,n2104 ,n1843);
    or g413(n2354 ,n2102 ,n1842);
    or g414(n2353 ,n2101 ,n1841);
    or g415(n2352 ,n2100 ,n1840);
    or g416(n2351 ,n2098 ,n1839);
    or g417(n2350 ,n2097 ,n1838);
    or g418(n2349 ,n2095 ,n1837);
    or g419(n2348 ,n2094 ,n1836);
    or g420(n2347 ,n2093 ,n1835);
    or g421(n2346 ,n2091 ,n1834);
    or g422(n2345 ,n2090 ,n1833);
    or g423(n2344 ,n2088 ,n1832);
    or g424(n2343 ,n2087 ,n1831);
    or g425(n2342 ,n2086 ,n1830);
    or g426(n2341 ,n2084 ,n1829);
    or g427(n2340 ,n2083 ,n1828);
    or g428(n2339 ,n2082 ,n1827);
    or g429(n2338 ,n2081 ,n1826);
    or g430(n2337 ,n2079 ,n1825);
    or g431(n2336 ,n2077 ,n1824);
    or g432(n2335 ,n2075 ,n1823);
    or g433(n2334 ,n2074 ,n1822);
    or g434(n2333 ,n2073 ,n1821);
    or g435(n2332 ,n2071 ,n1820);
    or g436(n2331 ,n2070 ,n1819);
    or g437(n2330 ,n2068 ,n1818);
    or g438(n2329 ,n2067 ,n1817);
    or g439(n2328 ,n2135 ,n1863);
    or g440(n2327 ,n2065 ,n1815);
    or g441(n2326 ,n2063 ,n1814);
    or g442(n2325 ,n2062 ,n1813);
    or g443(n2324 ,n2060 ,n1812);
    or g444(n2323 ,n2059 ,n1811);
    or g445(n2322 ,n2058 ,n1810);
    or g446(n2321 ,n2057 ,n1809);
    or g447(n2320 ,n2054 ,n1808);
    or g448(n2319 ,n2053 ,n1807);
    or g449(n2318 ,n2052 ,n1806);
    or g450(n2317 ,n2050 ,n1805);
    or g451(n2316 ,n2048 ,n1804);
    or g452(n2315 ,n2046 ,n1803);
    or g453(n2314 ,n2045 ,n1802);
    or g454(n2313 ,n2043 ,n1801);
    or g455(n2312 ,n1733 ,n1988);
    or g456(n2311 ,n1735 ,n1992);
    or g457(n2310 ,n1734 ,n1990);
    or g458(n2309 ,n1732 ,n1989);
    or g459(n2308 ,n1731 ,n1986);
    or g460(n2307 ,n1730 ,n1987);
    or g461(n2306 ,n1729 ,n1984);
    or g462(n2305 ,n1709 ,n1982);
    or g463(n2304 ,n1727 ,n1983);
    or g464(n2303 ,n1716 ,n1981);
    or g465(n2302 ,n1726 ,n1975);
    or g466(n2301 ,n1725 ,n1979);
    or g467(n2300 ,n1724 ,n1980);
    or g468(n2299 ,n1723 ,n1978);
    or g469(n2298 ,n1728 ,n1985);
    or g470(n2297 ,n1722 ,n1977);
    or g471(n2296 ,n1594 ,n1976);
    or g472(n2295 ,n1721 ,n1974);
    or g473(n2294 ,n1720 ,n1971);
    or g474(n2293 ,n1623 ,n1973);
    or g475(n2292 ,n1719 ,n1972);
    or g476(n2291 ,n1718 ,n1970);
    or g477(n2290 ,n1717 ,n1969);
    or g478(n2289 ,n1666 ,n1968);
    or g479(n2288 ,n1715 ,n1967);
    or g480(n2287 ,n1711 ,n1957);
    or g481(n2286 ,n1682 ,n1965);
    or g482(n2285 ,n1683 ,n1966);
    or g483(n2284 ,n1713 ,n1964);
    or g484(n2283 ,n1710 ,n1961);
    or g485(n2282 ,n1563 ,n1963);
    or g486(n2281 ,n1708 ,n1962);
    or g487(n2280 ,n1591 ,n1912);
    or g488(n2279 ,n1707 ,n1959);
    or g489(n2278 ,n1706 ,n1958);
    or g490(n2277 ,n1705 ,n1956);
    or g491(n2276 ,n1590 ,n1955);
    or g492(n2275 ,n1703 ,n1954);
    or g493(n2274 ,n1656 ,n1951);
    or g494(n2273 ,n1665 ,n1952);
    or g495(n2272 ,n1701 ,n1950);
    or g496(n2271 ,n1700 ,n1948);
    or g497(n2270 ,n1704 ,n1949);
    or g498(n2269 ,n1699 ,n1947);
    or g499(n2268 ,n1702 ,n1953);
    or g500(n2267 ,n1714 ,n1946);
    or g501(n2266 ,n1698 ,n1945);
    or g502(n2265 ,n1694 ,n1941);
    or g503(n2264 ,n1697 ,n1944);
    or g504(n2263 ,n1603 ,n1943);
    or g505(n2262 ,n1611 ,n1942);
    or g506(n2261 ,n1691 ,n1936);
    or g507(n2260 ,n1695 ,n1940);
    or g508(n2259 ,n1692 ,n1939);
    or g509(n2258 ,n1645 ,n1938);
    or g510(n2257 ,n1660 ,n1937);
    or g511(n2256 ,n1688 ,n1935);
    or g512(n2255 ,n1684 ,n1934);
    or g513(n2254 ,n1679 ,n1933);
    or g514(n2253 ,n1670 ,n1931);
    or g515(n2252 ,n1674 ,n1932);
    or g516(n2251 ,n1668 ,n1930);
    or g517(n2250 ,n1662 ,n1929);
    or g518(n2249 ,n1657 ,n1928);
    or g519(n2248 ,n1651 ,n1927);
    or g520(n2247 ,n1649 ,n1926);
    or g521(n2246 ,n1643 ,n1925);
    or g522(n2245 ,n1640 ,n1924);
    or g523(n2244 ,n1634 ,n1923);
    or g524(n2243 ,n1631 ,n1922);
    or g525(n2242 ,n1626 ,n1921);
    or g526(n2241 ,n1622 ,n1920);
    or g527(n2240 ,n1617 ,n1919);
    or g528(n2239 ,n1614 ,n1918);
    or g529(n2238 ,n1609 ,n1916);
    or g530(n2237 ,n1605 ,n1915);
    or g531(n2236 ,n1601 ,n1914);
    or g532(n2235 ,n1597 ,n1913);
    or g533(n2234 ,n1593 ,n1911);
    or g534(n2233 ,n1589 ,n1909);
    or g535(n2232 ,n1567 ,n1960);
    or g536(n2231 ,n1588 ,n1910);
    or g537(n2230 ,n1586 ,n1908);
    or g538(n2229 ,n1577 ,n1900);
    or g539(n2228 ,n1585 ,n1907);
    or g540(n2227 ,n1587 ,n1906);
    or g541(n2226 ,n1584 ,n1904);
    or g542(n2225 ,n1583 ,n1905);
    or g543(n2224 ,n1582 ,n1903);
    or g544(n2223 ,n1581 ,n1901);
    or g545(n2222 ,n1580 ,n1902);
    or g546(n2221 ,n1579 ,n1899);
    or g547(n2220 ,n1576 ,n1898);
    or g548(n2219 ,n1575 ,n1897);
    or g549(n2218 ,n1598 ,n1917);
    or g550(n2217 ,n1574 ,n1896);
    or g551(n2216 ,n1573 ,n1895);
    or g552(n2215 ,n1572 ,n1894);
    or g553(n2214 ,n1571 ,n1893);
    or g554(n2213 ,n1570 ,n1892);
    or g555(n2212 ,n1568 ,n1891);
    or g556(n2211 ,n1569 ,n1887);
    or g557(n2210 ,n1635 ,n1888);
    or g558(n2209 ,n1566 ,n1889);
    or g559(n2208 ,n1646 ,n1886);
    or g560(n2207 ,n1565 ,n1883);
    or g561(n2206 ,n1564 ,n1885);
    or g562(n2205 ,n1464 ,n1875);
    or g563(n2204 ,n1562 ,n1884);
    or g564(n2203 ,n1465 ,n1881);
    or g565(n2202 ,n1800 ,n1882);
    or g566(n2201 ,n1463 ,n1880);
    or g567(n2200 ,n1461 ,n1878);
    or g568(n2199 ,n1462 ,n1879);
    or g569(n2198 ,n1460 ,n1877);
    or g570(n2197 ,n1459 ,n1876);
    or g571(n2196 ,n1712 ,n1874);
    or g572(n2195 ,n1457 ,n1871);
    or g573(n2194 ,n1456 ,n1872);
    or g574(n2193 ,n1455 ,n1870);
    or g575(n2192 ,n1453 ,n1869);
    or g576(n2191 ,n1458 ,n1868);
    or g577(n2190 ,n1454 ,n1873);
    or g578(n2189 ,n1452 ,n1867);
    or g579(n2188 ,n1451 ,n1890);
    or g580(n2187 ,n1450 ,n1866);
    or g581(n2186 ,n1578 ,n1865);
    or g582(n2185 ,n1449 ,n1991);
    nor g583(n2184 ,n682 ,n1466);
    nor g584(n2183 ,n618 ,n1559);
    nor g585(n2182 ,n609 ,n1513);
    nor g586(n2181 ,n698 ,n1524);
    nor g587(n2180 ,n568 ,n1560);
    nor g588(n2179 ,n574 ,n1519);
    nor g589(n2178 ,n668 ,n1552);
    nor g590(n2177 ,n556 ,n1495);
    nor g591(n2176 ,n708 ,n1515);
    nor g592(n2175 ,n350 ,n1556);
    nor g593(n2174 ,n579 ,n1494);
    nor g594(n2173 ,n674 ,n1512);
    nor g595(n2172 ,n683 ,n1493);
    nor g596(n2171 ,n362 ,n1492);
    nor g597(n2170 ,n548 ,n1558);
    nor g598(n2169 ,n703 ,n1472);
    nor g599(n2168 ,n590 ,n1490);
    nor g600(n2167 ,n704 ,n1506);
    nor g601(n2166 ,n597 ,n1488);
    nor g602(n2165 ,n612 ,n1489);
    nor g603(n2164 ,n635 ,n1505);
    nor g604(n2163 ,n659 ,n1487);
    nor g605(n2162 ,n620 ,n1486);
    nor g606(n2161 ,n644 ,n1504);
    nor g607(n2160 ,n586 ,n1485);
    nor g608(n2159 ,n686 ,n1484);
    nor g609(n2158 ,n550 ,n1535);
    nor g610(n2157 ,n691 ,n1482);
    nor g611(n2156 ,n552 ,n1480);
    nor g612(n2155 ,n608 ,n1500);
    nor g613(n2154 ,n374 ,n1521);
    nor g614(n2153 ,n610 ,n1478);
    nor g615(n2152 ,n695 ,n1499);
    nor g616(n2151 ,n335 ,n1477);
    nor g617(n2150 ,n341 ,n1555);
    nor g618(n2149 ,n599 ,n1476);
    nor g619(n2148 ,n557 ,n1498);
    nor g620(n2147 ,n592 ,n1475);
    nor g621(n2146 ,n555 ,n1474);
    nor g622(n2145 ,n702 ,n1557);
    nor g623(n2144 ,n562 ,n1497);
    nor g624(n2143 ,n573 ,n1473);
    nor g625(n2142 ,n303 ,n1554);
    nor g626(n2141 ,n379 ,n1471);
    nor g627(n2140 ,n542 ,n1553);
    nor g628(n2139 ,n603 ,n1470);
    nor g629(n2138 ,n626 ,n1469);
    nor g630(n2137 ,n352 ,n1481);
    nor g631(n2136 ,n699 ,n1467);
    nor g632(n2135 ,n688 ,n1501);
    nor g633(n2134 ,n375 ,n1513);
    nor g634(n2133 ,n630 ,n1502);
    nor g635(n2132 ,n588 ,n1560);
    nor g636(n2131 ,n613 ,n1510);
    nor g637(n2130 ,n650 ,n1552);
    nor g638(n2129 ,n677 ,n1551);
    nor g639(n2128 ,n651 ,n1549);
    nor g640(n2127 ,n658 ,n1550);
    nor g641(n2126 ,n619 ,n1548);
    nor g642(n2125 ,n594 ,n1546);
    nor g643(n2124 ,n641 ,n1547);
    nor g644(n2123 ,n640 ,n1545);
    nor g645(n2122 ,n643 ,n1544);
    nor g646(n2121 ,n652 ,n1542);
    nor g647(n2120 ,n563 ,n1543);
    nor g648(n2119 ,n583 ,n1541);
    nor g649(n2118 ,n631 ,n1540);
    nor g650(n2117 ,n578 ,n1539);
    nor g651(n2116 ,n587 ,n1538);
    nor g652(n2115 ,n710 ,n1537);
    nor g653(n2114 ,n600 ,n1534);
    nor g654(n2113 ,n566 ,n1536);
    nor g655(n2112 ,n576 ,n1533);
    nor g656(n2111 ,n584 ,n1532);
    nor g657(n2110 ,n622 ,n1530);
    nor g658(n2109 ,n377 ,n1531);
    nor g659(n2108 ,n606 ,n1529);
    nor g660(n2107 ,n329 ,n1527);
    nor g661(n2106 ,n678 ,n1528);
    nor g662(n2105 ,n689 ,n1526);
    nor g663(n2104 ,n661 ,n1525);
    nor g664(n2103 ,n564 ,n1524);
    nor g665(n2102 ,n585 ,n1523);
    nor g666(n2101 ,n546 ,n1522);
    nor g667(n2100 ,n633 ,n1520);
    nor g668(n2099 ,n628 ,n1519);
    nor g669(n2098 ,n667 ,n1518);
    nor g670(n2097 ,n671 ,n1517);
    nor g671(n2096 ,n569 ,n1515);
    nor g672(n2095 ,n605 ,n1516);
    nor g673(n2094 ,n638 ,n1514);
    nor g674(n2093 ,n705 ,n1561);
    nor g675(n2092 ,n611 ,n1512);
    nor g676(n2091 ,n595 ,n1511);
    nor g677(n2090 ,n554 ,n1509);
    nor g678(n2089 ,n642 ,n1508);
    nor g679(n2088 ,n575 ,n1553);
    nor g680(n2087 ,n675 ,n1501);
    nor g681(n2086 ,n636 ,n1510);
    nor g682(n2085 ,n343 ,n1506);
    nor g683(n2084 ,n353 ,n1551);
    nor g684(n2083 ,n561 ,n1550);
    nor g685(n2082 ,n567 ,n1548);
    nor g686(n2081 ,n582 ,n1547);
    nor g687(n2080 ,n323 ,n1496);
    nor g688(n2079 ,n701 ,n1545);
    nor g689(n2078 ,n709 ,n1505);
    nor g690(n2077 ,n572 ,n1544);
    nor g691(n2076 ,n580 ,n1504);
    nor g692(n2075 ,n627 ,n1542);
    nor g693(n2074 ,n601 ,n1541);
    nor g694(n2073 ,n545 ,n1540);
    nor g695(n2072 ,n334 ,n1503);
    nor g696(n2071 ,n634 ,n1538);
    nor g697(n2070 ,n565 ,n1537);
    nor g698(n2069 ,n616 ,n1500);
    nor g699(n2068 ,n615 ,n1536);
    nor g700(n2067 ,n687 ,n1533);
    nor g701(n2066 ,n662 ,n1532);
    nor g702(n2065 ,n646 ,n1530);
    nor g703(n2064 ,n607 ,n1499);
    nor g704(n2063 ,n604 ,n1529);
    nor g705(n2062 ,n670 ,n1528);
    nor g706(n2061 ,n621 ,n1466);
    nor g707(n2060 ,n623 ,n1526);
    nor g708(n2059 ,n680 ,n1525);
    nor g709(n2058 ,n571 ,n1523);
    nor g710(n2057 ,n570 ,n1522);
    nor g711(n2056 ,n694 ,n1498);
    nor g712(n2055 ,n657 ,n1497);
    nor g713(n2054 ,n669 ,n1520);
    nor g714(n2053 ,n581 ,n1518);
    nor g715(n2052 ,n617 ,n1517);
    nor g716(n2051 ,n697 ,n1496);
    nor g717(n2050 ,n551 ,n1516);
    nor g718(n2049 ,n645 ,n1508);
    nor g719(n2048 ,n700 ,n1514);
    nor g720(n2047 ,n558 ,n1491);
    nor g721(n2046 ,n543 ,n1561);
    nor g722(n2045 ,n692 ,n1511);
    nor g723(n2044 ,n639 ,n1507);
    nor g724(n2043 ,n553 ,n1509);
    nor g725(n2042 ,n632 ,n1495);
    nor g726(n2041 ,n577 ,n1479);
    nor g727(n2040 ,n707 ,n1556);
    nor g728(n2039 ,n560 ,n1468);
    nor g729(n2038 ,n649 ,n1494);
    nor g730(n2037 ,n330 ,n1493);
    nor g731(n2036 ,n306 ,n1492);
    nor g732(n2035 ,n376 ,n1483);
    nor g733(n2034 ,n696 ,n1472);
    nor g734(n2033 ,n625 ,n1491);
    nor g735(n2032 ,n681 ,n1559);
    nor g736(n2031 ,n660 ,n1490);
    nor g737(n2030 ,n693 ,n1488);
    nor g738(n2029 ,n685 ,n1558);
    nor g739(n2028 ,n647 ,n1489);
    nor g740(n2027 ,n596 ,n1487);
    nor g741(n2026 ,n679 ,n1535);
    nor g742(n2025 ,n655 ,n1486);
    nor g743(n2024 ,n663 ,n1507);
    nor g744(n2023 ,n338 ,n1485);
    nor g745(n2022 ,n593 ,n1555);
    nor g746(n2021 ,n666 ,n1484);
    nor g747(n2020 ,n672 ,n1554);
    nor g748(n2019 ,n624 ,n1482);
    nor g749(n2018 ,n591 ,n1480);
    nor g750(n2017 ,n312 ,n1502);
    nor g751(n2016 ,n665 ,n1521);
    nor g752(n2015 ,n602 ,n1478);
    nor g753(n2014 ,n340 ,n1549);
    nor g754(n2013 ,n559 ,n1479);
    nor g755(n2012 ,n351 ,n1477);
    nor g756(n2011 ,n549 ,n1476);
    nor g757(n2010 ,n664 ,n1546);
    nor g758(n2009 ,n614 ,n1475);
    nor g759(n2008 ,n373 ,n1543);
    nor g760(n2007 ,n648 ,n1474);
    nor g761(n2006 ,n544 ,n1468);
    nor g762(n2005 ,n690 ,n1557);
    nor g763(n2004 ,n629 ,n1539);
    nor g764(n2003 ,n673 ,n1473);
    nor g765(n2002 ,n327 ,n1471);
    nor g766(n2001 ,n684 ,n1534);
    nor g767(n2000 ,n653 ,n1470);
    nor g768(n1999 ,n656 ,n1503);
    nor g769(n1998 ,n547 ,n1469);
    nor g770(n1997 ,n706 ,n1531);
    nor g771(n1996 ,n598 ,n1481);
    nor g772(n1995 ,n637 ,n1483);
    nor g773(n1994 ,n654 ,n1467);
    nor g774(n1993 ,n676 ,n1527);
    nor g775(n1992 ,n1016 ,n1448);
    nor g776(n1991 ,n1165 ,n1447);
    nor g777(n1990 ,n1065 ,n1446);
    nor g778(n1989 ,n1148 ,n1444);
    nor g779(n1988 ,n1092 ,n1445);
    nor g780(n1987 ,n1164 ,n1440);
    nor g781(n1986 ,n1127 ,n1442);
    nor g782(n1985 ,n1163 ,n1443);
    nor g783(n1984 ,n1129 ,n1412);
    nor g784(n1983 ,n1144 ,n1439);
    nor g785(n1982 ,n1140 ,n1419);
    nor g786(n1981 ,n1072 ,n1438);
    nor g787(n1980 ,n1150 ,n1437);
    nor g788(n1979 ,n1151 ,n1436);
    nor g789(n1978 ,n1162 ,n1441);
    nor g790(n1977 ,n1023 ,n1434);
    nor g791(n1976 ,n1030 ,n1372);
    nor g792(n1975 ,n1155 ,n1435);
    nor g793(n1974 ,n1149 ,n1433);
    nor g794(n1973 ,n1102 ,n1432);
    nor g795(n1972 ,n1067 ,n1431);
    nor g796(n1971 ,n1096 ,n1389);
    nor g797(n1970 ,n1063 ,n1388);
    nor g798(n1969 ,n1098 ,n1430);
    nor g799(n1968 ,n1086 ,n1390);
    nor g800(n1967 ,n1147 ,n1428);
    nor g801(n1966 ,n1118 ,n1427);
    nor g802(n1965 ,n1047 ,n1426);
    nor g803(n1964 ,n985 ,n1425);
    nor g804(n1963 ,n1137 ,n1424);
    nor g805(n1962 ,n1115 ,n1422);
    nor g806(n1961 ,n987 ,n1423);
    nor g807(n1960 ,n1034 ,n1421);
    nor g808(n1959 ,n1139 ,n1420);
    nor g809(n1958 ,n997 ,n1358);
    nor g810(n1957 ,n1012 ,n1418);
    nor g811(n1956 ,n1136 ,n1378);
    nor g812(n1955 ,n1161 ,n1364);
    nor g813(n1954 ,n1130 ,n1417);
    nor g814(n1953 ,n1128 ,n1414);
    nor g815(n1952 ,n1126 ,n1416);
    nor g816(n1951 ,n1095 ,n1415);
    nor g817(n1950 ,n1120 ,n1413);
    nor g818(n1949 ,n1133 ,n1411);
    nor g819(n1948 ,n1125 ,n1410);
    nor g820(n1947 ,n990 ,n1409);
    nor g821(n1946 ,n975 ,n1408);
    nor g822(n1945 ,n1145 ,n1406);
    nor g823(n1944 ,n1060 ,n1405);
    nor g824(n1943 ,n1018 ,n1404);
    nor g825(n1942 ,n1044 ,n1403);
    nor g826(n1941 ,n1124 ,n1407);
    nor g827(n1940 ,n1156 ,n1380);
    nor g828(n1939 ,n1169 ,n1402);
    nor g829(n1938 ,n1024 ,n1401);
    nor g830(n1937 ,n1103 ,n1400);
    nor g831(n1936 ,n1111 ,n1399);
    nor g832(n1935 ,n1159 ,n1398);
    nor g833(n1934 ,n1146 ,n1397);
    nor g834(n1933 ,n1113 ,n1396);
    nor g835(n1932 ,n1109 ,n1395);
    nor g836(n1931 ,n1104 ,n1394);
    nor g837(n1930 ,n1093 ,n1393);
    nor g838(n1929 ,n1090 ,n1392);
    nor g839(n1928 ,n1082 ,n1391);
    nor g840(n1927 ,n1079 ,n1387);
    nor g841(n1926 ,n1074 ,n1386);
    nor g842(n1925 ,n1066 ,n1384);
    nor g843(n1924 ,n979 ,n1383);
    nor g844(n1923 ,n1138 ,n1382);
    nor g845(n1922 ,n1049 ,n1381);
    nor g846(n1921 ,n1045 ,n1379);
    nor g847(n1920 ,n1039 ,n1377);
    nor g848(n1919 ,n1036 ,n1376);
    nor g849(n1918 ,n1033 ,n1375);
    nor g850(n1917 ,n1007 ,n1354);
    nor g851(n1916 ,n1029 ,n1374);
    nor g852(n1915 ,n998 ,n1373);
    nor g853(n1914 ,n1008 ,n1370);
    nor g854(n1913 ,n1019 ,n1369);
    nor g855(n1912 ,n1132 ,n1367);
    nor g856(n1911 ,n1123 ,n1368);
    nor g857(n1910 ,n1142 ,n1365);
    nor g858(n1909 ,n1015 ,n1366);
    nor g859(n1908 ,n1013 ,n1363);
    nor g860(n1907 ,n1009 ,n1362);
    nor g861(n1906 ,n1011 ,n1361);
    nor g862(n1905 ,n1006 ,n1360);
    nor g863(n1904 ,n983 ,n1326);
    nor g864(n1903 ,n984 ,n1359);
    nor g865(n1902 ,n993 ,n1357);
    nor g866(n1901 ,n991 ,n1355);
    nor g867(n1900 ,n1152 ,n1349);
    nor g868(n1899 ,n1003 ,n1353);
    nor g869(n1898 ,n1010 ,n1356);
    nor g870(n1897 ,n995 ,n1352);
    nor g871(n1896 ,n1021 ,n1351);
    nor g872(n1895 ,n1001 ,n1371);
    nor g873(n1894 ,n1025 ,n1350);
    nor g874(n1893 ,n1084 ,n1348);
    nor g875(n1892 ,n1000 ,n1347);
    nor g876(n1891 ,n1042 ,n1346);
    nor g877(n1890 ,n1002 ,n1322);
    nor g878(n1889 ,n1054 ,n1345);
    nor g879(n1888 ,n1058 ,n1344);
    nor g880(n1887 ,n999 ,n1343);
    nor g881(n1886 ,n1070 ,n1385);
    nor g882(n1885 ,n996 ,n1342);
    nor g883(n1884 ,n1107 ,n1340);
    nor g884(n1883 ,n1089 ,n1341);
    nor g885(n1882 ,n994 ,n1338);
    nor g886(n1881 ,n992 ,n1339);
    nor g887(n1880 ,n1121 ,n1336);
    nor g888(n1879 ,n989 ,n1333);
    nor g889(n1878 ,n988 ,n1334);
    nor g890(n1877 ,n1135 ,n1429);
    nor g891(n1876 ,n1131 ,n1332);
    nor g892(n1875 ,n1134 ,n1337);
    nor g893(n1874 ,n1154 ,n1331);
    nor g894(n1873 ,n976 ,n1324);
    nor g895(n1872 ,n1153 ,n1330);
    nor g896(n1871 ,n982 ,n1329);
    nor g897(n1870 ,n1116 ,n1328);
    nor g898(n1869 ,n1014 ,n1335);
    nor g899(n1868 ,n981 ,n1327);
    nor g900(n1867 ,n1158 ,n1325);
    nor g901(n1866 ,n1062 ,n1323);
    nor g902(n1865 ,n986 ,n1321);
    or g903(n1864 ,n1696 ,n1799);
    or g904(n1863 ,n1693 ,n1798);
    or g905(n1862 ,n1663 ,n1797);
    or g906(n1861 ,n1690 ,n1796);
    or g907(n1860 ,n1689 ,n1795);
    or g908(n1859 ,n1687 ,n1794);
    or g909(n1858 ,n1686 ,n1793);
    or g910(n1857 ,n1685 ,n1792);
    or g911(n1856 ,n1681 ,n1791);
    or g912(n1855 ,n1680 ,n1790);
    or g913(n1854 ,n1678 ,n1789);
    or g914(n1853 ,n1677 ,n1788);
    or g915(n1852 ,n1676 ,n1787);
    or g916(n1851 ,n1675 ,n1786);
    or g917(n1850 ,n1673 ,n1785);
    or g918(n1849 ,n1672 ,n1784);
    or g919(n1848 ,n1671 ,n1783);
    or g920(n1847 ,n1669 ,n1782);
    or g921(n1846 ,n1667 ,n1781);
    or g922(n1845 ,n1664 ,n1780);
    or g923(n1844 ,n1661 ,n1779);
    or g924(n1843 ,n1659 ,n1778);
    or g925(n1842 ,n1658 ,n1777);
    or g926(n1841 ,n1655 ,n1776);
    or g927(n1840 ,n1654 ,n1775);
    or g928(n1839 ,n1653 ,n1774);
    or g929(n1838 ,n1652 ,n1773);
    or g930(n1837 ,n1650 ,n1772);
    or g931(n1836 ,n1648 ,n1771);
    or g932(n1835 ,n1647 ,n1770);
    or g933(n1834 ,n1644 ,n1769);
    or g934(n1833 ,n1642 ,n1768);
    or g935(n1832 ,n1641 ,n1767);
    or g936(n1831 ,n1639 ,n1766);
    or g937(n1830 ,n1638 ,n1765);
    or g938(n1829 ,n1637 ,n1764);
    or g939(n1828 ,n1636 ,n1763);
    or g940(n1827 ,n1633 ,n1762);
    or g941(n1826 ,n1632 ,n1761);
    or g942(n1825 ,n1630 ,n1760);
    or g943(n1824 ,n1629 ,n1759);
    or g944(n1823 ,n1628 ,n1758);
    or g945(n1822 ,n1627 ,n1757);
    or g946(n1821 ,n1625 ,n1756);
    or g947(n1820 ,n1624 ,n1755);
    or g948(n1819 ,n1621 ,n1754);
    or g949(n1818 ,n1620 ,n1753);
    or g950(n1817 ,n1619 ,n1752);
    or g951(n1816 ,n1618 ,n1751);
    or g952(n1815 ,n1616 ,n1750);
    or g953(n1814 ,n1615 ,n1749);
    or g954(n1813 ,n1613 ,n1748);
    or g955(n1812 ,n1612 ,n1747);
    or g956(n1811 ,n1610 ,n1746);
    or g957(n1810 ,n1608 ,n1745);
    or g958(n1809 ,n1607 ,n1744);
    or g959(n1808 ,n1606 ,n1743);
    or g960(n1807 ,n1604 ,n1742);
    or g961(n1806 ,n1602 ,n1741);
    or g962(n1805 ,n1600 ,n1740);
    or g963(n1804 ,n1599 ,n1739);
    or g964(n1803 ,n1596 ,n1738);
    or g965(n1802 ,n1595 ,n1737);
    or g966(n1801 ,n1592 ,n1736);
    nor g967(n1800 ,n5[44] ,n1301);
    nor g968(n1799 ,n1099 ,n1274);
    nor g969(n1798 ,n1122 ,n1214);
    nor g970(n1797 ,n1087 ,n1273);
    nor g971(n1796 ,n978 ,n1272);
    nor g972(n1795 ,n977 ,n1271);
    nor g973(n1794 ,n1157 ,n1270);
    nor g974(n1793 ,n1097 ,n1269);
    nor g975(n1792 ,n1052 ,n1268);
    nor g976(n1791 ,n1143 ,n1267);
    nor g977(n1790 ,n1160 ,n1265);
    nor g978(n1789 ,n1114 ,n1264);
    nor g979(n1788 ,n1112 ,n1263);
    nor g980(n1787 ,n1110 ,n1262);
    nor g981(n1786 ,n1108 ,n1261);
    nor g982(n1785 ,n1106 ,n1260);
    nor g983(n1784 ,n1105 ,n1259);
    nor g984(n1783 ,n1101 ,n1258);
    nor g985(n1782 ,n1141 ,n1257);
    nor g986(n1781 ,n1094 ,n1256);
    nor g987(n1780 ,n1166 ,n1255);
    nor g988(n1779 ,n1091 ,n1266);
    nor g989(n1778 ,n1088 ,n1234);
    nor g990(n1777 ,n1085 ,n1233);
    nor g991(n1776 ,n1083 ,n1231);
    nor g992(n1775 ,n1081 ,n1229);
    nor g993(n1774 ,n1080 ,n1228);
    nor g994(n1773 ,n1078 ,n1226);
    nor g995(n1772 ,n1076 ,n1224);
    nor g996(n1771 ,n1075 ,n1222);
    nor g997(n1770 ,n1073 ,n1221);
    nor g998(n1769 ,n1071 ,n1219);
    nor g999(n1768 ,n1069 ,n1218);
    nor g1000(n1767 ,n1064 ,n1217);
    nor g1001(n1766 ,n1100 ,n1215);
    nor g1002(n1765 ,n1117 ,n1213);
    nor g1003(n1764 ,n1061 ,n1212);
    nor g1004(n1763 ,n1057 ,n1210);
    nor g1005(n1762 ,n1056 ,n1209);
    nor g1006(n1761 ,n1053 ,n1208);
    nor g1007(n1760 ,n1050 ,n1206);
    nor g1008(n1759 ,n1017 ,n1204);
    nor g1009(n1758 ,n1048 ,n1207);
    nor g1010(n1757 ,n1051 ,n1202);
    nor g1011(n1756 ,n1043 ,n1200);
    nor g1012(n1755 ,n1041 ,n1199);
    nor g1013(n1754 ,n1040 ,n1198);
    nor g1014(n1753 ,n1038 ,n1197);
    nor g1015(n1752 ,n1037 ,n1196);
    nor g1016(n1751 ,n1022 ,n1194);
    nor g1017(n1750 ,n1035 ,n1193);
    nor g1018(n1749 ,n1068 ,n1191);
    nor g1019(n1748 ,n1077 ,n1190);
    nor g1020(n1747 ,n1032 ,n1189);
    nor g1021(n1746 ,n1031 ,n1192);
    nor g1022(n1745 ,n1046 ,n1195);
    nor g1023(n1744 ,n1028 ,n1201);
    nor g1024(n1743 ,n1027 ,n1203);
    nor g1025(n1742 ,n1026 ,n1205);
    nor g1026(n1741 ,n1004 ,n1211);
    nor g1027(n1740 ,n1005 ,n1216);
    nor g1028(n1739 ,n1020 ,n1220);
    nor g1029(n1738 ,n1059 ,n1223);
    nor g1030(n1737 ,n980 ,n1225);
    nor g1031(n1736 ,n1119 ,n1227);
    nor g1032(n1735 ,n4[28] ,n1283);
    nor g1033(n1734 ,n4[29] ,n1282);
    nor g1034(n1733 ,n5[51] ,n1293);
    nor g1035(n1732 ,n4[30] ,n1281);
    nor g1036(n1731 ,n4[31] ,n1280);
    nor g1037(n1730 ,n5[52] ,n1292);
    nor g1038(n1729 ,n4[32] ,n1279);
    nor g1039(n1728 ,n5[5] ,n1308);
    nor g1040(n1727 ,n5[53] ,n1291);
    nor g1041(n1726 ,n5[6] ,n1305);
    nor g1042(n1725 ,n5[54] ,n1290);
    nor g1043(n1724 ,n4[35] ,n1306);
    nor g1044(n1723 ,n4[36] ,n1307);
    nor g1045(n1722 ,n5[55] ,n1289);
    nor g1046(n1721 ,n4[38] ,n1305);
    nor g1047(n1720 ,n5[7] ,n1304);
    nor g1048(n1719 ,n5[56] ,n1288);
    nor g1049(n1718 ,n4[40] ,n1277);
    nor g1050(n1717 ,n5[57] ,n1287);
    nor g1051(n1716 ,n4[34] ,n1286);
    nor g1052(n1715 ,n4[42] ,n1303);
    nor g1053(n1714 ,n4[55] ,n1289);
    nor g1054(n1713 ,n4[44] ,n1301);
    nor g1055(n1712 ,n4[21] ,n1291);
    nor g1056(n1711 ,n5[8] ,n1277);
    nor g1057(n1710 ,n5[59] ,n1284);
    nor g1058(n1709 ,n4[33] ,n1278);
    nor g1059(n1708 ,n4[46] ,n1298);
    nor g1060(n1707 ,n5[60] ,n1283);
    nor g1061(n1706 ,n4[48] ,n1296);
    nor g1062(n1705 ,n5[61] ,n1282);
    nor g1063(n1704 ,n4[53] ,n1291);
    nor g1064(n1703 ,n4[50] ,n1294);
    nor g1065(n1702 ,n5[9] ,n1299);
    nor g1066(n1701 ,n4[52] ,n1292);
    nor g1067(n1700 ,n5[63] ,n1280);
    nor g1068(n1699 ,n4[54] ,n1290);
    nor g1069(n1698 ,n4[56] ,n1288);
    nor g1070(n1697 ,n4[57] ,n1287);
    nor g1071(n1696 ,n3[0] ,n1279);
    nor g1072(n1695 ,n4[60] ,n1283);
    nor g1073(n1694 ,n5[10] ,n1303);
    nor g1074(n1693 ,n3[1] ,n1278);
    nor g1075(n1692 ,n4[61] ,n1282);
    nor g1076(n1691 ,n5[11] ,n1302);
    nor g1077(n1690 ,n3[3] ,n1306);
    nor g1078(n1689 ,n3[4] ,n1307);
    nor g1079(n1688 ,n5[12] ,n1301);
    nor g1080(n1687 ,n3[5] ,n1308);
    nor g1081(n1686 ,n3[6] ,n1305);
    nor g1082(n1685 ,n3[7] ,n1304);
    nor g1083(n1684 ,n5[13] ,n1300);
    nor g1084(n1683 ,n4[43] ,n1302);
    nor g1085(n1682 ,n5[58] ,n1285);
    nor g1086(n1681 ,n3[8] ,n1277);
    nor g1087(n1680 ,n3[9] ,n1299);
    nor g1088(n1679 ,n5[14] ,n1298);
    nor g1089(n1678 ,n3[10] ,n1303);
    nor g1090(n1677 ,n3[11] ,n1302);
    nor g1091(n1676 ,n3[12] ,n1301);
    nor g1092(n1675 ,n3[13] ,n1300);
    nor g1093(n1674 ,n5[15] ,n1297);
    nor g1094(n1673 ,n3[14] ,n1298);
    nor g1095(n1672 ,n3[15] ,n1297);
    nor g1096(n1671 ,n3[16] ,n1296);
    nor g1097(n1670 ,n5[16] ,n1296);
    nor g1098(n1669 ,n3[17] ,n1295);
    nor g1099(n1668 ,n5[17] ,n1295);
    nor g1100(n1667 ,n3[18] ,n1294);
    nor g1101(n1666 ,n4[41] ,n1299);
    nor g1102(n1665 ,n4[51] ,n1293);
    nor g1103(n1664 ,n3[19] ,n1293);
    nor g1104(n1663 ,n3[2] ,n1286);
    nor g1105(n1662 ,n5[18] ,n1294);
    nor g1106(n1661 ,n3[20] ,n1292);
    nor g1107(n1660 ,n4[63] ,n1280);
    nor g1108(n1659 ,n3[21] ,n1291);
    nor g1109(n1658 ,n3[22] ,n1290);
    nor g1110(n1657 ,n5[19] ,n1293);
    nor g1111(n1656 ,n5[62] ,n1281);
    nor g1112(n1655 ,n3[23] ,n1289);
    nor g1113(n1654 ,n3[24] ,n1288);
    nor g1114(n1653 ,n3[25] ,n1287);
    nor g1115(n1652 ,n3[26] ,n1285);
    nor g1116(n1651 ,n5[20] ,n1292);
    nor g1117(n1650 ,n3[27] ,n1284);
    nor g1118(n1649 ,n5[21] ,n1291);
    nor g1119(n1648 ,n3[28] ,n1283);
    nor g1120(n1647 ,n3[29] ,n1282);
    nor g1121(n1646 ,n4[14] ,n1298);
    nor g1122(n1645 ,n4[62] ,n1281);
    nor g1123(n1644 ,n3[30] ,n1281);
    nor g1124(n1643 ,n5[22] ,n1290);
    nor g1125(n1642 ,n3[31] ,n1280);
    nor g1126(n1641 ,n3[32] ,n1279);
    nor g1127(n1640 ,n5[23] ,n1289);
    nor g1128(n1639 ,n3[33] ,n1278);
    nor g1129(n1638 ,n3[34] ,n1286);
    nor g1130(n1637 ,n3[35] ,n1306);
    nor g1131(n1636 ,n3[36] ,n1307);
    nor g1132(n1635 ,n5[42] ,n1303);
    nor g1133(n1634 ,n5[24] ,n1288);
    nor g1134(n1633 ,n3[37] ,n1308);
    nor g1135(n1632 ,n3[38] ,n1305);
    nor g1136(n1631 ,n5[25] ,n1287);
    nor g1137(n1630 ,n3[39] ,n1304);
    nor g1138(n1629 ,n3[40] ,n1277);
    nor g1139(n1628 ,n3[41] ,n1299);
    nor g1140(n1627 ,n3[42] ,n1303);
    nor g1141(n1626 ,n5[26] ,n1285);
    nor g1142(n1625 ,n3[43] ,n1302);
    nor g1143(n1624 ,n3[44] ,n1301);
    nor g1144(n1623 ,n4[39] ,n1304);
    nor g1145(n1622 ,n5[27] ,n1284);
    nor g1146(n1621 ,n3[45] ,n1300);
    nor g1147(n1620 ,n3[46] ,n1298);
    nor g1148(n1619 ,n3[47] ,n1297);
    nor g1149(n1618 ,n3[48] ,n1296);
    nor g1150(n1617 ,n5[28] ,n1283);
    nor g1151(n1616 ,n3[49] ,n1295);
    nor g1152(n1615 ,n3[50] ,n1294);
    nor g1153(n1614 ,n5[29] ,n1282);
    nor g1154(n1613 ,n3[51] ,n1293);
    nor g1155(n1612 ,n3[52] ,n1292);
    nor g1156(n1611 ,n4[59] ,n1284);
    nor g1157(n1610 ,n3[53] ,n1291);
    nor g1158(n1609 ,n5[30] ,n1281);
    nor g1159(n1608 ,n3[54] ,n1290);
    nor g1160(n1607 ,n3[55] ,n1289);
    nor g1161(n1606 ,n3[56] ,n1288);
    nor g1162(n1605 ,n5[31] ,n1280);
    nor g1163(n1604 ,n3[57] ,n1287);
    nor g1164(n1603 ,n4[58] ,n1285);
    nor g1165(n1602 ,n3[58] ,n1285);
    nor g1166(n1601 ,n5[32] ,n1279);
    nor g1167(n1600 ,n3[59] ,n1284);
    nor g1168(n1599 ,n3[60] ,n1283);
    nor g1169(n1598 ,n5[0] ,n1279);
    nor g1170(n1597 ,n5[33] ,n1278);
    nor g1171(n1596 ,n3[61] ,n1282);
    nor g1172(n1595 ,n3[62] ,n1281);
    nor g1173(n1594 ,n4[37] ,n1308);
    nor g1174(n1593 ,n5[34] ,n1286);
    nor g1175(n1592 ,n3[63] ,n1280);
    nor g1176(n1591 ,n4[0] ,n1279);
    nor g1177(n1590 ,n4[49] ,n1295);
    nor g1178(n1589 ,n5[35] ,n1306);
    nor g1179(n1588 ,n4[1] ,n1278);
    nor g1180(n1587 ,n5[36] ,n1307);
    nor g1181(n1586 ,n4[2] ,n1286);
    nor g1182(n1585 ,n4[3] ,n1306);
    nor g1183(n1584 ,n4[4] ,n1307);
    nor g1184(n1583 ,n5[37] ,n1308);
    nor g1185(n1582 ,n4[5] ,n1308);
    nor g1186(n1581 ,n5[38] ,n1305);
    nor g1187(n1580 ,n4[6] ,n1305);
    nor g1188(n1579 ,n4[7] ,n1304);
    nor g1189(n1578 ,n4[27] ,n1284);
    nor g1190(n1577 ,n5[1] ,n1278);
    nor g1191(n1576 ,n5[39] ,n1304);
    nor g1192(n1575 ,n4[8] ,n1277);
    nor g1193(n1574 ,n4[9] ,n1299);
    nor g1194(n1573 ,n5[40] ,n1277);
    nor g1195(n1572 ,n4[10] ,n1303);
    nor g1196(n1571 ,n4[11] ,n1302);
    nor g1197(n1570 ,n5[41] ,n1299);
    nor g1198(n1569 ,n5[2] ,n1286);
    nor g1199(n1568 ,n4[12] ,n1301);
    nor g1200(n1567 ,n4[47] ,n1297);
    nor g1201(n1566 ,n4[13] ,n1300);
    nor g1202(n1565 ,n5[43] ,n1302);
    nor g1203(n1564 ,n4[15] ,n1297);
    nor g1204(n1563 ,n4[45] ,n1300);
    nor g1205(n1562 ,n4[16] ,n1296);
    nor g1206(n1465 ,n4[17] ,n1295);
    nor g1207(n1464 ,n5[3] ,n1306);
    nor g1208(n1463 ,n4[18] ,n1294);
    nor g1209(n1462 ,n5[45] ,n1300);
    nor g1210(n1461 ,n4[19] ,n1293);
    nor g1211(n1460 ,n4[20] ,n1292);
    nor g1212(n1459 ,n5[46] ,n1298);
    nor g1213(n1458 ,n4[24] ,n1288);
    nor g1214(n1457 ,n5[47] ,n1297);
    nor g1215(n1456 ,n4[22] ,n1290);
    nor g1216(n1455 ,n4[23] ,n1289);
    nor g1217(n1454 ,n5[4] ,n1307);
    nor g1218(n1453 ,n5[48] ,n1296);
    nor g1219(n1452 ,n4[25] ,n1287);
    nor g1220(n1451 ,n5[49] ,n1295);
    nor g1221(n1450 ,n4[26] ,n1285);
    nor g1222(n1449 ,n5[50] ,n1294);
    or g1223(n1448 ,n767 ,n1275);
    or g1224(n1447 ,n884 ,n1276);
    or g1225(n1446 ,n821 ,n1275);
    or g1226(n1445 ,n870 ,n1276);
    or g1227(n1444 ,n787 ,n1275);
    or g1228(n1443 ,n784 ,n1276);
    or g1229(n1442 ,n872 ,n1275);
    or g1230(n1441 ,n907 ,n1275);
    or g1231(n1440 ,n876 ,n1276);
    or g1232(n1439 ,n881 ,n1276);
    or g1233(n1438 ,n887 ,n1275);
    or g1234(n1437 ,n894 ,n1275);
    or g1235(n1436 ,n901 ,n1276);
    or g1236(n1435 ,n889 ,n1276);
    or g1237(n1434 ,n781 ,n1276);
    or g1238(n1433 ,n774 ,n1275);
    or g1239(n1432 ,n822 ,n1275);
    or g1240(n1431 ,n789 ,n1276);
    or g1241(n1430 ,n837 ,n1276);
    or g1242(n1429 ,n771 ,n1275);
    or g1243(n1428 ,n856 ,n1275);
    or g1244(n1427 ,n860 ,n1275);
    or g1245(n1426 ,n891 ,n1276);
    or g1246(n1425 ,n903 ,n1275);
    or g1247(n1424 ,n880 ,n1275);
    or g1248(n1423 ,n863 ,n1276);
    or g1249(n1422 ,n818 ,n1275);
    or g1250(n1421 ,n717 ,n1275);
    or g1251(n1420 ,n745 ,n1276);
    or g1252(n1419 ,n897 ,n1275);
    or g1253(n1418 ,n761 ,n1276);
    or g1254(n1417 ,n801 ,n1275);
    or g1255(n1416 ,n869 ,n1275);
    or g1256(n1415 ,n865 ,n1276);
    or g1257(n1414 ,n751 ,n1276);
    or g1258(n1413 ,n812 ,n1275);
    or g1259(n1412 ,n814 ,n1275);
    or g1260(n1411 ,n772 ,n1275);
    or g1261(n1410 ,n795 ,n1276);
    or g1262(n1409 ,n734 ,n1275);
    or g1263(n1408 ,n720 ,n1275);
    or g1264(n1407 ,n743 ,n1276);
    or g1265(n1406 ,n896 ,n1275);
    or g1266(n1405 ,n763 ,n1275);
    or g1267(n1404 ,n851 ,n1275);
    or g1268(n1403 ,n769 ,n1275);
    or g1269(n1402 ,n804 ,n1275);
    or g1270(n1401 ,n866 ,n1275);
    or g1271(n1400 ,n839 ,n1275);
    or g1272(n1399 ,n861 ,n1276);
    or g1273(n1398 ,n859 ,n1276);
    or g1274(n1397 ,n846 ,n1276);
    or g1275(n1396 ,n741 ,n1276);
    or g1276(n1395 ,n847 ,n1276);
    or g1277(n1394 ,n840 ,n1276);
    or g1278(n1393 ,n835 ,n1276);
    or g1279(n1392 ,n726 ,n1276);
    or g1280(n1391 ,n824 ,n1276);
    or g1281(n1390 ,n831 ,n1275);
    or g1282(n1389 ,n886 ,n1276);
    or g1283(n1388 ,n813 ,n1275);
    or g1284(n1387 ,n817 ,n1276);
    or g1285(n1386 ,n793 ,n1276);
    or g1286(n1385 ,n791 ,n1275);
    or g1287(n1384 ,n807 ,n1276);
    or g1288(n1383 ,n796 ,n1276);
    or g1289(n1382 ,n780 ,n1276);
    or g1290(n1381 ,n754 ,n1276);
    or g1291(n1380 ,n836 ,n1275);
    or g1292(n1379 ,n832 ,n1276);
    or g1293(n1378 ,n864 ,n1276);
    or g1294(n1377 ,n899 ,n1276);
    or g1295(n1376 ,n775 ,n1276);
    or g1296(n1375 ,n828 ,n1276);
    or g1297(n1374 ,n719 ,n1276);
    or g1298(n1373 ,n747 ,n1276);
    or g1299(n1372 ,n735 ,n1275);
    or g1300(n1371 ,n748 ,n1276);
    or g1301(n1370 ,n885 ,n1276);
    or g1302(n1369 ,n941 ,n1276);
    or g1303(n1368 ,n905 ,n1276);
    or g1304(n1367 ,n752 ,n1275);
    or g1305(n1366 ,n857 ,n1276);
    or g1306(n1365 ,n750 ,n1275);
    or g1307(n1364 ,n757 ,n1275);
    or g1308(n1363 ,n890 ,n1275);
    or g1309(n1362 ,n802 ,n1275);
    or g1310(n1361 ,n892 ,n1276);
    or g1311(n1360 ,n718 ,n1276);
    or g1312(n1359 ,n722 ,n1275);
    or g1313(n1358 ,n898 ,n1275);
    or g1314(n1357 ,n888 ,n1275);
    or g1315(n1356 ,n738 ,n1276);
    or g1316(n1355 ,n731 ,n1276);
    or g1317(n1354 ,n746 ,n1276);
    or g1318(n1353 ,n733 ,n1275);
    or g1319(n1352 ,n768 ,n1275);
    or g1320(n1351 ,n737 ,n1275);
    or g1321(n1350 ,n766 ,n1275);
    or g1322(n1349 ,n755 ,n1276);
    or g1323(n1348 ,n773 ,n1275);
    or g1324(n1347 ,n883 ,n1276);
    or g1325(n1346 ,n786 ,n1275);
    or g1326(n1345 ,n797 ,n1275);
    or g1327(n1344 ,n724 ,n1276);
    or g1328(n1343 ,n816 ,n1276);
    or g1329(n1342 ,n715 ,n1275);
    or g1330(n1341 ,n858 ,n1276);
    or g1331(n1340 ,n723 ,n1275);
    or g1332(n1339 ,n855 ,n1275);
    or g1333(n1338 ,n871 ,n1276);
    or g1334(n1337 ,n877 ,n1276);
    or g1335(n1336 ,n867 ,n1275);
    or g1336(n1335 ,n744 ,n1276);
    or g1337(n1334 ,n862 ,n1275);
    or g1338(n1333 ,n875 ,n1276);
    or g1339(n1332 ,n882 ,n1276);
    or g1340(n1331 ,n842 ,n1275);
    or g1341(n1330 ,n902 ,n1275);
    or g1342(n1329 ,n904 ,n1276);
    or g1343(n1328 ,n893 ,n1275);
    or g1344(n1327 ,n728 ,n1275);
    or g1345(n1326 ,n895 ,n1275);
    or g1346(n1325 ,n825 ,n1275);
    or g1347(n1324 ,n849 ,n1276);
    or g1348(n1323 ,n800 ,n1275);
    or g1349(n1322 ,n873 ,n1276);
    or g1350(n1321 ,n749 ,n1275);
    nor g1351(n1561 ,n1253 ,n1185);
    nor g1352(n1560 ,n277 ,n1254);
    nor g1353(n1559 ,n276 ,n1309);
    nor g1354(n1558 ,n276 ,n1250);
    nor g1355(n1557 ,n277 ,n1244);
    nor g1356(n1556 ,n277 ,n1241);
    nor g1357(n1555 ,n276 ,n1311);
    nor g1358(n1554 ,n276 ,n1320);
    nor g1359(n1553 ,n1242 ,n1185);
    nor g1360(n1552 ,n277 ,n1251);
    nor g1361(n1551 ,n1239 ,n1185);
    nor g1362(n1550 ,n1238 ,n1185);
    nor g1363(n1549 ,n276 ,n1312);
    nor g1364(n1548 ,n1240 ,n1185);
    nor g1365(n1547 ,n1309 ,n1185);
    nor g1366(n1546 ,n276 ,n1318);
    nor g1367(n1545 ,n1250 ,n1185);
    nor g1368(n1544 ,n1314 ,n1185);
    nor g1369(n1543 ,n276 ,n1316);
    nor g1370(n1542 ,n1311 ,n1185);
    nor g1371(n1541 ,n1320 ,n1185);
    nor g1372(n1540 ,n1243 ,n1185);
    nor g1373(n1539 ,n276 ,n1319);
    nor g1374(n1538 ,n1312 ,n1185);
    nor g1375(n1537 ,n1318 ,n1185);
    nor g1376(n1536 ,n1316 ,n1185);
    nor g1377(n1535 ,n276 ,n1314);
    nor g1378(n1534 ,n276 ,n1317);
    nor g1379(n1533 ,n1319 ,n1185);
    nor g1380(n1532 ,n1317 ,n1185);
    nor g1381(n1531 ,n276 ,n1313);
    nor g1382(n1530 ,n1313 ,n1185);
    nor g1383(n1529 ,n1315 ,n1185);
    nor g1384(n1528 ,n1235 ,n1185);
    nor g1385(n1527 ,n276 ,n1315);
    nor g1386(n1526 ,n1237 ,n1185);
    nor g1387(n1525 ,n1244 ,n1185);
    nor g1388(n1524 ,n276 ,n1235);
    nor g1389(n1523 ,n1245 ,n1185);
    nor g1390(n1522 ,n1246 ,n1185);
    nor g1391(n1521 ,n277 ,n1319);
    nor g1392(n1520 ,n1247 ,n1185);
    nor g1393(n1519 ,n276 ,n1237);
    nor g1394(n1518 ,n1248 ,n1185);
    nor g1395(n1517 ,n1249 ,n1185);
    nor g1396(n1516 ,n1236 ,n1185);
    nor g1397(n1515 ,n276 ,n1244);
    nor g1398(n1514 ,n1252 ,n1185);
    nor g1399(n1513 ,n277 ,n1253);
    nor g1400(n1512 ,n276 ,n1245);
    nor g1401(n1511 ,n1254 ,n1185);
    nor g1402(n1510 ,n1310 ,n1185);
    nor g1403(n1509 ,n1251 ,n1185);
    nor g1404(n1508 ,n276 ,n1246);
    nor g1405(n1507 ,n276 ,n1310);
    nor g1406(n1506 ,n276 ,n1247);
    nor g1407(n1505 ,n276 ,n1248);
    nor g1408(n1504 ,n276 ,n1249);
    nor g1409(n1503 ,n276 ,n1236);
    nor g1410(n1502 ,n276 ,n1243);
    nor g1411(n1501 ,n1241 ,n1185);
    nor g1412(n1500 ,n276 ,n1252);
    nor g1413(n1499 ,n276 ,n1253);
    nor g1414(n1498 ,n276 ,n1254);
    nor g1415(n1497 ,n276 ,n1251);
    nor g1416(n1496 ,n276 ,n1242);
    nor g1417(n1495 ,n277 ,n1242);
    nor g1418(n1494 ,n277 ,n1310);
    nor g1419(n1493 ,n277 ,n1239);
    nor g1420(n1492 ,n277 ,n1238);
    nor g1421(n1491 ,n276 ,n1241);
    nor g1422(n1490 ,n277 ,n1309);
    nor g1423(n1489 ,n277 ,n1314);
    nor g1424(n1488 ,n277 ,n1250);
    nor g1425(n1487 ,n277 ,n1311);
    nor g1426(n1486 ,n277 ,n1320);
    nor g1427(n1485 ,n277 ,n1243);
    nor g1428(n1484 ,n277 ,n1312);
    nor g1429(n1483 ,n276 ,n1240);
    nor g1430(n1482 ,n277 ,n1318);
    nor g1431(n1481 ,n277 ,n1249);
    nor g1432(n1480 ,n277 ,n1316);
    nor g1433(n1479 ,n276 ,n1239);
    nor g1434(n1478 ,n277 ,n1317);
    nor g1435(n1477 ,n277 ,n1313);
    nor g1436(n1476 ,n277 ,n1315);
    nor g1437(n1475 ,n277 ,n1235);
    nor g1438(n1474 ,n277 ,n1237);
    nor g1439(n1473 ,n277 ,n1245);
    nor g1440(n1472 ,n277 ,n1240);
    nor g1441(n1471 ,n277 ,n1246);
    nor g1442(n1470 ,n277 ,n1247);
    nor g1443(n1469 ,n277 ,n1248);
    nor g1444(n1468 ,n276 ,n1238);
    nor g1445(n1467 ,n277 ,n1236);
    nor g1446(n1466 ,n277 ,n1252);
    or g1447(n1274 ,n794 ,n1187);
    or g1448(n1273 ,n878 ,n1187);
    or g1449(n1272 ,n736 ,n1187);
    or g1450(n1271 ,n730 ,n1187);
    or g1451(n1270 ,n753 ,n1187);
    or g1452(n1269 ,n739 ,n1187);
    or g1453(n1268 ,n879 ,n1187);
    or g1454(n1267 ,n756 ,n1187);
    or g1455(n1266 ,n830 ,n1187);
    or g1456(n1265 ,n844 ,n1187);
    or g1457(n1264 ,n854 ,n1187);
    or g1458(n1263 ,n853 ,n1187);
    or g1459(n1262 ,n850 ,n1187);
    or g1460(n1261 ,n848 ,n1187);
    or g1461(n1260 ,n826 ,n1187);
    or g1462(n1259 ,n843 ,n1187);
    or g1463(n1258 ,n721 ,n1187);
    or g1464(n1257 ,n838 ,n1187);
    or g1465(n1256 ,n834 ,n1187);
    or g1466(n1255 ,n806 ,n1187);
    nor g1467(n1320 ,n8[10] ,n279);
    nor g1468(n1319 ,n8[15] ,n279);
    nor g1469(n1318 ,n8[13] ,n279);
    nor g1470(n1317 ,n8[16] ,n279);
    nor g1471(n1316 ,n8[14] ,n279);
    nor g1472(n1315 ,n8[18] ,n279);
    nor g1473(n1314 ,n8[8] ,n279);
    nor g1474(n1313 ,n8[17] ,n279);
    nor g1475(n1312 ,n8[12] ,n279);
    nor g1476(n1311 ,n8[9] ,n279);
    nor g1477(n1310 ,n8[2] ,n279);
    nor g1478(n1309 ,n8[6] ,n279);
    or g1479(n1308 ,n289 ,n278);
    or g1480(n1307 ,n533 ,n278);
    or g1481(n1306 ,n538 ,n278);
    or g1482(n1305 ,n521 ,n278);
    or g1483(n1304 ,n531 ,n278);
    or g1484(n1303 ,n526 ,n278);
    or g1485(n1302 ,n522 ,n278);
    or g1486(n1301 ,n516 ,n278);
    or g1487(n1300 ,n529 ,n278);
    or g1488(n1299 ,n520 ,n278);
    or g1489(n1298 ,n291 ,n278);
    or g1490(n1297 ,n515 ,n278);
    or g1491(n1296 ,n525 ,n278);
    or g1492(n1295 ,n534 ,n278);
    or g1493(n1294 ,n539 ,n278);
    or g1494(n1293 ,n513 ,n278);
    or g1495(n1292 ,n524 ,n278);
    or g1496(n1291 ,n532 ,n278);
    or g1497(n1290 ,n536 ,n278);
    or g1498(n1289 ,n518 ,n278);
    or g1499(n1288 ,n535 ,n278);
    or g1500(n1287 ,n528 ,n278);
    or g1501(n1286 ,n519 ,n278);
    or g1502(n1285 ,n517 ,n278);
    or g1503(n1284 ,n537 ,n278);
    or g1504(n1283 ,n530 ,n278);
    or g1505(n1282 ,n527 ,n278);
    or g1506(n1281 ,n523 ,n278);
    or g1507(n1280 ,n293 ,n278);
    or g1508(n1279 ,n292 ,n278);
    or g1509(n1278 ,n290 ,n278);
    or g1510(n1277 ,n514 ,n278);
    or g1511(n1276 ,n1181 ,n1184);
    or g1512(n1275 ,n1179 ,n1183);
    or g1513(n1234 ,n829 ,n1187);
    or g1514(n1233 ,n732 ,n1187);
    nor g1515(n1232 ,n287 ,n1182);
    or g1516(n1231 ,n758 ,n1187);
    nor g1517(n1230 ,n288 ,n1186);
    or g1518(n1229 ,n823 ,n1187);
    or g1519(n1228 ,n819 ,n1187);
    or g1520(n1227 ,n742 ,n1187);
    or g1521(n1226 ,n845 ,n1187);
    or g1522(n1225 ,n841 ,n1187);
    or g1523(n1224 ,n815 ,n1187);
    or g1524(n1223 ,n820 ,n1187);
    or g1525(n1222 ,n811 ,n1187);
    or g1526(n1221 ,n810 ,n1187);
    or g1527(n1220 ,n777 ,n1187);
    or g1528(n1219 ,n809 ,n1187);
    or g1529(n1218 ,n805 ,n1187);
    or g1530(n1217 ,n833 ,n1187);
    or g1531(n1216 ,n759 ,n1187);
    or g1532(n1215 ,n906 ,n1187);
    or g1533(n1214 ,n798 ,n1187);
    or g1534(n1213 ,n799 ,n1187);
    or g1535(n1212 ,n868 ,n1187);
    or g1536(n1211 ,n740 ,n1187);
    or g1537(n1210 ,n792 ,n1187);
    or g1538(n1209 ,n790 ,n1187);
    or g1539(n1208 ,n788 ,n1187);
    or g1540(n1207 ,n776 ,n1187);
    or g1541(n1206 ,n803 ,n1187);
    or g1542(n1205 ,n729 ,n1187);
    or g1543(n1204 ,n785 ,n1187);
    or g1544(n1203 ,n727 ,n1187);
    or g1545(n1202 ,n783 ,n1187);
    or g1546(n1201 ,n716 ,n1187);
    or g1547(n1200 ,n782 ,n1187);
    or g1548(n1199 ,n900 ,n1187);
    or g1549(n1198 ,n874 ,n1187);
    or g1550(n1197 ,n779 ,n1187);
    or g1551(n1196 ,n764 ,n1187);
    or g1552(n1195 ,n725 ,n1187);
    or g1553(n1194 ,n762 ,n1187);
    or g1554(n1193 ,n778 ,n1187);
    or g1555(n1192 ,n765 ,n1187);
    or g1556(n1191 ,n770 ,n1187);
    or g1557(n1190 ,n808 ,n1187);
    or g1558(n1189 ,n852 ,n1187);
    nor g1559(n1254 ,n8[30] ,n279);
    nor g1560(n1253 ,n8[29] ,n279);
    nor g1561(n1252 ,n8[28] ,n279);
    nor g1562(n1251 ,n8[31] ,n279);
    nor g1563(n1250 ,n8[7] ,n279);
    nor g1564(n1249 ,n8[26] ,n279);
    nor g1565(n1248 ,n8[25] ,n279);
    nor g1566(n1247 ,n8[24] ,n279);
    nor g1567(n1246 ,n8[23] ,n279);
    nor g1568(n1245 ,n8[22] ,n279);
    nor g1569(n1244 ,n8[21] ,n279);
    nor g1570(n1243 ,n8[11] ,n279);
    nor g1571(n1242 ,n10[0] ,n279);
    nor g1572(n1241 ,n10[1] ,n279);
    nor g1573(n1240 ,n8[5] ,n279);
    nor g1574(n1239 ,n8[3] ,n279);
    nor g1575(n1238 ,n8[4] ,n279);
    nor g1576(n1237 ,n8[20] ,n279);
    nor g1577(n1236 ,n8[27] ,n279);
    nor g1578(n1235 ,n8[19] ,n279);
    not g1579(n279 ,n1188);
    not g1580(n278 ,n1188);
    nor g1581(n1186 ,n1177 ,n1175);
    nor g1582(n1188 ,n942 ,n1176);
    or g1583(n1187 ,n714 ,n1176);
    not g1584(n277 ,n1184);
    not g1585(n276 ,n1183);
    xnor g1586(n1182 ,n1171 ,n9[0]);
    nor g1587(n1185 ,n288 ,n1174);
    or g1588(n1184 ,n287 ,n1178);
    or g1589(n1183 ,n287 ,n1180);
    not g1590(n1181 ,n1180);
    not g1591(n1179 ,n1178);
    nor g1592(n1177 ,n541 ,n1171);
    nor g1593(n1180 ,n541 ,n1170);
    nor g1594(n1178 ,n540 ,n1170);
    nor g1595(n1175 ,n1170 ,n1173);
    nor g1596(n1174 ,n1172 ,n1170);
    or g1597(n1176 ,n287 ,n1170);
    not g1598(n1173 ,n1172);
    not g1599(n1170 ,n1171);
    xnor g1600(n1172 ,n540 ,n9[1]);
    nor g1601(n1171 ,n1168 ,n1055);
    nor g1602(n1169 ,n527 ,n507);
    or g1603(n1168 ,n589 ,n711);
    nor g1604(n1167 ,n364 ,n287);
    nor g1605(n1166 ,n513 ,n301);
    nor g1606(n1165 ,n539 ,n391);
    nor g1607(n1164 ,n524 ,n417);
    nor g1608(n1163 ,n289 ,n429);
    nor g1609(n1162 ,n533 ,n508);
    nor g1610(n1161 ,n534 ,n499);
    nor g1611(n1160 ,n520 ,n355);
    nor g1612(n1159 ,n516 ,n458);
    nor g1613(n1158 ,n528 ,n472);
    nor g1614(n1157 ,n289 ,n349);
    nor g1615(n1156 ,n530 ,n496);
    nor g1616(n1155 ,n521 ,n442);
    nor g1617(n1154 ,n532 ,n497);
    nor g1618(n1153 ,n536 ,n468);
    nor g1619(n1152 ,n441 ,n290);
    nor g1620(n1151 ,n536 ,n437);
    nor g1621(n1150 ,n538 ,n505);
    nor g1622(n1149 ,n521 ,n487);
    nor g1623(n1148 ,n523 ,n490);
    nor g1624(n1147 ,n526 ,n382);
    nor g1625(n1146 ,n529 ,n398);
    nor g1626(n1145 ,n535 ,n387);
    nor g1627(n1144 ,n532 ,n485);
    nor g1628(n1143 ,n514 ,n295);
    nor g1629(n1142 ,n446 ,n290);
    nor g1630(n1141 ,n534 ,n300);
    nor g1631(n1140 ,n392 ,n290);
    nor g1632(n1139 ,n530 ,n413);
    nor g1633(n1138 ,n535 ,n390);
    nor g1634(n1137 ,n529 ,n488);
    nor g1635(n1136 ,n527 ,n422);
    nor g1636(n1135 ,n524 ,n448);
    nor g1637(n1134 ,n538 ,n394);
    nor g1638(n1133 ,n532 ,n495);
    nor g1639(n1132 ,n460 ,n292);
    nor g1640(n1131 ,n291 ,n455);
    nor g1641(n1130 ,n539 ,n438);
    nor g1642(n1129 ,n424 ,n292);
    nor g1643(n1128 ,n520 ,n404);
    nor g1644(n1127 ,n293 ,n463);
    nor g1645(n1126 ,n513 ,n471);
    nor g1646(n1125 ,n293 ,n457);
    nor g1647(n1124 ,n526 ,n433);
    nor g1648(n1123 ,n519 ,n397);
    nor g1649(n1122 ,n314 ,n290);
    nor g1650(n1121 ,n539 ,n486);
    nor g1651(n1120 ,n524 ,n426);
    nor g1652(n1119 ,n293 ,n346);
    nor g1653(n1118 ,n522 ,n479);
    nor g1654(n1117 ,n519 ,n320);
    nor g1655(n1116 ,n518 ,n450);
    nor g1656(n1115 ,n291 ,n465);
    nor g1657(n1114 ,n526 ,n326);
    nor g1658(n1113 ,n291 ,n427);
    nor g1659(n1112 ,n522 ,n363);
    nor g1660(n1111 ,n522 ,n477);
    nor g1661(n1110 ,n516 ,n308);
    nor g1662(n1109 ,n515 ,n464);
    nor g1663(n1108 ,n529 ,n310);
    nor g1664(n1107 ,n525 ,n484);
    nor g1665(n1106 ,n291 ,n369);
    nor g1666(n1105 ,n515 ,n358);
    nor g1667(n1104 ,n525 ,n452);
    nor g1668(n1103 ,n293 ,n449);
    nor g1669(n1102 ,n531 ,n443);
    nor g1670(n1101 ,n525 ,n342);
    nor g1671(n1100 ,n356 ,n290);
    nor g1672(n1099 ,n313 ,n292);
    nor g1673(n1098 ,n528 ,n384);
    nor g1674(n1097 ,n521 ,n371);
    nor g1675(n1096 ,n531 ,n444);
    nor g1676(n1095 ,n523 ,n416);
    nor g1677(n1094 ,n539 ,n299);
    nor g1678(n1093 ,n534 ,n428);
    nor g1679(n1092 ,n513 ,n423);
    nor g1680(n1091 ,n524 ,n378);
    nor g1681(n1090 ,n539 ,n406);
    nor g1682(n1089 ,n522 ,n466);
    nor g1683(n1088 ,n532 ,n297);
    nor g1684(n1087 ,n519 ,n332);
    nor g1685(n1086 ,n520 ,n474);
    nor g1686(n1085 ,n536 ,n325);
    nor g1687(n1084 ,n522 ,n476);
    nor g1688(n1083 ,n518 ,n344);
    nor g1689(n1082 ,n513 ,n400);
    nor g1690(n1081 ,n535 ,n360);
    nor g1691(n1080 ,n528 ,n381);
    nor g1692(n1079 ,n524 ,n454);
    nor g1693(n1078 ,n517 ,n298);
    nor g1694(n1077 ,n513 ,n364);
    nor g1695(n1076 ,n537 ,n296);
    nor g1696(n1075 ,n530 ,n337);
    nor g1697(n1074 ,n532 ,n462);
    nor g1698(n1073 ,n527 ,n324);
    nor g1699(n1072 ,n519 ,n480);
    nor g1700(n1071 ,n523 ,n361);
    nor g1701(n1070 ,n291 ,n451);
    nor g1702(n1069 ,n293 ,n354);
    nor g1703(n1068 ,n539 ,n302);
    nor g1704(n1067 ,n535 ,n407);
    nor g1705(n1066 ,n536 ,n509);
    nor g1706(n1065 ,n527 ,n421);
    nor g1707(n1064 ,n372 ,n292);
    nor g1708(n1063 ,n514 ,n478);
    nor g1709(n1062 ,n517 ,n445);
    nor g1710(n1061 ,n538 ,n365);
    nor g1711(n1060 ,n528 ,n396);
    nor g1712(n1059 ,n527 ,n318);
    nor g1713(n1058 ,n526 ,n411);
    nor g1714(n1057 ,n533 ,n294);
    nor g1715(n1056 ,n289 ,n319);
    or g1716(n1055 ,n713 ,n712);
    nor g1717(n1054 ,n529 ,n401);
    nor g1718(n1053 ,n521 ,n317);
    nor g1719(n1052 ,n531 ,n368);
    nor g1720(n1051 ,n526 ,n348);
    nor g1721(n1050 ,n531 ,n347);
    nor g1722(n1049 ,n528 ,n481);
    nor g1723(n1048 ,n520 ,n357);
    nor g1724(n1047 ,n517 ,n461);
    nor g1725(n1046 ,n536 ,n380);
    nor g1726(n1045 ,n517 ,n506);
    nor g1727(n1044 ,n537 ,n453);
    nor g1728(n1043 ,n522 ,n304);
    nor g1729(n1042 ,n516 ,n415);
    nor g1730(n1041 ,n516 ,n333);
    nor g1731(n1040 ,n529 ,n366);
    nor g1732(n1039 ,n537 ,n473);
    nor g1733(n1038 ,n291 ,n307);
    nor g1734(n1037 ,n515 ,n305);
    nor g1735(n1036 ,n530 ,n493);
    nor g1736(n1035 ,n534 ,n359);
    nor g1737(n1034 ,n515 ,n459);
    nor g1738(n1033 ,n527 ,n470);
    nor g1739(n1032 ,n524 ,n311);
    nor g1740(n1031 ,n532 ,n331);
    nor g1741(n1030 ,n289 ,n494);
    nor g1742(n1029 ,n523 ,n435);
    nor g1743(n1028 ,n518 ,n339);
    nor g1744(n1027 ,n535 ,n370);
    nor g1745(n1026 ,n528 ,n345);
    nor g1746(n1025 ,n526 ,n388);
    nor g1747(n1024 ,n523 ,n482);
    nor g1748(n1023 ,n518 ,n504);
    nor g1749(n1022 ,n525 ,n321);
    nor g1750(n1021 ,n520 ,n412);
    nor g1751(n1020 ,n530 ,n309);
    nor g1752(n1019 ,n385 ,n290);
    nor g1753(n1018 ,n517 ,n440);
    nor g1754(n1017 ,n514 ,n328);
    nor g1755(n1016 ,n530 ,n383);
    nor g1756(n1015 ,n538 ,n419);
    nor g1757(n1014 ,n525 ,n491);
    nor g1758(n1013 ,n519 ,n425);
    nor g1759(n1012 ,n514 ,n475);
    nor g1760(n1011 ,n533 ,n410);
    nor g1761(n1010 ,n531 ,n469);
    nor g1762(n1009 ,n538 ,n409);
    nor g1763(n1008 ,n418 ,n292);
    nor g1764(n1007 ,n439 ,n292);
    nor g1765(n1006 ,n289 ,n500);
    nor g1766(n1005 ,n537 ,n315);
    nor g1767(n1004 ,n517 ,n316);
    nor g1768(n1003 ,n531 ,n393);
    nor g1769(n1002 ,n534 ,n399);
    nor g1770(n1001 ,n514 ,n456);
    nor g1771(n1000 ,n520 ,n431);
    nor g1772(n999 ,n519 ,n432);
    nor g1773(n998 ,n293 ,n395);
    nor g1774(n997 ,n525 ,n492);
    nor g1775(n996 ,n515 ,n436);
    nor g1776(n995 ,n514 ,n498);
    nor g1777(n994 ,n516 ,n386);
    nor g1778(n993 ,n521 ,n430);
    nor g1779(n992 ,n534 ,n403);
    nor g1780(n991 ,n521 ,n402);
    nor g1781(n990 ,n536 ,n420);
    nor g1782(n989 ,n529 ,n414);
    nor g1783(n988 ,n513 ,n447);
    nor g1784(n987 ,n537 ,n503);
    nor g1785(n986 ,n537 ,n405);
    nor g1786(n985 ,n516 ,n467);
    nor g1787(n984 ,n289 ,n483);
    nor g1788(n983 ,n533 ,n408);
    nor g1789(n982 ,n515 ,n489);
    nor g1790(n981 ,n535 ,n502);
    nor g1791(n980 ,n523 ,n336);
    nor g1792(n979 ,n518 ,n389);
    nor g1793(n978 ,n538 ,n322);
    nor g1794(n977 ,n533 ,n367);
    nor g1795(n976 ,n533 ,n501);
    nor g1796(n975 ,n518 ,n434);
    nor g1797(n974 ,n370 ,n281);
    nor g1798(n973 ,n299 ,n288);
    nor g1799(n972 ,n307 ,n288);
    nor g1800(n971 ,n349 ,n287);
    nor g1801(n970 ,n368 ,n287);
    nor g1802(n969 ,n308 ,n282);
    nor g1803(n968 ,n304 ,n282);
    nor g1804(n967 ,n346 ,n281);
    nor g1805(n966 ,n296 ,n282);
    nor g1806(n965 ,n510 ,n280);
    nor g1807(n964 ,n309 ,n284);
    nor g1808(n963 ,n305 ,n280);
    nor g1809(n962 ,n361 ,n280);
    nor g1810(n961 ,n512 ,n284);
    nor g1811(n960 ,n511 ,n286);
    nor g1812(n959 ,n324 ,n284);
    nor g1813(n958 ,n358 ,n285);
    nor g1814(n957 ,n294 ,n280);
    nor g1815(n956 ,n336 ,n285);
    nor g1816(n955 ,n302 ,n281);
    nor g1817(n954 ,n314 ,n285);
    nor g1818(n953 ,n369 ,n285);
    nor g1819(n952 ,n310 ,n282);
    nor g1820(n951 ,n348 ,n282);
    nor g1821(n950 ,n339 ,n285);
    nor g1822(n949 ,n326 ,n280);
    nor g1823(n948 ,n328 ,n284);
    nor g1824(n947 ,n347 ,n286);
    nor g1825(n946 ,n337 ,n284);
    nor g1826(n945 ,n321 ,n280);
    nor g1827(n944 ,n316 ,n281);
    nor g1828(n943 ,n371 ,n282);
    or g1829(n942 ,n540 ,n541);
    nor g1830(n941 ,n2539 ,n10[1]);
    nor g1831(n940 ,n315 ,n286);
    nor g1832(n939 ,n300 ,n286);
    nor g1833(n938 ,n317 ,n288);
    nor g1834(n937 ,n378 ,n288);
    nor g1835(n936 ,n363 ,n283);
    nor g1836(n935 ,n354 ,n283);
    nor g1837(n934 ,n313 ,n283);
    nor g1838(n933 ,n372 ,n283);
    nor g1839(n932 ,n318 ,n287);
    nor g1840(n931 ,n365 ,n287);
    nor g1841(n930 ,n356 ,n284);
    nor g1842(n929 ,n301 ,n283);
    nor g1843(n928 ,n344 ,n285);
    nor g1844(n927 ,n331 ,n285);
    nor g1845(n926 ,n367 ,n285);
    nor g1846(n925 ,n319 ,n284);
    nor g1847(n924 ,n366 ,n282);
    nor g1848(n923 ,n332 ,n282);
    nor g1849(n922 ,n311 ,n281);
    nor g1850(n921 ,n298 ,n287);
    nor g1851(n920 ,n342 ,n283);
    nor g1852(n919 ,n380 ,n286);
    nor g1853(n918 ,n297 ,n284);
    nor g1854(n917 ,n325 ,n283);
    nor g1855(n916 ,n360 ,n281);
    nor g1856(n915 ,n359 ,n280);
    nor g1857(n914 ,n357 ,n287);
    nor g1858(n913 ,n322 ,n288);
    nor g1859(n912 ,n333 ,n286);
    nor g1860(n911 ,n355 ,n286);
    nor g1861(n910 ,n381 ,n280);
    nor g1862(n909 ,n345 ,n281);
    nor g1863(n908 ,n295 ,n286);
    nor g1864(n907 ,n8[4] ,n2[100]);
    nor g1865(n906 ,n2[33] ,n10[1]);
    nor g1866(n905 ,n8[2] ,n2540);
    nor g1867(n904 ,n8[15] ,n2553);
    nor g1868(n903 ,n8[12] ,n2[108]);
    nor g1869(n902 ,n8[22] ,n2[86]);
    nor g1870(n901 ,n8[22] ,n2560);
    nor g1871(n900 ,n8[12] ,n2[44]);
    nor g1872(n899 ,n8[27] ,n2533);
    nor g1873(n898 ,n8[16] ,n2[112]);
    nor g1874(n897 ,n2[97] ,n10[1]);
    nor g1875(n896 ,n8[24] ,n2[120]);
    nor g1876(n895 ,n8[4] ,n2[68]);
    nor g1877(n894 ,n8[3] ,n2[99]);
    nor g1878(n893 ,n8[23] ,n2[87]);
    nor g1879(n892 ,n8[4] ,n2542);
    nor g1880(n891 ,n8[26] ,n2564);
    nor g1881(n890 ,n8[2] ,n2[66]);
    nor g1882(n889 ,n8[6] ,n2512);
    nor g1883(n888 ,n8[6] ,n2[70]);
    nor g1884(n887 ,n8[2] ,n2[98]);
    nor g1885(n886 ,n8[7] ,n2513);
    nor g1886(n885 ,n2538 ,n10[0]);
    nor g1887(n884 ,n8[18] ,n2556);
    nor g1888(n883 ,n8[9] ,n2547);
    nor g1889(n882 ,n8[14] ,n2552);
    nor g1890(n881 ,n8[21] ,n2559);
    nor g1891(n880 ,n8[13] ,n2[109]);
    nor g1892(n879 ,n8[7] ,n2[7]);
    nor g1893(n878 ,n8[2] ,n2[2]);
    nor g1894(n877 ,n8[3] ,n2509);
    nor g1895(n876 ,n8[20] ,n2558);
    nor g1896(n875 ,n8[13] ,n2551);
    nor g1897(n874 ,n8[13] ,n2[45]);
    nor g1898(n873 ,n8[17] ,n2555);
    nor g1899(n872 ,n8[31] ,n2[95]);
    nor g1900(n871 ,n8[12] ,n2550);
    nor g1901(n870 ,n8[19] ,n2557);
    nor g1902(n869 ,n8[19] ,n2[115]);
    nor g1903(n868 ,n8[3] ,n2[35]);
    nor g1904(n867 ,n8[18] ,n2[82]);
    nor g1905(n866 ,n8[30] ,n2[126]);
    nor g1906(n865 ,n8[30] ,n2568);
    nor g1907(n864 ,n8[29] ,n2567);
    nor g1908(n863 ,n8[27] ,n2565);
    nor g1909(n862 ,n8[19] ,n2[83]);
    nor g1910(n861 ,n8[11] ,n2517);
    nor g1911(n860 ,n8[11] ,n2[107]);
    nor g1912(n859 ,n8[12] ,n2518);
    nor g1913(n858 ,n8[11] ,n2549);
    nor g1914(n857 ,n8[3] ,n2541);
    nor g1915(n856 ,n8[10] ,n2[106]);
    nor g1916(n855 ,n8[17] ,n2[81]);
    nor g1917(n854 ,n8[10] ,n2[10]);
    nor g1918(n853 ,n8[11] ,n2[11]);
    nor g1919(n852 ,n8[20] ,n2[52]);
    nor g1920(n851 ,n8[26] ,n2[122]);
    nor g1921(n850 ,n8[12] ,n2[12]);
    nor g1922(n849 ,n8[4] ,n2510);
    nor g1923(n848 ,n8[13] ,n2[13]);
    nor g1924(n847 ,n8[15] ,n2521);
    nor g1925(n846 ,n8[13] ,n2519);
    nor g1926(n845 ,n8[26] ,n2[26]);
    nor g1927(n844 ,n8[9] ,n2[9]);
    nor g1928(n843 ,n8[15] ,n2[15]);
    nor g1929(n842 ,n8[21] ,n2[85]);
    nor g1930(n841 ,n8[30] ,n2[62]);
    nor g1931(n840 ,n8[16] ,n2522);
    nor g1932(n839 ,n8[31] ,n2[127]);
    nor g1933(n838 ,n8[17] ,n2[17]);
    nor g1934(n837 ,n8[25] ,n2563);
    nor g1935(n836 ,n8[28] ,n2[124]);
    nor g1936(n835 ,n8[17] ,n2523);
    nor g1937(n834 ,n8[18] ,n2[18]);
    nor g1938(n833 ,n2[32] ,n10[0]);
    nor g1939(n832 ,n8[26] ,n2532);
    nor g1940(n831 ,n8[9] ,n2[105]);
    nor g1941(n830 ,n8[20] ,n2[20]);
    nor g1942(n829 ,n8[21] ,n2[21]);
    nor g1943(n828 ,n8[29] ,n2535);
    nor g1944(n827 ,n320 ,n281);
    nor g1945(n826 ,n8[14] ,n2[14]);
    nor g1946(n825 ,n8[25] ,n2[89]);
    nor g1947(n824 ,n8[19] ,n2525);
    nor g1948(n823 ,n8[24] ,n2[24]);
    nor g1949(n822 ,n8[7] ,n2[103]);
    nor g1950(n821 ,n8[29] ,n2[93]);
    nor g1951(n820 ,n8[29] ,n2[61]);
    nor g1952(n819 ,n8[25] ,n2[25]);
    nor g1953(n818 ,n8[14] ,n2[110]);
    nor g1954(n817 ,n8[20] ,n2526);
    nor g1955(n816 ,n8[2] ,n2508);
    nor g1956(n815 ,n8[27] ,n2[27]);
    nor g1957(n814 ,n2[96] ,n10[0]);
    nor g1958(n813 ,n8[8] ,n2[104]);
    nor g1959(n812 ,n8[20] ,n2[116]);
    nor g1960(n811 ,n8[28] ,n2[28]);
    nor g1961(n810 ,n8[29] ,n2[29]);
    nor g1962(n809 ,n8[30] ,n2[30]);
    nor g1963(n808 ,n8[19] ,n2[51]);
    nor g1964(n807 ,n8[22] ,n2528);
    nor g1965(n806 ,n8[19] ,n2[19]);
    nor g1966(n805 ,n8[31] ,n2[31]);
    nor g1967(n804 ,n8[29] ,n2[125]);
    nor g1968(n803 ,n8[7] ,n2[39]);
    nor g1969(n802 ,n8[3] ,n2[67]);
    nor g1970(n801 ,n8[18] ,n2[114]);
    nor g1971(n800 ,n8[26] ,n2[90]);
    nor g1972(n799 ,n8[2] ,n2[34]);
    nor g1973(n798 ,n2[1] ,n10[1]);
    nor g1974(n797 ,n8[13] ,n2[77]);
    nor g1975(n796 ,n8[23] ,n2529);
    nor g1976(n795 ,n8[31] ,n2569);
    nor g1977(n794 ,n2[0] ,n10[0]);
    nor g1978(n793 ,n8[21] ,n2527);
    nor g1979(n792 ,n8[4] ,n2[36]);
    nor g1980(n791 ,n8[14] ,n2[78]);
    nor g1981(n790 ,n8[5] ,n2[37]);
    nor g1982(n789 ,n8[24] ,n2562);
    nor g1983(n788 ,n8[6] ,n2[38]);
    nor g1984(n787 ,n8[30] ,n2[94]);
    nor g1985(n786 ,n8[12] ,n2[76]);
    nor g1986(n785 ,n8[8] ,n2[40]);
    nor g1987(n784 ,n8[5] ,n2511);
    nor g1988(n783 ,n8[10] ,n2[42]);
    nor g1989(n782 ,n8[11] ,n2[43]);
    nor g1990(n781 ,n8[23] ,n2561);
    nor g1991(n780 ,n8[24] ,n2530);
    nor g1992(n779 ,n8[14] ,n2[46]);
    nor g1993(n778 ,n8[17] ,n2[49]);
    nor g1994(n777 ,n8[28] ,n2[60]);
    nor g1995(n776 ,n8[9] ,n2[41]);
    nor g1996(n775 ,n8[28] ,n2534);
    nor g1997(n774 ,n8[6] ,n2[102]);
    nor g1998(n773 ,n8[11] ,n2[75]);
    nor g1999(n772 ,n8[21] ,n2[117]);
    nor g2000(n771 ,n8[20] ,n2[84]);
    nor g2001(n770 ,n8[18] ,n2[50]);
    nor g2002(n769 ,n8[27] ,n2[123]);
    nor g2003(n768 ,n8[8] ,n2[72]);
    nor g2004(n767 ,n8[28] ,n2[92]);
    nor g2005(n766 ,n8[10] ,n2[74]);
    nor g2006(n765 ,n8[21] ,n2[53]);
    nor g2007(n764 ,n8[15] ,n2[47]);
    nor g2008(n763 ,n8[25] ,n2[121]);
    nor g2009(n762 ,n8[16] ,n2[48]);
    nor g2010(n761 ,n8[8] ,n2514);
    nor g2011(n760 ,n6[0] ,n288);
    nor g2012(n759 ,n8[27] ,n2[59]);
    nor g2013(n758 ,n8[23] ,n2[23]);
    nor g2014(n757 ,n8[17] ,n2[113]);
    nor g2015(n756 ,n8[8] ,n2[8]);
    nor g2016(n755 ,n2507 ,n10[1]);
    nor g2017(n754 ,n8[25] ,n2531);
    nor g2018(n753 ,n8[5] ,n2[5]);
    nor g2019(n752 ,n2[64] ,n10[0]);
    nor g2020(n751 ,n8[9] ,n2515);
    nor g2021(n750 ,n2[65] ,n10[1]);
    nor g2022(n749 ,n8[27] ,n2[91]);
    nor g2023(n748 ,n8[8] ,n2546);
    nor g2024(n747 ,n8[31] ,n2537);
    nor g2025(n746 ,n2506 ,n10[0]);
    nor g2026(n745 ,n8[28] ,n2566);
    nor g2027(n744 ,n8[16] ,n2554);
    nor g2028(n743 ,n8[10] ,n2516);
    nor g2029(n742 ,n8[31] ,n2[63]);
    nor g2030(n741 ,n8[14] ,n2520);
    nor g2031(n740 ,n8[26] ,n2[58]);
    nor g2032(n739 ,n8[6] ,n2[6]);
    nor g2033(n738 ,n8[7] ,n2545);
    nor g2034(n737 ,n8[9] ,n2[73]);
    nor g2035(n736 ,n8[3] ,n2[3]);
    nor g2036(n735 ,n8[5] ,n2[101]);
    nor g2037(n734 ,n8[22] ,n2[118]);
    nor g2038(n733 ,n8[7] ,n2[71]);
    nor g2039(n732 ,n8[22] ,n2[22]);
    nor g2040(n731 ,n8[6] ,n2544);
    nor g2041(n730 ,n8[4] ,n2[4]);
    nor g2042(n729 ,n8[25] ,n2[57]);
    nor g2043(n728 ,n8[24] ,n2[88]);
    nor g2044(n727 ,n8[24] ,n2[56]);
    nor g2045(n726 ,n8[18] ,n2524);
    nor g2046(n725 ,n8[22] ,n2[54]);
    nor g2047(n724 ,n8[10] ,n2548);
    nor g2048(n723 ,n8[16] ,n2[80]);
    nor g2049(n722 ,n8[5] ,n2[69]);
    nor g2050(n721 ,n8[16] ,n2[16]);
    nor g2051(n720 ,n8[23] ,n2[119]);
    nor g2052(n719 ,n8[30] ,n2536);
    nor g2053(n718 ,n8[5] ,n2543);
    nor g2054(n717 ,n8[15] ,n2[111]);
    nor g2055(n716 ,n8[23] ,n2[55]);
    nor g2056(n715 ,n8[15] ,n2[79]);
    or g2057(n714 ,n9[0] ,n9[1]);
    not g2058(n713 ,n6[2]);
    not g2059(n712 ,n6[3]);
    not g2060(n711 ,n6[1]);
    not g2061(n710 ,n3[13]);
    not g2062(n709 ,n5[25]);
    not g2063(n708 ,n5[53]);
    not g2064(n707 ,n4[1]);
    not g2065(n706 ,n5[49]);
    not g2066(n705 ,n3[29]);
    not g2067(n704 ,n5[56]);
    not g2068(n703 ,n4[37]);
    not g2069(n702 ,n4[53]);
    not g2070(n701 ,n3[39]);
    not g2071(n700 ,n3[60]);
    not g2072(n699 ,n4[59]);
    not g2073(n698 ,n5[51]);
    not g2074(n697 ,n5[32]);
    not g2075(n696 ,n4[5]);
    not g2076(n695 ,n5[61]);
    not g2077(n694 ,n5[30]);
    not g2078(n693 ,n4[7]);
    not g2079(n692 ,n3[62]);
    not g2080(n691 ,n4[45]);
    not g2081(n690 ,n4[21]);
    not g2082(n689 ,n3[20]);
    not g2083(n688 ,n3[1]);
    not g2084(n687 ,n3[47]);
    not g2085(n686 ,n4[44]);
    not g2086(n685 ,n5[39]);
    not g2087(n684 ,n5[48]);
    not g2088(n683 ,n4[35]);
    not g2089(n682 ,n4[28]);
    not g2090(n681 ,n5[38]);
    not g2091(n680 ,n3[53]);
    not g2092(n679 ,n5[40]);
    not g2093(n678 ,n3[19]);
    not g2094(n677 ,n3[3]);
    not g2095(n676 ,n5[50]);
    not g2096(n675 ,n3[33]);
    not g2097(n674 ,n5[54]);
    not g2098(n673 ,n4[22]);
    not g2099(n672 ,n5[42]);
    not g2100(n671 ,n3[26]);
    not g2101(n670 ,n3[51]);
    not g2102(n669 ,n3[56]);
    not g2103(n668 ,n4[31]);
    not g2104(n667 ,n3[25]);
    not g2105(n666 ,n4[12]);
    not g2106(n665 ,n4[15]);
    not g2107(n664 ,n5[45]);
    not g2108(n663 ,n5[2]);
    not g2109(n662 ,n3[48]);
    not g2110(n661 ,n3[21]);
    not g2111(n660 ,n4[6]);
    not g2112(n659 ,n4[41]);
    not g2113(n658 ,n3[4]);
    not g2114(n657 ,n5[31]);
    not g2115(n656 ,n5[59]);
    not g2116(n655 ,n4[10]);
    not g2117(n654 ,n4[27]);
    not g2118(n653 ,n4[24]);
    not g2119(n652 ,n3[9]);
    not g2120(n651 ,n5[12]);
    not g2121(n650 ,n4[63]);
    not g2122(n649 ,n4[2]);
    not g2123(n648 ,n4[20]);
    not g2124(n647 ,n4[8]);
    not g2125(n646 ,n3[49]);
    not g2126(n645 ,n5[55]);
    not g2127(n644 ,n5[58]);
    not g2128(n643 ,n3[8]);
    not g2129(n642 ,n5[23]);
    not g2130(n641 ,n3[6]);
    not g2131(n640 ,n3[7]);
    not g2132(n639 ,n5[34]);
    not g2133(n638 ,n3[28]);
    not g2134(n637 ,n5[5]);
    not g2135(n636 ,n3[34]);
    not g2136(n635 ,n5[57]);
    not g2137(n634 ,n3[44]);
    not g2138(n633 ,n3[24]);
    not g2139(n632 ,n4[0]);
    not g2140(n631 ,n3[11]);
    not g2141(n630 ,n5[11]);
    not g2142(n629 ,n5[47]);
    not g2143(n628 ,n5[20]);
    not g2144(n627 ,n3[41]);
    not g2145(n626 ,n4[57]);
    not g2146(n625 ,n5[1]);
    not g2147(n624 ,n4[13]);
    not g2148(n623 ,n3[52]);
    not g2149(n622 ,n3[17]);
    not g2150(n621 ,n4[60]);
    not g2151(n620 ,n4[42]);
    not g2152(n619 ,n3[5]);
    not g2153(n618 ,n5[6]);
    not g2154(n617 ,n3[58]);
    not g2155(n616 ,n5[28]);
    not g2156(n615 ,n3[46]);
    not g2157(n614 ,n4[19]);
    not g2158(n613 ,n3[2]);
    not g2159(n612 ,n4[40]);
    not g2160(n611 ,n5[22]);
    not g2161(n610 ,n4[48]);
    not g2162(n609 ,n4[29]);
    not g2163(n608 ,n5[60]);
    not g2164(n607 ,n5[29]);
    not g2165(n606 ,n3[18]);
    not g2166(n605 ,n3[27]);
    not g2167(n604 ,n3[50]);
    not g2168(n603 ,n4[56]);
    not g2169(n602 ,n4[16]);
    not g2170(n601 ,n3[42]);
    not g2171(n600 ,n5[16]);
    not g2172(n599 ,n4[50]);
    not g2173(n598 ,n4[26]);
    not g2174(n597 ,n4[39]);
    not g2175(n596 ,n4[9]);
    not g2176(n595 ,n3[30]);
    not g2177(n594 ,n5[13]);
    not g2178(n593 ,n5[41]);
    not g2179(n592 ,n4[51]);
    not g2180(n591 ,n4[14]);
    not g2181(n590 ,n4[38]);
    not g2182(n589 ,n6[0]);
    not g2183(n588 ,n4[62]);
    not g2184(n587 ,n3[12]);
    not g2185(n586 ,n4[43]);
    not g2186(n585 ,n3[22]);
    not g2187(n584 ,n3[16]);
    not g2188(n583 ,n3[10]);
    not g2189(n582 ,n3[38]);
    not g2190(n581 ,n3[57]);
    not g2191(n580 ,n5[26]);
    not g2192(n579 ,n4[34]);
    not g2193(n578 ,n5[15]);
    not g2194(n577 ,n5[35]);
    not g2195(n576 ,n3[15]);
    not g2196(n575 ,n3[32]);
    not g2197(n574 ,n5[52]);
    not g2198(n573 ,n4[54]);
    not g2199(n572 ,n3[40]);
    not g2200(n571 ,n3[54]);
    not g2201(n570 ,n3[55]);
    not g2202(n569 ,n5[21]);
    not g2203(n568 ,n4[30]);
    not g2204(n567 ,n3[37]);
    not g2205(n566 ,n3[14]);
    not g2206(n565 ,n3[45]);
    not g2207(n564 ,n5[19]);
    not g2208(n563 ,n5[14]);
    not g2209(n562 ,n5[63]);
    not g2210(n561 ,n3[36]);
    not g2211(n560 ,n5[36]);
    not g2212(n559 ,n5[3]);
    not g2213(n558 ,n5[33]);
    not g2214(n557 ,n5[62]);
    not g2215(n556 ,n4[32]);
    not g2216(n555 ,n4[52]);
    not g2217(n554 ,n3[31]);
    not g2218(n553 ,n3[63]);
    not g2219(n552 ,n4[46]);
    not g2220(n551 ,n3[59]);
    not g2221(n550 ,n5[8]);
    not g2222(n549 ,n4[18]);
    not g2223(n548 ,n5[7]);
    not g2224(n547 ,n4[25]);
    not g2225(n546 ,n3[23]);
    not g2226(n545 ,n3[43]);
    not g2227(n544 ,n5[4]);
    not g2228(n543 ,n3[61]);
    not g2229(n542 ,n3[0]);
    not g2230(n541 ,n9[1]);
    not g2231(n540 ,n9[0]);
    not g2232(n539 ,n8[18]);
    not g2233(n538 ,n8[3]);
    not g2234(n537 ,n8[27]);
    not g2235(n536 ,n8[22]);
    not g2236(n535 ,n8[24]);
    not g2237(n534 ,n8[17]);
    not g2238(n533 ,n8[4]);
    not g2239(n532 ,n8[21]);
    not g2240(n531 ,n8[7]);
    not g2241(n530 ,n8[28]);
    not g2242(n529 ,n8[13]);
    not g2243(n528 ,n8[25]);
    not g2244(n527 ,n8[29]);
    not g2245(n526 ,n8[10]);
    not g2246(n525 ,n8[16]);
    not g2247(n524 ,n8[20]);
    not g2248(n523 ,n8[30]);
    not g2249(n522 ,n8[11]);
    not g2250(n521 ,n8[6]);
    not g2251(n520 ,n8[9]);
    not g2252(n519 ,n8[2]);
    not g2253(n518 ,n8[23]);
    not g2254(n517 ,n8[26]);
    not g2255(n516 ,n8[12]);
    not g2256(n515 ,n8[15]);
    not g2257(n514 ,n8[8]);
    not g2258(n513 ,n8[19]);
    not g2259(n512 ,n2571);
    not g2260(n511 ,n2572);
    not g2261(n510 ,n2570);
    not g2262(n509 ,n2528);
    not g2263(n508 ,n2[100]);
    not g2264(n507 ,n2[125]);
    not g2265(n506 ,n2532);
    not g2266(n505 ,n2[99]);
    not g2267(n504 ,n2561);
    not g2268(n503 ,n2565);
    not g2269(n502 ,n2[88]);
    not g2270(n501 ,n2510);
    not g2271(n500 ,n2543);
    not g2272(n499 ,n2[113]);
    not g2273(n498 ,n2[72]);
    not g2274(n497 ,n2[85]);
    not g2275(n496 ,n2[124]);
    not g2276(n495 ,n2[117]);
    not g2277(n494 ,n2[101]);
    not g2278(n493 ,n2534);
    not g2279(n492 ,n2[112]);
    not g2280(n491 ,n2554);
    not g2281(n490 ,n2[94]);
    not g2282(n489 ,n2553);
    not g2283(n488 ,n2[109]);
    not g2284(n487 ,n2[102]);
    not g2285(n486 ,n2[82]);
    not g2286(n485 ,n2559);
    not g2287(n484 ,n2[80]);
    not g2288(n483 ,n2[69]);
    not g2289(n482 ,n2[126]);
    not g2290(n481 ,n2531);
    not g2291(n480 ,n2[98]);
    not g2292(n479 ,n2[107]);
    not g2293(n478 ,n2[104]);
    not g2294(n477 ,n2517);
    not g2295(n476 ,n2[75]);
    not g2296(n475 ,n2514);
    not g2297(n474 ,n2[105]);
    not g2298(n473 ,n2533);
    not g2299(n472 ,n2[89]);
    not g2300(n471 ,n2[115]);
    not g2301(n470 ,n2535);
    not g2302(n469 ,n2545);
    not g2303(n468 ,n2[86]);
    not g2304(n467 ,n2[108]);
    not g2305(n466 ,n2549);
    not g2306(n465 ,n2[110]);
    not g2307(n464 ,n2521);
    not g2308(n463 ,n2[95]);
    not g2309(n462 ,n2527);
    not g2310(n461 ,n2564);
    not g2311(n460 ,n2[64]);
    not g2312(n459 ,n2[111]);
    not g2313(n458 ,n2518);
    not g2314(n457 ,n2569);
    not g2315(n456 ,n2546);
    not g2316(n455 ,n2552);
    not g2317(n454 ,n2526);
    not g2318(n453 ,n2[123]);
    not g2319(n452 ,n2522);
    not g2320(n451 ,n2[78]);
    not g2321(n450 ,n2[87]);
    not g2322(n449 ,n2[127]);
    not g2323(n448 ,n2[84]);
    not g2324(n447 ,n2[83]);
    not g2325(n446 ,n2[65]);
    not g2326(n445 ,n2[90]);
    not g2327(n444 ,n2513);
    not g2328(n443 ,n2[103]);
    not g2329(n442 ,n2512);
    not g2330(n441 ,n2507);
    not g2331(n440 ,n2[122]);
    not g2332(n439 ,n2506);
    not g2333(n438 ,n2[114]);
    not g2334(n437 ,n2560);
    not g2335(n436 ,n2[79]);
    not g2336(n435 ,n2536);
    not g2337(n434 ,n2[119]);
    not g2338(n433 ,n2516);
    not g2339(n432 ,n2508);
    not g2340(n431 ,n2547);
    not g2341(n430 ,n2[70]);
    not g2342(n429 ,n2511);
    not g2343(n428 ,n2523);
    not g2344(n427 ,n2520);
    not g2345(n426 ,n2[116]);
    not g2346(n425 ,n2[66]);
    not g2347(n424 ,n2[96]);
    not g2348(n423 ,n2557);
    not g2349(n422 ,n2567);
    not g2350(n421 ,n2[93]);
    not g2351(n420 ,n2[118]);
    not g2352(n419 ,n2541);
    not g2353(n418 ,n2538);
    not g2354(n417 ,n2558);
    not g2355(n416 ,n2568);
    not g2356(n415 ,n2[76]);
    not g2357(n414 ,n2551);
    not g2358(n413 ,n2566);
    not g2359(n412 ,n2[73]);
    not g2360(n411 ,n2548);
    not g2361(n410 ,n2542);
    not g2362(n409 ,n2[67]);
    not g2363(n408 ,n2[68]);
    not g2364(n407 ,n2562);
    not g2365(n406 ,n2524);
    not g2366(n405 ,n2[91]);
    not g2367(n404 ,n2515);
    not g2368(n403 ,n2[81]);
    not g2369(n402 ,n2544);
    not g2370(n401 ,n2[77]);
    not g2371(n400 ,n2525);
    not g2372(n399 ,n2555);
    not g2373(n398 ,n2519);
    not g2374(n397 ,n2540);
    not g2375(n396 ,n2[121]);
    not g2376(n395 ,n2537);
    not g2377(n394 ,n2509);
    not g2378(n393 ,n2[71]);
    not g2379(n392 ,n2[97]);
    not g2380(n391 ,n2556);
    not g2381(n390 ,n2530);
    not g2382(n389 ,n2529);
    not g2383(n388 ,n2[74]);
    not g2384(n387 ,n2[120]);
    not g2385(n386 ,n2550);
    not g2386(n385 ,n2539);
    not g2387(n384 ,n2563);
    not g2388(n383 ,n2[92]);
    not g2389(n382 ,n2[106]);
    not g2390(n381 ,n2[25]);
    not g2391(n380 ,n2[54]);
    not g2392(n379 ,n4[55]);
    not g2393(n378 ,n2[20]);
    not g2394(n377 ,n5[17]);
    not g2395(n376 ,n5[37]);
    not g2396(n375 ,n4[61]);
    not g2397(n374 ,n4[47]);
    not g2398(n373 ,n5[46]);
    not g2399(n372 ,n2[32]);
    not g2400(n371 ,n2[6]);
    not g2401(n370 ,n2[56]);
    not g2402(n369 ,n2[14]);
    not g2403(n368 ,n2[7]);
    not g2404(n367 ,n2[4]);
    not g2405(n366 ,n2[45]);
    not g2406(n365 ,n2[35]);
    not g2407(n364 ,n2[51]);
    not g2408(n363 ,n2[11]);
    not g2409(n362 ,n4[36]);
    not g2410(n361 ,n2[30]);
    not g2411(n360 ,n2[24]);
    not g2412(n359 ,n2[49]);
    not g2413(n358 ,n2[15]);
    not g2414(n357 ,n2[41]);
    not g2415(n356 ,n2[33]);
    not g2416(n355 ,n2[9]);
    not g2417(n354 ,n2[31]);
    not g2418(n353 ,n3[35]);
    not g2419(n352 ,n4[58]);
    not g2420(n351 ,n4[17]);
    not g2421(n350 ,n4[33]);
    not g2422(n349 ,n2[5]);
    not g2423(n348 ,n2[42]);
    not g2424(n347 ,n2[39]);
    not g2425(n346 ,n2[63]);
    not g2426(n345 ,n2[57]);
    not g2427(n344 ,n2[23]);
    not g2428(n343 ,n5[24]);
    not g2429(n342 ,n2[16]);
    not g2430(n341 ,n5[9]);
    not g2431(n340 ,n5[44]);
    not g2432(n339 ,n2[55]);
    not g2433(n338 ,n4[11]);
    not g2434(n337 ,n2[28]);
    not g2435(n336 ,n2[62]);
    not g2436(n335 ,n4[49]);
    not g2437(n334 ,n5[27]);
    not g2438(n333 ,n2[44]);
    not g2439(n332 ,n2[2]);
    not g2440(n331 ,n2[53]);
    not g2441(n330 ,n4[3]);
    not g2442(n329 ,n5[18]);
    not g2443(n328 ,n2[40]);
    not g2444(n327 ,n4[23]);
    not g2445(n326 ,n2[10]);
    not g2446(n325 ,n2[22]);
    not g2447(n324 ,n2[29]);
    not g2448(n323 ,n5[0]);
    not g2449(n322 ,n2[3]);
    not g2450(n321 ,n2[48]);
    not g2451(n320 ,n2[34]);
    not g2452(n319 ,n2[37]);
    not g2453(n318 ,n2[61]);
    not g2454(n317 ,n2[38]);
    not g2455(n316 ,n2[58]);
    not g2456(n315 ,n2[59]);
    not g2457(n314 ,n2[1]);
    not g2458(n313 ,n2[0]);
    not g2459(n312 ,n5[43]);
    not g2460(n311 ,n2[52]);
    not g2461(n310 ,n2[13]);
    not g2462(n309 ,n2[60]);
    not g2463(n308 ,n2[12]);
    not g2464(n307 ,n2[46]);
    not g2465(n306 ,n4[4]);
    not g2466(n305 ,n2[47]);
    not g2467(n304 ,n2[43]);
    not g2468(n303 ,n5[10]);
    not g2469(n302 ,n2[50]);
    not g2470(n301 ,n2[19]);
    not g2471(n300 ,n2[17]);
    not g2472(n299 ,n2[18]);
    not g2473(n298 ,n2[26]);
    not g2474(n297 ,n2[21]);
    not g2475(n296 ,n2[27]);
    not g2476(n295 ,n2[8]);
    not g2477(n294 ,n2[36]);
    not g2478(n293 ,n8[31]);
    not g2479(n292 ,n10[0]);
    not g2480(n291 ,n8[14]);
    not g2481(n290 ,n10[1]);
    not g2482(n289 ,n8[5]);
    not g2483(n288 ,n2505);
    not g2484(n287 ,n2505);
    not g2485(n286 ,n2505);
    not g2486(n285 ,n2505);
    not g2487(n284 ,n2505);
    not g2488(n283 ,n2505);
    not g2489(n282 ,n2505);
    not g2490(n281 ,n2505);
    not g2491(n280 ,n2505);
    xnor g2492(n2569 ,n79 ,n267);
    nor g2493(n267 ,n52 ,n266);
    xnor g2494(n2568 ,n95 ,n265);
    nor g2495(n266 ,n95 ,n265);
    nor g2496(n265 ,n41 ,n264);
    xnor g2497(n2567 ,n116 ,n263);
    nor g2498(n264 ,n116 ,n263);
    nor g2499(n263 ,n70 ,n262);
    xnor g2500(n2566 ,n98 ,n261);
    nor g2501(n262 ,n98 ,n261);
    nor g2502(n261 ,n44 ,n260);
    xnor g2503(n2565 ,n103 ,n259);
    nor g2504(n260 ,n103 ,n259);
    nor g2505(n259 ,n56 ,n258);
    xnor g2506(n2564 ,n125 ,n257);
    nor g2507(n258 ,n125 ,n257);
    nor g2508(n257 ,n37 ,n256);
    xnor g2509(n2563 ,n108 ,n255);
    nor g2510(n256 ,n108 ,n255);
    nor g2511(n255 ,n71 ,n254);
    xnor g2512(n2562 ,n97 ,n253);
    nor g2513(n254 ,n97 ,n253);
    nor g2514(n253 ,n17 ,n252);
    xnor g2515(n2561 ,n136 ,n251);
    nor g2516(n252 ,n136 ,n251);
    nor g2517(n251 ,n36 ,n250);
    xnor g2518(n2560 ,n90 ,n249);
    nor g2519(n250 ,n90 ,n249);
    nor g2520(n249 ,n63 ,n248);
    xnor g2521(n2559 ,n131 ,n247);
    nor g2522(n248 ,n131 ,n247);
    nor g2523(n247 ,n48 ,n246);
    xnor g2524(n2558 ,n126 ,n245);
    nor g2525(n246 ,n126 ,n245);
    nor g2526(n245 ,n40 ,n244);
    xnor g2527(n2557 ,n120 ,n243);
    nor g2528(n244 ,n120 ,n243);
    nor g2529(n243 ,n32 ,n242);
    xnor g2530(n2556 ,n112 ,n241);
    nor g2531(n242 ,n112 ,n241);
    nor g2532(n241 ,n28 ,n240);
    xnor g2533(n2555 ,n101 ,n239);
    nor g2534(n240 ,n101 ,n239);
    nor g2535(n239 ,n22 ,n238);
    xnor g2536(n2554 ,n110 ,n237);
    nor g2537(n238 ,n110 ,n237);
    nor g2538(n237 ,n15 ,n236);
    xnor g2539(n2553 ,n86 ,n235);
    nor g2540(n236 ,n86 ,n235);
    nor g2541(n235 ,n58 ,n234);
    xnor g2542(n2552 ,n81 ,n233);
    nor g2543(n234 ,n81 ,n233);
    nor g2544(n233 ,n76 ,n232);
    xnor g2545(n2551 ,n83 ,n231);
    nor g2546(n232 ,n83 ,n231);
    nor g2547(n231 ,n57 ,n230);
    xnor g2548(n2550 ,n89 ,n229);
    nor g2549(n230 ,n89 ,n229);
    nor g2550(n229 ,n64 ,n228);
    xnor g2551(n2549 ,n138 ,n227);
    nor g2552(n228 ,n138 ,n227);
    nor g2553(n227 ,n31 ,n226);
    xnor g2554(n2548 ,n134 ,n225);
    nor g2555(n226 ,n134 ,n225);
    nor g2556(n225 ,n50 ,n224);
    xnor g2557(n2547 ,n129 ,n223);
    nor g2558(n224 ,n129 ,n223);
    nor g2559(n223 ,n26 ,n222);
    xnor g2560(n2546 ,n99 ,n221);
    nor g2561(n222 ,n99 ,n221);
    nor g2562(n221 ,n42 ,n220);
    xnor g2563(n2545 ,n123 ,n219);
    nor g2564(n220 ,n123 ,n219);
    nor g2565(n219 ,n67 ,n218);
    xnor g2566(n2544 ,n119 ,n217);
    nor g2567(n218 ,n119 ,n217);
    nor g2568(n217 ,n34 ,n216);
    xnor g2569(n2543 ,n114 ,n215);
    nor g2570(n216 ,n114 ,n215);
    nor g2571(n215 ,n39 ,n214);
    xnor g2572(n2542 ,n111 ,n213);
    nor g2573(n214 ,n111 ,n213);
    nor g2574(n213 ,n54 ,n212);
    xnor g2575(n2541 ,n109 ,n211);
    nor g2576(n212 ,n109 ,n211);
    nor g2577(n211 ,n18 ,n210);
    xnor g2578(n2540 ,n105 ,n209);
    nor g2579(n210 ,n105 ,n209);
    nor g2580(n209 ,n24 ,n208);
    xnor g2581(n2539 ,n100 ,n207);
    nor g2582(n208 ,n100 ,n207);
    nor g2583(n207 ,n47 ,n206);
    xnor g2584(n2538 ,n93 ,n205);
    nor g2585(n206 ,n93 ,n205);
    nor g2586(n205 ,n73 ,n204);
    xnor g2587(n2537 ,n88 ,n203);
    nor g2588(n204 ,n88 ,n203);
    nor g2589(n203 ,n74 ,n202);
    xnor g2590(n2536 ,n85 ,n201);
    nor g2591(n202 ,n85 ,n201);
    nor g2592(n201 ,n16 ,n200);
    xnor g2593(n2535 ,n80 ,n199);
    nor g2594(n200 ,n80 ,n199);
    nor g2595(n199 ,n53 ,n198);
    xnor g2596(n2534 ,n82 ,n197);
    nor g2597(n198 ,n82 ,n197);
    nor g2598(n197 ,n68 ,n196);
    xnor g2599(n2533 ,n84 ,n195);
    nor g2600(n196 ,n84 ,n195);
    nor g2601(n195 ,n65 ,n194);
    xnor g2602(n2532 ,n87 ,n193);
    nor g2603(n194 ,n87 ,n193);
    nor g2604(n193 ,n45 ,n192);
    xnor g2605(n2531 ,n92 ,n191);
    nor g2606(n192 ,n92 ,n191);
    nor g2607(n191 ,n43 ,n190);
    xnor g2608(n2530 ,n91 ,n189);
    nor g2609(n190 ,n91 ,n189);
    nor g2610(n189 ,n19 ,n188);
    xnor g2611(n2529 ,n140 ,n187);
    nor g2612(n188 ,n140 ,n187);
    nor g2613(n187 ,n62 ,n186);
    xnor g2614(n2528 ,n137 ,n185);
    nor g2615(n186 ,n137 ,n185);
    nor g2616(n185 ,n59 ,n184);
    xnor g2617(n2527 ,n135 ,n183);
    nor g2618(n184 ,n135 ,n183);
    nor g2619(n183 ,n55 ,n182);
    xnor g2620(n2526 ,n133 ,n181);
    nor g2621(n182 ,n133 ,n181);
    nor g2622(n181 ,n51 ,n180);
    xnor g2623(n2525 ,n132 ,n179);
    nor g2624(n180 ,n132 ,n179);
    nor g2625(n179 ,n49 ,n178);
    xnor g2626(n2524 ,n130 ,n177);
    nor g2627(n178 ,n130 ,n177);
    nor g2628(n177 ,n30 ,n176);
    xnor g2629(n2523 ,n127 ,n175);
    nor g2630(n176 ,n127 ,n175);
    nor g2631(n175 ,n21 ,n174);
    xnor g2632(n2522 ,n106 ,n173);
    nor g2633(n174 ,n106 ,n173);
    nor g2634(n173 ,n23 ,n172);
    xnor g2635(n2521 ,n124 ,n171);
    nor g2636(n172 ,n124 ,n171);
    nor g2637(n171 ,n66 ,n170);
    xnor g2638(n2520 ,n122 ,n169);
    nor g2639(n170 ,n122 ,n169);
    nor g2640(n169 ,n38 ,n168);
    xnor g2641(n2519 ,n121 ,n167);
    nor g2642(n168 ,n121 ,n167);
    nor g2643(n167 ,n35 ,n166);
    xnor g2644(n2518 ,n118 ,n165);
    nor g2645(n166 ,n118 ,n165);
    nor g2646(n165 ,n69 ,n164);
    xnor g2647(n2517 ,n117 ,n163);
    nor g2648(n164 ,n117 ,n163);
    nor g2649(n163 ,n33 ,n162);
    xnor g2650(n2516 ,n115 ,n161);
    nor g2651(n162 ,n115 ,n161);
    nor g2652(n161 ,n46 ,n160);
    xnor g2653(n2515 ,n113 ,n159);
    nor g2654(n160 ,n113 ,n159);
    nor g2655(n159 ,n29 ,n158);
    xnor g2656(n2514 ,n128 ,n157);
    nor g2657(n158 ,n128 ,n157);
    nor g2658(n157 ,n60 ,n156);
    xnor g2659(n2513 ,n94 ,n155);
    nor g2660(n156 ,n94 ,n155);
    nor g2661(n155 ,n27 ,n154);
    xnor g2662(n2512 ,n139 ,n153);
    nor g2663(n154 ,n139 ,n153);
    nor g2664(n153 ,n25 ,n152);
    xnor g2665(n2511 ,n107 ,n151);
    nor g2666(n152 ,n107 ,n151);
    nor g2667(n151 ,n75 ,n150);
    xnor g2668(n2510 ,n104 ,n149);
    nor g2669(n150 ,n104 ,n149);
    nor g2670(n149 ,n72 ,n148);
    xor g2671(n2509 ,n102 ,n146);
    nor g2672(n148 ,n102 ,n147);
    not g2673(n147 ,n146);
    nor g2674(n146 ,n61 ,n145);
    xnor g2675(n2508 ,n141 ,n143);
    nor g2676(n145 ,n141 ,n144);
    not g2677(n144 ,n143);
    nor g2678(n143 ,n20 ,n142);
    xnor g2679(n2507 ,n96 ,n78);
    nor g2680(n142 ,n78 ,n96);
    nor g2681(n2506 ,n78 ,n77);
    xnor g2682(n141 ,n2[2] ,n2[66]);
    xnor g2683(n140 ,n2[23] ,n2[87]);
    xnor g2684(n139 ,n2[6] ,n2[70]);
    xnor g2685(n138 ,n2[43] ,n2[107]);
    xnor g2686(n137 ,n2[22] ,n2[86]);
    xnor g2687(n136 ,n2[55] ,n2[119]);
    xnor g2688(n135 ,n2[21] ,n2[85]);
    xnor g2689(n134 ,n2[42] ,n2[106]);
    xnor g2690(n133 ,n2[20] ,n2[84]);
    xnor g2691(n132 ,n2[19] ,n2[83]);
    xnor g2692(n131 ,n2[53] ,n2[117]);
    xnor g2693(n130 ,n2[18] ,n2[82]);
    xnor g2694(n129 ,n2[41] ,n2[105]);
    xnor g2695(n128 ,n2[8] ,n2[72]);
    xnor g2696(n127 ,n2[17] ,n2[81]);
    xnor g2697(n126 ,n2[52] ,n2[116]);
    xnor g2698(n125 ,n2[58] ,n2[122]);
    xnor g2699(n124 ,n2[15] ,n2[79]);
    xnor g2700(n123 ,n2[39] ,n2[103]);
    xnor g2701(n122 ,n2[14] ,n2[78]);
    xnor g2702(n121 ,n2[13] ,n2[77]);
    xnor g2703(n120 ,n2[51] ,n2[115]);
    xnor g2704(n119 ,n2[38] ,n2[102]);
    xnor g2705(n118 ,n2[12] ,n2[76]);
    xnor g2706(n117 ,n2[11] ,n2[75]);
    xnor g2707(n116 ,n2[61] ,n2[125]);
    xnor g2708(n115 ,n2[10] ,n2[74]);
    xnor g2709(n114 ,n2[37] ,n2[101]);
    xnor g2710(n113 ,n2[9] ,n2[73]);
    xnor g2711(n112 ,n2[50] ,n2[114]);
    xnor g2712(n111 ,n2[36] ,n2[100]);
    xnor g2713(n110 ,n2[48] ,n2[112]);
    xnor g2714(n109 ,n2[35] ,n2[99]);
    xnor g2715(n108 ,n2[57] ,n2[121]);
    xnor g2716(n107 ,n2[5] ,n2[69]);
    xnor g2717(n106 ,n2[16] ,n2[80]);
    xnor g2718(n105 ,n2[34] ,n2[98]);
    xnor g2719(n104 ,n2[4] ,n2[68]);
    xnor g2720(n103 ,n2[59] ,n2[123]);
    xnor g2721(n102 ,n2[3] ,n2[67]);
    xnor g2722(n101 ,n2[49] ,n2[113]);
    xnor g2723(n100 ,n2[33] ,n2[97]);
    xnor g2724(n99 ,n2[40] ,n2[104]);
    xnor g2725(n98 ,n2[60] ,n2[124]);
    xnor g2726(n97 ,n2[56] ,n2[120]);
    xnor g2727(n96 ,n2[1] ,n2[65]);
    xnor g2728(n95 ,n2[62] ,n2[126]);
    xnor g2729(n94 ,n2[7] ,n2[71]);
    xnor g2730(n93 ,n2[32] ,n2[96]);
    xnor g2731(n92 ,n2[25] ,n2[89]);
    xnor g2732(n91 ,n2[24] ,n2[88]);
    xnor g2733(n90 ,n2[54] ,n2[118]);
    xnor g2734(n89 ,n2[44] ,n2[108]);
    xnor g2735(n88 ,n2[31] ,n2[95]);
    xnor g2736(n87 ,n2[26] ,n2[90]);
    xnor g2737(n86 ,n2[47] ,n2[111]);
    xnor g2738(n85 ,n2[30] ,n2[94]);
    xnor g2739(n84 ,n2[27] ,n2[91]);
    xnor g2740(n83 ,n2[45] ,n2[109]);
    xnor g2741(n82 ,n2[28] ,n2[92]);
    xnor g2742(n81 ,n2[46] ,n2[110]);
    xnor g2743(n80 ,n2[29] ,n2[93]);
    xnor g2744(n79 ,n2[63] ,n2[127]);
    nor g2745(n77 ,n2[0] ,n2[64]);
    nor g2746(n76 ,n2[45] ,n2[109]);
    nor g2747(n75 ,n2[4] ,n2[68]);
    nor g2748(n74 ,n2[30] ,n2[94]);
    nor g2749(n73 ,n2[31] ,n2[95]);
    nor g2750(n72 ,n2[3] ,n2[67]);
    nor g2751(n71 ,n2[56] ,n2[120]);
    nor g2752(n70 ,n2[60] ,n2[124]);
    nor g2753(n69 ,n2[11] ,n2[75]);
    nor g2754(n68 ,n2[27] ,n2[91]);
    nor g2755(n67 ,n2[38] ,n2[102]);
    nor g2756(n66 ,n2[14] ,n2[78]);
    nor g2757(n65 ,n2[26] ,n2[90]);
    nor g2758(n64 ,n2[43] ,n2[107]);
    nor g2759(n63 ,n2[53] ,n2[117]);
    nor g2760(n62 ,n2[22] ,n2[86]);
    nor g2761(n61 ,n13 ,n12);
    nor g2762(n60 ,n2[7] ,n2[71]);
    nor g2763(n59 ,n2[21] ,n2[85]);
    nor g2764(n58 ,n2[46] ,n2[110]);
    nor g2765(n57 ,n2[44] ,n2[108]);
    nor g2766(n56 ,n2[58] ,n2[122]);
    nor g2767(n55 ,n2[20] ,n2[84]);
    nor g2768(n54 ,n2[35] ,n2[99]);
    nor g2769(n53 ,n2[28] ,n2[92]);
    nor g2770(n52 ,n2[62] ,n2[126]);
    nor g2771(n51 ,n2[19] ,n2[83]);
    nor g2772(n50 ,n2[41] ,n2[105]);
    nor g2773(n49 ,n2[18] ,n2[82]);
    nor g2774(n48 ,n2[52] ,n2[116]);
    nor g2775(n47 ,n2[32] ,n2[96]);
    nor g2776(n78 ,n14 ,n11);
    nor g2777(n46 ,n2[9] ,n2[73]);
    nor g2778(n45 ,n2[25] ,n2[89]);
    nor g2779(n44 ,n2[59] ,n2[123]);
    nor g2780(n43 ,n2[24] ,n2[88]);
    nor g2781(n42 ,n2[39] ,n2[103]);
    nor g2782(n41 ,n2[61] ,n2[125]);
    nor g2783(n40 ,n2[51] ,n2[115]);
    nor g2784(n39 ,n2[36] ,n2[100]);
    nor g2785(n38 ,n2[13] ,n2[77]);
    nor g2786(n37 ,n2[57] ,n2[121]);
    nor g2787(n36 ,n2[54] ,n2[118]);
    nor g2788(n35 ,n2[12] ,n2[76]);
    nor g2789(n34 ,n2[37] ,n2[101]);
    nor g2790(n33 ,n2[10] ,n2[74]);
    nor g2791(n32 ,n2[50] ,n2[114]);
    nor g2792(n31 ,n2[42] ,n2[106]);
    nor g2793(n30 ,n2[17] ,n2[81]);
    nor g2794(n29 ,n2[8] ,n2[72]);
    nor g2795(n28 ,n2[49] ,n2[113]);
    nor g2796(n27 ,n2[6] ,n2[70]);
    nor g2797(n26 ,n2[40] ,n2[104]);
    nor g2798(n25 ,n2[5] ,n2[69]);
    nor g2799(n24 ,n2[33] ,n2[97]);
    nor g2800(n23 ,n2[15] ,n2[79]);
    nor g2801(n22 ,n2[48] ,n2[112]);
    nor g2802(n21 ,n2[16] ,n2[80]);
    nor g2803(n20 ,n2[1] ,n2[65]);
    nor g2804(n19 ,n2[23] ,n2[87]);
    nor g2805(n18 ,n2[34] ,n2[98]);
    nor g2806(n17 ,n2[55] ,n2[119]);
    nor g2807(n16 ,n2[29] ,n2[93]);
    nor g2808(n15 ,n2[47] ,n2[111]);
    not g2809(n14 ,n2[0]);
    not g2810(n13 ,n2[2]);
    not g2811(n12 ,n2[66]);
    not g2812(n11 ,n2[64]);
    xor g2813(n2570 ,n6[3] ,n275);
    nor g2814(n2571 ,n274 ,n275);
    nor g2815(n275 ,n270 ,n273);
    nor g2816(n274 ,n6[2] ,n272);
    nor g2817(n2572 ,n272 ,n271);
    not g2818(n273 ,n272);
    nor g2819(n272 ,n268 ,n269);
    nor g2820(n271 ,n6[1] ,n6[0]);
    not g2821(n270 ,n6[2]);
    not g2822(n269 ,n6[0]);
    not g2823(n268 ,n6[1]);
    or g2824(n10[1] ,n8[1] ,n2616);
    or g2825(n10[0] ,n8[0] ,n2616);
    nor g2826(n2616 ,n2611 ,n2615);
    or g2827(n2615 ,n2608 ,n2614);
    or g2828(n2614 ,n2605 ,n2613);
    or g2829(n2613 ,n2612 ,n2610);
    or g2830(n2612 ,n2607 ,n2609);
    or g2831(n2611 ,n2604 ,n2606);
    or g2832(n2610 ,n2603 ,n2602);
    or g2833(n2609 ,n2595 ,n2588);
    or g2834(n2608 ,n2596 ,n2594);
    or g2835(n2607 ,n2597 ,n2601);
    or g2836(n2606 ,n2587 ,n2590);
    or g2837(n2605 ,n2591 ,n2599);
    or g2838(n2604 ,n2592 ,n2598);
    or g2839(n2603 ,n2600 ,n2589);
    or g2840(n2602 ,n2586 ,n2593);
    or g2841(n2601 ,n2576 ,n7[6]);
    or g2842(n2600 ,n2583 ,n2582);
    or g2843(n2599 ,n2585 ,n7[24]);
    or g2844(n2598 ,n2579 ,n7[17]);
    or g2845(n2597 ,n2573 ,n2574);
    or g2846(n2596 ,n2577 ,n7[22]);
    or g2847(n2595 ,n2575 ,n7[2]);
    or g2848(n2594 ,n2580 ,n7[20]);
    or g2849(n2593 ,n7[9] ,n7[8]);
    or g2850(n2592 ,n2581 ,n7[18]);
    or g2851(n2591 ,n2584 ,n7[26]);
    or g2852(n2590 ,n7[29] ,n7[28]);
    or g2853(n2589 ,n2578 ,n7[15]);
    or g2854(n2588 ,n7[1] ,n7[0]);
    or g2855(n2587 ,n7[31] ,n7[30]);
    or g2856(n2586 ,n7[11] ,n7[10]);
    not g2857(n2585 ,n7[25]);
    not g2858(n2584 ,n7[27]);
    not g2859(n2583 ,n7[13]);
    not g2860(n2582 ,n7[12]);
    not g2861(n2581 ,n7[19]);
    not g2862(n2580 ,n7[21]);
    not g2863(n2579 ,n7[16]);
    not g2864(n2578 ,n7[14]);
    not g2865(n2577 ,n7[23]);
    not g2866(n2576 ,n7[7]);
    not g2867(n2575 ,n7[3]);
    not g2868(n2574 ,n7[4]);
    not g2869(n2573 ,n7[5]);
endmodule
