module top(n0, n1, n7, n8, n9, n2, n3, n4, n5, n14, n15, n6, n16, n17, n10, n11, n12, n13);
    input n0, n1, n2, n3, n4, n5, n6;
    input [6:0] n7;
    input [7:0] n8;
    output [7:0] n9, n10, n11, n12, n13;
    output n14, n15, n16, n17;
    wire n0, n1, n2, n3, n4, n5, n6;
    wire [6:0] n7;
    wire [7:0] n8;
    wire [7:0] n9, n10, n11, n12, n13;
    wire n14, n15, n16, n17;
    wire [3:0] n18;
    wire [15:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [4:0] n22;
    wire [3:0] n23;
    wire [3:0] n24;
    wire [7:0] n25;
    wire [2:0] n26;
    wire [4:0] n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738;
    buf g0(n27[4], 1'b0);
    buf g1(n27[3], 1'b0);
    buf g2(n27[2], 1'b0);
    buf g3(n27[1], 1'b0);
    buf g4(n27[0], 1'b0);
    buf g5(n23[3], 1'b0);
    buf g6(n13[0], n10[0]);
    buf g7(n13[1], n10[1]);
    buf g8(n13[2], n10[0]);
    buf g9(n13[3], n10[1]);
    buf g10(n13[4], 1'b0);
    buf g11(n13[5], n10[7]);
    buf g12(n12[0], n11[0]);
    buf g13(n12[1], n11[1]);
    buf g14(n12[2], n11[2]);
    buf g15(n12[3], 1'b0);
    buf g16(n12[4], 1'b0);
    buf g17(n12[5], 1'b0);
    buf g18(n12[6], 1'b0);
    buf g19(n12[7], 1'b0);
    buf g20(n11[3], 1'b0);
    buf g21(n11[4], 1'b0);
    buf g22(n11[5], 1'b0);
    buf g23(n11[6], 1'b0);
    buf g24(n11[7], 1'b0);
    buf g25(n10[6], 1'b0);
    buf g26(n17, 1'b0);
    not g27(n698 ,n1);
    not g28(n697 ,n5);
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n686), .Q(n18[0]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n687), .Q(n18[1]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n684), .Q(n18[2]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n685), .Q(n18[3]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n437), .Q(n16));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n480), .Q(n19[0]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n514), .Q(n19[1]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n513), .Q(n19[2]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n512), .Q(n19[3]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n511), .Q(n19[4]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n510), .Q(n19[5]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n509), .Q(n19[6]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n508), .Q(n19[7]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n507), .Q(n19[8]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n506), .Q(n19[9]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n505), .Q(n19[10]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n504), .Q(n19[11]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n503), .Q(n19[12]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n515), .Q(n19[13]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n523), .Q(n19[14]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n502), .Q(n19[15]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n300), .Q(n10[0]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n301), .Q(n10[1]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n302), .Q(n10[7]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n269), .Q(n13[6]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n277), .Q(n13[7]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n604), .Q(n11[0]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n658), .Q(n11[1]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n448), .Q(n11[2]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n468), .Q(n9[0]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n469), .Q(n9[1]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n470), .Q(n9[2]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n457), .Q(n9[3]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n455), .Q(n9[4]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n460), .Q(n9[5]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n459), .Q(n9[6]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n458), .Q(n9[7]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n695), .Q(n20[0]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n696), .Q(n20[1]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n694), .Q(n20[2]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n693), .Q(n20[3]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n692), .Q(n20[4]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n691), .Q(n20[5]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n690), .Q(n20[6]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n689), .Q(n20[7]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n641), .Q(n21[0]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n640), .Q(n21[1]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n639), .Q(n21[2]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n638), .Q(n21[3]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n637), .Q(n21[4]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n636), .Q(n21[5]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n635), .Q(n21[6]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n634), .Q(n21[7]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n665), .Q(n22[0]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n379), .Q(n22[0]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n642), .Q(n22[1]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n378), .Q(n22[1]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n650), .Q(n22[2]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n377), .Q(n22[2]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n649), .Q(n22[3]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n376), .Q(n22[3]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n648), .Q(n22[4]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n375), .Q(n22[4]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n452), .Q(n23[3]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n647), .Q(n24[0]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n646), .Q(n24[1]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n645), .Q(n24[2]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n644), .Q(n24[3]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n666), .Q(n25[0]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n656), .Q(n25[1]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n653), .Q(n25[2]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n655), .Q(n25[3]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n654), .Q(n25[4]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n652), .Q(n25[5]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n657), .Q(n25[6]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n661), .Q(n25[7]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n548), .Q(n14));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n607), .Q(n15));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n643), .Q(n26[0]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n660), .Q(n26[1]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n651), .Q(n26[2]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n444), .Q(n10[2]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n445), .Q(n10[3]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n446), .Q(n10[4]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n447), .Q(n10[5]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n427), .Q(n27[0]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n441), .Q(n27[1]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n440), .Q(n27[2]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n439), .Q(n27[3]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n438), .Q(n27[4]));
    or g119(n696 ,n674 ,n682);
    or g120(n695 ,n675 ,n683);
    or g121(n694 ,n673 ,n681);
    or g122(n693 ,n672 ,n679);
    or g123(n692 ,n671 ,n680);
    or g124(n691 ,n670 ,n678);
    or g125(n690 ,n669 ,n677);
    or g126(n689 ,n676 ,n688);
    nor g127(n688 ,n141 ,n667);
    or g128(n687 ,n554 ,n664);
    or g129(n686 ,n553 ,n659);
    or g130(n685 ,n589 ,n662);
    or g131(n684 ,n552 ,n663);
    nor g132(n683 ,n201 ,n667);
    nor g133(n682 ,n198 ,n667);
    nor g134(n681 ,n205 ,n667);
    nor g135(n680 ,n137 ,n667);
    nor g136(n679 ,n202 ,n667);
    nor g137(n678 ,n197 ,n667);
    nor g138(n677 ,n200 ,n667);
    nor g139(n676 ,n228 ,n668);
    nor g140(n675 ,n232 ,n668);
    nor g141(n674 ,n257 ,n668);
    nor g142(n673 ,n245 ,n668);
    nor g143(n672 ,n260 ,n668);
    nor g144(n671 ,n233 ,n668);
    nor g145(n670 ,n229 ,n668);
    nor g146(n669 ,n250 ,n668);
    not g147(n667 ,n668);
    nor g148(n666 ,n698 ,n603);
    nor g149(n665 ,n698 ,n594);
    nor g150(n664 ,n171 ,n133);
    nor g151(n663 ,n158 ,n133);
    nor g152(n662 ,n173 ,n133);
    nor g153(n661 ,n698 ,n595);
    or g154(n660 ,n533 ,n610);
    nor g155(n659 ,n282 ,n606);
    nor g156(n658 ,n698 ,n597);
    nor g157(n657 ,n698 ,n596);
    nor g158(n656 ,n698 ,n602);
    nor g159(n655 ,n698 ,n600);
    nor g160(n654 ,n698 ,n599);
    nor g161(n653 ,n698 ,n601);
    nor g162(n652 ,n698 ,n598);
    nor g163(n668 ,n267 ,n605);
    or g164(n651 ,n535 ,n609);
    nor g165(n650 ,n698 ,n592);
    nor g166(n649 ,n698 ,n591);
    nor g167(n648 ,n698 ,n590);
    or g168(n647 ,n611 ,n568);
    or g169(n646 ,n632 ,n631);
    or g170(n645 ,n630 ,n629);
    or g171(n644 ,n628 ,n627);
    or g172(n643 ,n536 ,n608);
    nor g173(n642 ,n698 ,n593);
    or g174(n641 ,n618 ,n626);
    or g175(n640 ,n617 ,n625);
    or g176(n639 ,n616 ,n624);
    or g177(n638 ,n615 ,n623);
    or g178(n637 ,n614 ,n622);
    or g179(n636 ,n613 ,n621);
    or g180(n635 ,n612 ,n620);
    or g181(n634 ,n633 ,n619);
    nor g182(n633 ,n227 ,n563);
    nor g183(n632 ,n207 ,n565);
    nor g184(n631 ,n174 ,n566);
    nor g185(n630 ,n203 ,n565);
    nor g186(n629 ,n151 ,n566);
    nor g187(n628 ,n199 ,n565);
    nor g188(n627 ,n169 ,n566);
    nor g189(n626 ,n201 ,n562);
    nor g190(n625 ,n198 ,n562);
    nor g191(n624 ,n205 ,n562);
    nor g192(n623 ,n202 ,n562);
    nor g193(n622 ,n137 ,n562);
    nor g194(n621 ,n197 ,n562);
    nor g195(n620 ,n200 ,n562);
    nor g196(n619 ,n141 ,n562);
    nor g197(n618 ,n146 ,n563);
    nor g198(n617 ,n234 ,n563);
    nor g199(n616 ,n230 ,n563);
    nor g200(n615 ,n243 ,n563);
    nor g201(n614 ,n258 ,n563);
    nor g202(n613 ,n246 ,n563);
    nor g203(n612 ,n231 ,n563);
    nor g204(n611 ,n204 ,n565);
    nor g205(n610 ,n195 ,n567);
    nor g206(n609 ,n135 ,n567);
    nor g207(n608 ,n472 ,n549);
    or g208(n607 ,n547 ,n530);
    or g209(n606 ,n18[0] ,n564);
    or g210(n605 ,n24[3] ,n569);
    nor g211(n604 ,n698 ,n561);
    nor g212(n603 ,n575 ,n583);
    nor g213(n602 ,n574 ,n582);
    nor g214(n601 ,n573 ,n581);
    nor g215(n600 ,n572 ,n580);
    nor g216(n599 ,n571 ,n579);
    nor g217(n598 ,n570 ,n578);
    nor g218(n597 ,n11[1] ,n551);
    nor g219(n596 ,n560 ,n577);
    nor g220(n595 ,n550 ,n576);
    nor g221(n594 ,n559 ,n587);
    nor g222(n593 ,n558 ,n588);
    nor g223(n592 ,n557 ,n586);
    nor g224(n591 ,n556 ,n585);
    nor g225(n590 ,n555 ,n584);
    nor g226(n589 ,n219 ,n543);
    nor g227(n588 ,n177 ,n541);
    nor g228(n587 ,n162 ,n541);
    nor g229(n586 ,n185 ,n541);
    nor g230(n585 ,n165 ,n541);
    nor g231(n584 ,n154 ,n541);
    nor g232(n583 ,n147 ,n539);
    nor g233(n582 ,n201 ,n539);
    nor g234(n581 ,n198 ,n539);
    nor g235(n580 ,n205 ,n539);
    nor g236(n579 ,n202 ,n539);
    nor g237(n578 ,n137 ,n539);
    nor g238(n577 ,n197 ,n539);
    nor g239(n576 ,n200 ,n539);
    nor g240(n575 ,n201 ,n540);
    nor g241(n574 ,n198 ,n540);
    nor g242(n573 ,n205 ,n540);
    nor g243(n572 ,n202 ,n540);
    nor g244(n571 ,n137 ,n540);
    nor g245(n570 ,n197 ,n540);
    not g246(n569 ,n568);
    not g247(n562 ,n563);
    nor g248(n561 ,n11[0] ,n537);
    nor g249(n560 ,n200 ,n540);
    nor g250(n559 ,n226 ,n542);
    nor g251(n558 ,n236 ,n542);
    nor g252(n557 ,n237 ,n542);
    nor g253(n556 ,n244 ,n542);
    nor g254(n555 ,n242 ,n542);
    nor g255(n554 ,n136 ,n543);
    nor g256(n553 ,n194 ,n543);
    nor g257(n552 ,n193 ,n543);
    nor g258(n551 ,n288 ,n532);
    nor g259(n550 ,n141 ,n540);
    or g260(n549 ,n26[0] ,n546);
    or g261(n548 ,n521 ,n531);
    nor g262(n547 ,n492 ,n534);
    nor g263(n568 ,n24[0] ,n544);
    or g264(n567 ,n698 ,n545);
    or g265(n565 ,n698 ,n542);
    or g266(n564 ,n698 ,n538);
    nor g267(n563 ,n340 ,n544);
    not g268(n546 ,n545);
    not g269(n541 ,n542);
    not g270(n539 ,n540);
    nor g271(n537 ,n289 ,n525);
    nor g272(n536 ,n285 ,n529);
    nor g273(n535 ,n698 ,n522);
    or g274(n534 ,n254 ,n520);
    or g275(n533 ,n387 ,n519);
    or g276(n532 ,n26[1] ,n525);
    or g277(n531 ,n517 ,n527);
    or g278(n530 ,n527 ,n516);
    nor g279(n545 ,n528 ,n518);
    or g280(n544 ,n285 ,n524);
    or g281(n543 ,n395 ,n526);
    nor g282(n542 ,n192 ,n524);
    nor g283(n540 ,n26[0] ,n524);
    not g284(n529 ,n528);
    or g285(n523 ,n392 ,n495);
    or g286(n522 ,n290 ,n491);
    nor g287(n521 ,n196 ,n490);
    nor g288(n520 ,n372 ,n474);
    nor g289(n519 ,n384 ,n479);
    nor g290(n518 ,n371 ,n473);
    nor g291(n517 ,n14 ,n491);
    nor g292(n516 ,n476 ,n493);
    nor g293(n528 ,n363 ,n478);
    or g294(n527 ,n395 ,n475);
    nor g295(n526 ,n284 ,n477);
    or g296(n525 ,n147 ,n481);
    or g297(n524 ,n279 ,n494);
    or g298(n515 ,n407 ,n496);
    or g299(n514 ,n404 ,n498);
    or g300(n513 ,n403 ,n499);
    or g301(n512 ,n402 ,n500);
    or g302(n511 ,n401 ,n501);
    or g303(n510 ,n400 ,n488);
    or g304(n509 ,n399 ,n489);
    or g305(n508 ,n398 ,n487);
    or g306(n507 ,n426 ,n486);
    or g307(n506 ,n393 ,n485);
    or g308(n505 ,n391 ,n484);
    or g309(n504 ,n390 ,n483);
    or g310(n503 ,n406 ,n482);
    or g311(n502 ,n408 ,n497);
    nor g312(n501 ,n181 ,n461);
    nor g313(n500 ,n152 ,n461);
    nor g314(n499 ,n190 ,n461);
    nor g315(n498 ,n155 ,n461);
    nor g316(n497 ,n183 ,n461);
    nor g317(n496 ,n166 ,n461);
    nor g318(n495 ,n150 ,n461);
    or g319(n494 ,n140 ,n462);
    not g320(n493 ,n492);
    not g321(n491 ,n490);
    nor g322(n489 ,n186 ,n461);
    nor g323(n488 ,n164 ,n461);
    nor g324(n487 ,n167 ,n461);
    nor g325(n486 ,n184 ,n461);
    nor g326(n485 ,n179 ,n461);
    nor g327(n484 ,n157 ,n461);
    nor g328(n483 ,n182 ,n461);
    nor g329(n482 ,n172 ,n461);
    or g330(n481 ,n192 ,n471);
    or g331(n480 ,n405 ,n456);
    or g332(n479 ,n285 ,n462);
    or g333(n478 ,n192 ,n463);
    or g334(n477 ,n26[0] ,n471);
    nor g335(n476 ,n467 ,n453);
    nor g336(n475 ,n26[0] ,n466);
    or g337(n474 ,n319 ,n462);
    nor g338(n473 ,n380 ,n454);
    or g339(n472 ,n698 ,n465);
    nor g340(n492 ,n343 ,n471);
    nor g341(n490 ,n282 ,n464);
    or g342(n470 ,n420 ,n432);
    or g343(n469 ,n422 ,n433);
    or g344(n468 ,n424 ,n435);
    nor g345(n467 ,n136 ,n436);
    or g346(n471 ,n196 ,n450);
    not g347(n466 ,n465);
    not g348(n464 ,n463);
    or g349(n460 ,n414 ,n442);
    or g350(n459 ,n410 ,n429);
    or g351(n458 ,n412 ,n428);
    or g352(n457 ,n418 ,n431);
    nor g353(n456 ,n19[0] ,n451);
    or g354(n455 ,n416 ,n430);
    or g355(n454 ,n282 ,n450);
    nor g356(n453 ,n18[1] ,n434);
    or g357(n452 ,n356 ,n443);
    nor g358(n465 ,n283 ,n450);
    nor g359(n463 ,n284 ,n450);
    or g360(n462 ,n26[1] ,n450);
    or g361(n461 ,n451 ,n449);
    not g362(n450 ,n449);
    nor g363(n448 ,n698 ,n373);
    nor g364(n447 ,n698 ,n383);
    nor g365(n446 ,n698 ,n381);
    nor g366(n445 ,n698 ,n425);
    nor g367(n444 ,n698 ,n397);
    nor g368(n443 ,n159 ,n394);
    or g369(n451 ,n341 ,n395);
    nor g370(n449 ,n389 ,n388);
    or g371(n442 ,n350 ,n409);
    nor g372(n441 ,n698 ,n382);
    nor g373(n440 ,n698 ,n370);
    nor g374(n439 ,n698 ,n368);
    nor g375(n438 ,n698 ,n369);
    nor g376(n437 ,n698 ,n367);
    or g377(n436 ,n275 ,n386);
    or g378(n435 ,n355 ,n423);
    nor g379(n434 ,n374 ,n385);
    or g380(n433 ,n354 ,n421);
    or g381(n432 ,n349 ,n419);
    or g382(n431 ,n351 ,n417);
    or g383(n430 ,n348 ,n415);
    or g384(n429 ,n353 ,n413);
    or g385(n428 ,n352 ,n411);
    nor g386(n427 ,n698 ,n366);
    nor g387(n426 ,n220 ,n336);
    or g388(n425 ,n148 ,n342);
    nor g389(n424 ,n232 ,n337);
    nor g390(n423 ,n146 ,n365);
    nor g391(n422 ,n257 ,n337);
    nor g392(n421 ,n234 ,n365);
    nor g393(n420 ,n245 ,n337);
    nor g394(n419 ,n230 ,n365);
    nor g395(n418 ,n243 ,n365);
    nor g396(n417 ,n260 ,n337);
    nor g397(n416 ,n258 ,n365);
    nor g398(n415 ,n233 ,n337);
    nor g399(n414 ,n229 ,n337);
    nor g400(n413 ,n231 ,n365);
    nor g401(n412 ,n228 ,n337);
    nor g402(n411 ,n227 ,n365);
    nor g403(n410 ,n250 ,n337);
    nor g404(n409 ,n246 ,n365);
    nor g405(n408 ,n213 ,n336);
    nor g406(n407 ,n211 ,n336);
    nor g407(n406 ,n216 ,n336);
    nor g408(n405 ,n206 ,n336);
    nor g409(n404 ,n223 ,n336);
    nor g410(n403 ,n142 ,n336);
    nor g411(n402 ,n222 ,n336);
    nor g412(n401 ,n214 ,n336);
    nor g413(n400 ,n139 ,n336);
    nor g414(n399 ,n208 ,n336);
    nor g415(n398 ,n210 ,n336);
    or g416(n397 ,n145 ,n345);
    nor g417(n393 ,n218 ,n336);
    nor g418(n392 ,n221 ,n336);
    nor g419(n391 ,n215 ,n336);
    nor g420(n390 ,n209 ,n336);
    or g421(n389 ,n329 ,n330);
    or g422(n388 ,n325 ,n323);
    nor g423(n387 ,n698 ,n343);
    nor g424(n386 ,n308 ,n317);
    nor g425(n385 ,n273 ,n331);
    nor g426(n384 ,n3 ,n335);
    or g427(n383 ,n27[4] ,n342);
    nor g428(n382 ,n334 ,n360);
    or g429(n381 ,n22[4] ,n345);
    nor g430(n380 ,n284 ,n338);
    nor g431(n379 ,n698 ,n320);
    nor g432(n378 ,n698 ,n324);
    nor g433(n377 ,n698 ,n326);
    nor g434(n376 ,n698 ,n327);
    nor g435(n375 ,n698 ,n328);
    nor g436(n374 ,n18[0] ,n318);
    nor g437(n373 ,n11[2] ,n341);
    or g438(n372 ,n270 ,n332);
    or g439(n371 ,n26[0] ,n362);
    nor g440(n370 ,n346 ,n359);
    nor g441(n369 ,n333 ,n357);
    nor g442(n368 ,n364 ,n358);
    nor g443(n367 ,n322 ,n321);
    nor g444(n366 ,n347 ,n361);
    or g445(n396 ,n282 ,n338);
    or g446(n395 ,n698 ,n344);
    nor g447(n364 ,n240 ,n316);
    nor g448(n363 ,n144 ,n283);
    nor g449(n362 ,n144 ,n281);
    nor g450(n361 ,n160 ,n315);
    nor g451(n360 ,n191 ,n315);
    nor g452(n359 ,n187 ,n315);
    nor g453(n358 ,n189 ,n315);
    nor g454(n357 ,n176 ,n315);
    nor g455(n356 ,n138 ,n280);
    nor g456(n355 ,n225 ,n280);
    nor g457(n354 ,n253 ,n280);
    nor g458(n353 ,n248 ,n280);
    nor g459(n352 ,n241 ,n280);
    nor g460(n351 ,n143 ,n280);
    nor g461(n350 ,n235 ,n280);
    nor g462(n349 ,n249 ,n280);
    nor g463(n348 ,n239 ,n280);
    nor g464(n347 ,n259 ,n316);
    nor g465(n346 ,n149 ,n316);
    or g466(n365 ,n138 ,n286);
    not g467(n340 ,n339);
    or g468(n335 ,n135 ,n271);
    nor g469(n334 ,n255 ,n316);
    nor g470(n332 ,n192 ,n288);
    or g471(n331 ,n194 ,n265);
    or g472(n330 ,n312 ,n274);
    or g473(n329 ,n313 ,n297);
    nor g474(n328 ,n304 ,n296);
    nor g475(n327 ,n306 ,n293);
    nor g476(n326 ,n307 ,n298);
    or g477(n325 ,n261 ,n268);
    nor g478(n324 ,n305 ,n292);
    or g479(n323 ,n266 ,n262);
    nor g480(n322 ,n224 ,n282);
    nor g481(n321 ,n192 ,n281);
    nor g482(n320 ,n314 ,n294);
    nor g483(n319 ,n26[0] ,n287);
    nor g484(n318 ,n309 ,n295);
    or g485(n317 ,n18[0] ,n299);
    or g486(n345 ,n276 ,n278);
    nor g487(n344 ,n26[1] ,n291);
    or g488(n343 ,n26[0] ,n289);
    or g489(n342 ,n264 ,n263);
    nor g490(n341 ,n192 ,n283);
    nor g491(n339 ,n311 ,n310);
    nor g492(n338 ,n303 ,n272);
    or g493(n337 ,n23[3] ,n286);
    or g494(n336 ,n283 ,n285);
    not g495(n315 ,n316);
    nor g496(n314 ,n134 ,n163);
    or g497(n313 ,n142 ,n222);
    or g498(n312 ,n214 ,n139);
    or g499(n311 ,n204 ,n207);
    or g500(n310 ,n203 ,n199);
    nor g501(n309 ,n193 ,n175);
    nor g502(n308 ,n193 ,n188);
    nor g503(n307 ,n134 ,n178);
    nor g504(n306 ,n134 ,n180);
    nor g505(n305 ,n134 ,n153);
    nor g506(n304 ,n134 ,n161);
    or g507(n303 ,n194 ,n136);
    nor g508(n302 ,n224 ,n698);
    nor g509(n301 ,n212 ,n698);
    nor g510(n300 ,n217 ,n698);
    nor g511(n299 ,n170 ,n18[2]);
    nor g512(n298 ,n238 ,n733);
    or g513(n297 ,n206 ,n19[1]);
    nor g514(n296 ,n256 ,n733);
    nor g515(n295 ,n156 ,n18[2]);
    nor g516(n294 ,n251 ,n733);
    nor g517(n293 ,n247 ,n733);
    nor g518(n292 ,n252 ,n733);
    nor g519(n316 ,n697 ,n168);
    not g520(n291 ,n290);
    not g521(n288 ,n287);
    not g522(n283 ,n284);
    not g523(n281 ,n282);
    or g524(n279 ,n196 ,n135);
    or g525(n278 ,n22[3] ,n22[2]);
    nor g526(n277 ,n195 ,n698);
    or g527(n276 ,n22[1] ,n22[0]);
    nor g528(n275 ,n194 ,n7[3]);
    or g529(n274 ,n19[6] ,n19[7]);
    nor g530(n273 ,n193 ,n7[1]);
    or g531(n272 ,n193 ,n18[3]);
    nor g532(n271 ,n4 ,n722);
    nor g533(n270 ,n135 ,n14);
    nor g534(n269 ,n192 ,n698);
    or g535(n268 ,n19[10] ,n19[11]);
    or g536(n267 ,n24[1] ,n24[2]);
    or g537(n266 ,n19[12] ,n19[13]);
    nor g538(n265 ,n18[2] ,n7[5]);
    or g539(n264 ,n27[1] ,n27[0]);
    or g540(n263 ,n27[3] ,n27[2]);
    or g541(n262 ,n19[14] ,n19[15]);
    or g542(n261 ,n19[8] ,n19[9]);
    nor g543(n290 ,n26[0] ,n26[2]);
    or g544(n289 ,n195 ,n26[2]);
    nor g545(n287 ,n135 ,n4);
    or g546(n286 ,n698 ,n134);
    or g547(n285 ,n192 ,n698);
    nor g548(n284 ,n195 ,n135);
    nor g549(n282 ,n26[1] ,n26[2]);
    or g550(n280 ,n698 ,n733);
    not g551(n260 ,n20[3]);
    not g552(n259 ,n27[0]);
    not g553(n258 ,n21[4]);
    not g554(n257 ,n20[1]);
    not g555(n256 ,n22[4]);
    not g556(n255 ,n27[1]);
    not g557(n254 ,n15);
    not g558(n253 ,n9[1]);
    not g559(n252 ,n22[1]);
    not g560(n251 ,n22[0]);
    not g561(n250 ,n20[6]);
    not g562(n249 ,n9[2]);
    not g563(n248 ,n9[6]);
    not g564(n247 ,n22[3]);
    not g565(n246 ,n21[5]);
    not g566(n245 ,n20[2]);
    not g567(n244 ,n22[3]);
    not g568(n243 ,n21[3]);
    not g569(n242 ,n22[4]);
    not g570(n241 ,n9[7]);
    not g571(n240 ,n27[3]);
    not g572(n239 ,n9[4]);
    not g573(n238 ,n22[2]);
    not g574(n237 ,n22[2]);
    not g575(n236 ,n22[1]);
    not g576(n235 ,n9[5]);
    not g577(n234 ,n21[1]);
    not g578(n233 ,n20[4]);
    not g579(n232 ,n20[0]);
    not g580(n231 ,n21[6]);
    not g581(n230 ,n21[2]);
    not g582(n229 ,n20[5]);
    not g583(n228 ,n20[7]);
    not g584(n227 ,n21[7]);
    not g585(n226 ,n22[0]);
    not g586(n225 ,n9[0]);
    not g587(n224 ,n16);
    not g588(n223 ,n19[1]);
    not g589(n222 ,n19[3]);
    not g590(n221 ,n19[14]);
    not g591(n220 ,n19[8]);
    not g592(n219 ,n18[3]);
    not g593(n218 ,n19[9]);
    not g594(n217 ,n11[0]);
    not g595(n216 ,n19[12]);
    not g596(n215 ,n19[10]);
    not g597(n214 ,n19[4]);
    not g598(n213 ,n19[15]);
    not g599(n212 ,n11[1]);
    not g600(n211 ,n19[13]);
    not g601(n210 ,n19[7]);
    not g602(n209 ,n19[11]);
    not g603(n208 ,n19[6]);
    not g604(n207 ,n24[1]);
    not g605(n206 ,n19[0]);
    not g606(n205 ,n25[2]);
    not g607(n204 ,n24[0]);
    not g608(n203 ,n24[2]);
    not g609(n202 ,n25[3]);
    not g610(n201 ,n25[0]);
    not g611(n200 ,n25[6]);
    not g612(n199 ,n24[3]);
    not g613(n198 ,n25[1]);
    not g614(n197 ,n25[5]);
    not g615(n196 ,n14);
    not g616(n195 ,n26[1]);
    not g617(n194 ,n18[0]);
    not g618(n193 ,n18[2]);
    not g619(n192 ,n26[0]);
    not g620(n191 ,n737);
    not g621(n190 ,n704);
    not g622(n189 ,n735);
    not g623(n188 ,n7[0]);
    not g624(n187 ,n736);
    not g625(n186 ,n708);
    not g626(n185 ,n730);
    not g627(n184 ,n710);
    not g628(n183 ,n717);
    not g629(n182 ,n713);
    not g630(n181 ,n706);
    not g631(n180 ,n724);
    not g632(n179 ,n711);
    not g633(n178 ,n725);
    not g634(n177 ,n731);
    not g635(n176 ,n734);
    not g636(n175 ,n7[2]);
    not g637(n174 ,n699);
    not g638(n173 ,n702);
    not g639(n172 ,n714);
    not g640(n171 ,n718);
    not g641(n170 ,n7[4]);
    not g642(n169 ,n701);
    not g643(n168 ,n721);
    not g644(n167 ,n709);
    not g645(n166 ,n715);
    not g646(n165 ,n729);
    not g647(n164 ,n707);
    not g648(n163 ,n727);
    not g649(n162 ,n732);
    not g650(n161 ,n723);
    not g651(n160 ,n738);
    not g652(n159 ,n720);
    not g653(n158 ,n719);
    not g654(n157 ,n712);
    not g655(n156 ,n7[6]);
    not g656(n155 ,n703);
    not g657(n154 ,n728);
    not g658(n153 ,n726);
    not g659(n152 ,n705);
    not g660(n151 ,n700);
    not g661(n150 ,n716);
    not g662(n149 ,n27[2]);
    not g663(n148 ,n27[4]);
    not g664(n147 ,n6);
    not g665(n146 ,n21[0]);
    not g666(n145 ,n22[4]);
    not g667(n144 ,n2);
    not g668(n143 ,n9[3]);
    not g669(n142 ,n19[2]);
    not g670(n141 ,n25[7]);
    not g671(n140 ,n4);
    not g672(n139 ,n19[5]);
    not g673(n138 ,n23[3]);
    not g674(n137 ,n25[4]);
    not g675(n136 ,n18[1]);
    not g676(n135 ,n26[2]);
    not g677(n134 ,n733);
    or g678(n133 ,n396 ,n564);
    xor g679(n723 ,n22[4] ,n32);
    xor g680(n724 ,n22[3] ,n30);
    nor g681(n32 ,n22[3] ,n31);
    xor g682(n725 ,n22[2] ,n28);
    not g683(n31 ,n30);
    nor g684(n30 ,n22[2] ,n29);
    xnor g685(n726 ,n22[1] ,n22[0]);
    not g686(n29 ,n28);
    nor g687(n28 ,n22[1] ,n22[0]);
    not g688(n727 ,n22[0]);
    or g689(n722 ,n34 ,n35);
    or g690(n35 ,n27[3] ,n33);
    or g691(n34 ,n27[2] ,n27[0]);
    or g692(n33 ,n27[4] ,n27[1]);
    or g693(n733 ,n37 ,n38);
    or g694(n38 ,n22[3] ,n36);
    or g695(n37 ,n22[2] ,n22[0]);
    or g696(n36 ,n22[4] ,n22[1]);
    xor g697(n717 ,n19[15] ,n94);
    nor g698(n716 ,n93 ,n94);
    nor g699(n94 ,n50 ,n92);
    nor g700(n93 ,n19[14] ,n91);
    nor g701(n715 ,n90 ,n91);
    not g702(n92 ,n91);
    nor g703(n91 ,n40 ,n89);
    nor g704(n90 ,n19[13] ,n88);
    nor g705(n714 ,n87 ,n88);
    not g706(n89 ,n88);
    nor g707(n88 ,n53 ,n86);
    nor g708(n87 ,n19[12] ,n85);
    nor g709(n713 ,n84 ,n85);
    not g710(n86 ,n85);
    nor g711(n85 ,n49 ,n83);
    nor g712(n84 ,n19[11] ,n82);
    nor g713(n712 ,n81 ,n82);
    not g714(n83 ,n82);
    nor g715(n82 ,n51 ,n80);
    nor g716(n81 ,n19[10] ,n79);
    nor g717(n711 ,n78 ,n79);
    not g718(n80 ,n79);
    nor g719(n79 ,n48 ,n77);
    nor g720(n78 ,n19[9] ,n76);
    nor g721(n710 ,n75 ,n76);
    not g722(n77 ,n76);
    nor g723(n76 ,n45 ,n74);
    nor g724(n75 ,n19[8] ,n73);
    nor g725(n709 ,n72 ,n73);
    not g726(n74 ,n73);
    nor g727(n73 ,n46 ,n71);
    nor g728(n72 ,n19[7] ,n70);
    nor g729(n708 ,n69 ,n70);
    not g730(n71 ,n70);
    nor g731(n70 ,n39 ,n68);
    nor g732(n69 ,n19[6] ,n67);
    nor g733(n707 ,n66 ,n67);
    not g734(n68 ,n67);
    nor g735(n67 ,n44 ,n65);
    nor g736(n66 ,n19[5] ,n64);
    nor g737(n706 ,n63 ,n64);
    not g738(n65 ,n64);
    nor g739(n64 ,n42 ,n62);
    nor g740(n63 ,n19[4] ,n61);
    nor g741(n705 ,n60 ,n61);
    not g742(n62 ,n61);
    nor g743(n61 ,n41 ,n59);
    nor g744(n60 ,n19[3] ,n58);
    nor g745(n704 ,n57 ,n58);
    not g746(n59 ,n58);
    nor g747(n58 ,n43 ,n56);
    nor g748(n57 ,n19[2] ,n55);
    nor g749(n703 ,n55 ,n54);
    not g750(n56 ,n55);
    nor g751(n55 ,n47 ,n52);
    nor g752(n54 ,n19[1] ,n19[0]);
    not g753(n53 ,n19[12]);
    not g754(n52 ,n19[0]);
    not g755(n51 ,n19[10]);
    not g756(n50 ,n19[14]);
    not g757(n49 ,n19[11]);
    not g758(n48 ,n19[9]);
    not g759(n47 ,n19[1]);
    not g760(n46 ,n19[7]);
    not g761(n45 ,n19[8]);
    not g762(n44 ,n19[5]);
    not g763(n43 ,n19[2]);
    not g764(n42 ,n19[4]);
    not g765(n41 ,n19[3]);
    not g766(n40 ,n19[13]);
    not g767(n39 ,n19[6]);
    xor g768(n702 ,n18[3] ,n102);
    nor g769(n719 ,n101 ,n102);
    nor g770(n102 ,n97 ,n100);
    nor g771(n101 ,n18[2] ,n99);
    nor g772(n718 ,n99 ,n98);
    not g773(n100 ,n99);
    nor g774(n99 ,n95 ,n96);
    nor g775(n98 ,n18[1] ,n18[0]);
    not g776(n97 ,n18[2]);
    not g777(n96 ,n18[0]);
    not g778(n95 ,n18[1]);
    xor g779(n701 ,n24[3] ,n110);
    nor g780(n700 ,n109 ,n110);
    nor g781(n110 ,n105 ,n108);
    nor g782(n109 ,n24[2] ,n107);
    nor g783(n699 ,n107 ,n106);
    not g784(n108 ,n107);
    nor g785(n107 ,n103 ,n104);
    nor g786(n106 ,n24[1] ,n24[0]);
    not g787(n105 ,n24[2]);
    not g788(n104 ,n24[0]);
    not g789(n103 ,n24[1]);
    xor g790(n728 ,n22[4] ,n121);
    nor g791(n729 ,n120 ,n121);
    nor g792(n121 ,n112 ,n119);
    nor g793(n120 ,n22[3] ,n118);
    nor g794(n730 ,n117 ,n118);
    not g795(n119 ,n118);
    nor g796(n118 ,n113 ,n116);
    nor g797(n117 ,n22[2] ,n115);
    nor g798(n731 ,n115 ,n114);
    not g799(n116 ,n115);
    nor g800(n115 ,n111 ,n732);
    nor g801(n114 ,n22[1] ,n22[0]);
    not g802(n113 ,n22[2]);
    not g803(n732 ,n22[0]);
    not g804(n112 ,n22[3]);
    not g805(n111 ,n22[1]);
    nor g806(n735 ,n131 ,n132);
    nor g807(n132 ,n123 ,n130);
    nor g808(n131 ,n27[3] ,n129);
    nor g809(n736 ,n128 ,n129);
    not g810(n130 ,n129);
    nor g811(n129 ,n124 ,n127);
    nor g812(n128 ,n27[2] ,n126);
    nor g813(n737 ,n126 ,n125);
    not g814(n127 ,n126);
    nor g815(n126 ,n122 ,n738);
    nor g816(n125 ,n27[1] ,n27[0]);
    not g817(n124 ,n27[2]);
    not g818(n738 ,n27[0]);
    not g819(n123 ,n27[3]);
    not g820(n122 ,n27[1]);
    not g821(n721 ,n27[4]);
    buf g822(n720 ,n23[3]);
    buf g823(n333 ,n27[4]);
    buf g824(n394 ,n286);
    buf g825(n734 ,n132);
    not g826(n538 ,n526);
    buf g827(n566 ,n544);
endmodule
