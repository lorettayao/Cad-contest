module top(n0, n1, n2, n6, n3, n7, n5, n12, n4, n8, n9, n10, n11, n13, n14, n15, n16);
    input n0, n1, n2, n3, n4;
    input [7:0] n5;
    output n6, n7, n8, n9, n10, n11;
    output [7:0] n12, n13, n14, n15;
    output [15:0] n16;
    wire n0, n1, n2, n3, n4;
    wire [7:0] n5;
    wire n6, n7, n8, n9, n10, n11;
    wire [7:0] n12, n13, n14, n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [2:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [4:0] n21;
    wire [3:0] n22;
    wire [3:0] n23;
    wire [7:0] n24;
    wire [2:0] n25;
    wire [15:0] n26;
    wire [2:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [7:0] n37;
    wire [7:0] n38;
    wire [7:0] n39;
    wire [7:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [4:0] n44;
    wire [3:0] n45;
    wire [3:0] n46;
    wire [7:0] n47;
    wire [2:0] n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526, n527, n528;
    wire n529, n530, n531, n532, n533, n534, n535, n536;
    wire n537, n538, n539, n540, n541, n542, n543, n544;
    wire n545, n546, n547, n548, n549, n550, n551, n552;
    wire n553, n554, n555, n556, n557, n558, n559, n560;
    wire n561, n562, n563, n564, n565, n566, n567, n568;
    wire n569, n570, n571, n572, n573, n574, n575, n576;
    wire n577, n578, n579, n580, n581, n582, n583, n584;
    wire n585, n586, n587, n588, n589, n590, n591, n592;
    wire n593, n594, n595, n596, n597, n598, n599, n600;
    wire n601, n602, n603, n604, n605, n606, n607, n608;
    wire n609, n610, n611, n612, n613, n614, n615, n616;
    wire n617, n618, n619, n620, n621, n622, n623, n624;
    wire n625, n626, n627, n628, n629, n630, n631, n632;
    wire n633, n634, n635, n636, n637, n638, n639, n640;
    wire n641, n642, n643, n644, n645, n646, n647, n648;
    wire n649, n650, n651, n652, n653, n654, n655, n656;
    wire n657, n658, n659, n660, n661, n662, n663, n664;
    wire n665, n666, n667, n668, n669, n670, n671, n672;
    wire n673, n674, n675, n676, n677, n678, n679, n680;
    wire n681, n682, n683, n684, n685, n686, n687, n688;
    wire n689, n690, n691, n692, n693, n694, n695, n696;
    wire n697, n698, n699, n700, n701, n702, n703, n704;
    wire n705, n706, n707, n708, n709, n710, n711, n712;
    wire n713, n714, n715, n716, n717, n718, n719, n720;
    wire n721, n722, n723, n724, n725, n726, n727, n728;
    wire n729, n730, n731, n732, n733, n734, n735, n736;
    wire n737, n738, n739, n740, n741, n742, n743, n744;
    wire n745, n746, n747, n748, n749, n750, n751, n752;
    wire n753, n754, n755, n756, n757, n758, n759, n760;
    wire n761, n762, n763, n764, n765, n766, n767, n768;
    wire n769, n770, n771, n772, n773, n774, n775, n776;
    wire n777, n778, n779, n780, n781, n782, n783, n784;
    wire n785, n786, n787, n788, n789, n790, n791, n792;
    wire n793, n794, n795, n796, n797, n798, n799, n800;
    wire n801, n802, n803, n804, n805, n806, n807, n808;
    wire n809, n810, n811, n812, n813, n814, n815, n816;
    wire n817, n818, n819, n820, n821, n822, n823, n824;
    wire n825, n826, n827, n828, n829, n830, n831, n832;
    wire n833, n834, n835, n836, n837, n838, n839, n840;
    wire n841, n842, n843, n844, n845, n846, n847, n848;
    wire n849, n850, n851, n852, n853, n854, n855, n856;
    wire n857, n858, n859, n860, n861, n862, n863, n864;
    wire n865, n866, n867, n868, n869, n870, n871, n872;
    wire n873, n874, n875, n876, n877, n878, n879, n880;
    wire n881, n882, n883, n884, n885, n886, n887, n888;
    wire n889, n890, n891, n892, n893, n894, n895, n896;
    wire n897, n898, n899, n900, n901, n902, n903, n904;
    wire n905, n906, n907, n908, n909, n910, n911, n912;
    wire n913, n914, n915, n916, n917, n918, n919, n920;
    wire n921, n922, n923, n924, n925, n926, n927, n928;
    wire n929, n930, n931, n932, n933, n934, n935, n936;
    wire n937, n938, n939, n940, n941, n942, n943, n944;
    wire n945, n946, n947, n948, n949, n950, n951, n952;
    wire n953, n954, n955, n956, n957, n958, n959, n960;
    wire n961, n962, n963, n964, n965, n966, n967, n968;
    wire n969, n970, n971, n972, n973, n974, n975, n976;
    wire n977, n978, n979, n980, n981, n982, n983, n984;
    wire n985, n986, n987, n988, n989, n990, n991, n992;
    wire n993, n994, n995, n996, n997, n998, n999, n1000;
    wire n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
    wire n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
    wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
    wire n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
    wire n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
    wire n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
    wire n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
    wire n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064;
    wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
    wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
    wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
    wire n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096;
    wire n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
    wire n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;
    wire n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120;
    wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
    wire n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136;
    wire n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
    wire n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152;
    wire n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
    wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168;
    wire n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176;
    wire n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184;
    wire n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192;
    wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
    wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
    wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
    wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
    wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
    wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
    wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
    wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
    wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
    wire n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
    wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
    wire n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288;
    wire n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;
    wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;
    wire n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;
    wire n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;
    wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
    wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
    wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;
    wire n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;
    wire n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;
    wire n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368;
    wire n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;
    wire n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384;
    wire n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392;
    wire n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400;
    wire n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408;
    wire n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416;
    wire n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424;
    wire n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432;
    wire n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440;
    wire n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448;
    wire n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456;
    wire n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464;
    wire n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472;
    wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480;
    wire n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488;
    wire n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496;
    wire n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504;
    wire n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512;
    wire n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520;
    wire n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528;
    wire n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536;
    wire n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544;
    wire n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552;
    wire n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560;
    wire n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568;
    wire n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576;
    wire n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584;
    wire n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592;
    wire n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600;
    wire n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608;
    wire n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616;
    wire n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624;
    wire n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632;
    wire n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640;
    wire n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648;
    wire n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656;
    wire n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664;
    wire n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672;
    wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
    wire n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688;
    wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
    wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
    wire n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712;
    wire n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720;
    wire n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728;
    wire n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736;
    wire n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744;
    wire n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752;
    wire n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760;
    wire n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768;
    wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
    wire n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;
    wire n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792;
    wire n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800;
    wire n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808;
    wire n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816;
    wire n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824;
    wire n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832;
    wire n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840;
    wire n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848;
    wire n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856;
    wire n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864;
    wire n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872;
    wire n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880;
    wire n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888;
    wire n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896;
    wire n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904;
    wire n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912;
    wire n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920;
    wire n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928;
    wire n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936;
    wire n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944;
    buf g0(n46[3], 1'b0);
    buf g1(n46[2], 1'b0);
    buf g2(n46[1], 1'b0);
    buf g3(n46[0], 1'b0);
    buf g4(n22[3], 1'b0);
    buf g5(n22[2], 1'b0);
    buf g6(n22[1], 1'b0);
    buf g7(n22[0], 1'b0);
    buf g8(n16[0], 1'b0);
    buf g9(n16[1], 1'b0);
    buf g10(n16[2], 1'b0);
    buf g11(n16[3], 1'b0);
    buf g12(n16[4], 1'b0);
    buf g13(n16[5], 1'b0);
    buf g14(n16[6], 1'b0);
    buf g15(n16[7], 1'b0);
    buf g16(n16[8], 1'b0);
    buf g17(n16[9], 1'b0);
    buf g18(n16[10], 1'b0);
    buf g19(n16[11], 1'b0);
    buf g20(n16[12], 1'b0);
    buf g21(n16[13], 1'b0);
    buf g22(n16[14], 1'b0);
    buf g23(n16[15], 1'b0);
    buf g24(n15[0], 1'b0);
    buf g25(n15[1], 1'b0);
    buf g26(n15[2], 1'b0);
    buf g27(n15[3], n13[1]);
    buf g28(n15[4], n13[2]);
    buf g29(n15[5], n13[5]);
    buf g30(n14[0], 1'b0);
    buf g31(n14[2], 1'b0);
    buf g32(n14[3], 1'b0);
    buf g33(n14[4], 1'b0);
    buf g34(n14[5], 1'b0);
    buf g35(n14[6], 1'b0);
    buf g36(n14[7], 1'b0);
    buf g37(n13[0], 1'b0);
    not g38(n1879 ,n1937);
    not g39(n1878 ,n1919);
    not g40(n1877 ,n4);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n575), .Q(n7));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n14[1]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n618), .Q(n13[1]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n794), .Q(n13[2]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n797), .Q(n13[5]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n619), .Q(n15[6]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n621), .Q(n15[7]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1485), .Q(n17[0]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1487), .Q(n17[1]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1496), .Q(n17[2]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1512), .Q(n17[3]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1517), .Q(n17[4]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1520), .Q(n17[5]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1504), .Q(n17[6]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1503), .Q(n17[7]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1505), .Q(n17[8]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1502), .Q(n17[9]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1499), .Q(n17[10]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n18[0]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n18[1]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n18[2]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n11));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n896), .Q(n12[0]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n888), .Q(n12[1]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n889), .Q(n12[2]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n890), .Q(n12[3]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n895), .Q(n12[4]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n893), .Q(n12[5]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n898), .Q(n12[6]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n891), .Q(n12[7]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n9));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n19[0]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n19[1]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n19[2]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n19[3]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n19[4]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n19[5]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n19[6]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n19[7]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n20[0]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1693), .Q(n20[1]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1688), .Q(n20[2]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1684), .Q(n20[3]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1678), .Q(n20[4]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n20[5]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n20[6]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1673), .Q(n20[7]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1509), .Q(n21[0]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n708), .Q(n21[0]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1508), .Q(n21[1]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n707), .Q(n21[1]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1507), .Q(n21[2]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n724), .Q(n21[2]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1506), .Q(n21[3]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n706), .Q(n21[3]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1513), .Q(n21[4]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n711), .Q(n21[4]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n874), .Q(n22[0]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n894), .Q(n22[1]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n884), .Q(n22[2]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n900), .Q(n22[3]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1501), .Q(n23[0]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1500), .Q(n23[1]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1498), .Q(n23[2]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1497), .Q(n23[3]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n989), .Q(n24[0]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n988), .Q(n24[1]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n987), .Q(n24[2]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n986), .Q(n24[3]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n985), .Q(n24[4]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n990), .Q(n24[5]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n984), .Q(n24[6]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n991), .Q(n24[7]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n25[0]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n25[1]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n25[2]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n796), .Q(n13[3]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n795), .Q(n13[4]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n634), .Q(n13[6]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n620), .Q(n13[7]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n983), .Q(n26[0]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n982), .Q(n26[1]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n981), .Q(n26[2]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n980), .Q(n26[3]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n979), .Q(n26[4]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n978), .Q(n26[5]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n977), .Q(n26[6]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n976), .Q(n26[7]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n975), .Q(n26[8]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n974), .Q(n26[9]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n973), .Q(n26[10]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1493), .Q(n27[0]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1494), .Q(n27[1]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1492), .Q(n27[2]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n10));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1510), .Q(n8));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1339), .Q(n28[0]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1338), .Q(n28[1]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1336), .Q(n28[2]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1389), .Q(n28[3]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1396), .Q(n28[4]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1455), .Q(n28[5]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1448), .Q(n28[6]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n28[7]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n29[0]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1331), .Q(n29[1]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n29[2]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n29[3]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1337), .Q(n29[4]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n29[5]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1325), .Q(n29[6]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n29[7]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n30[0]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1340), .Q(n30[1]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n30[2]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n30[3]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n30[4]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n30[5]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n30[6]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1445), .Q(n30[7]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1386), .Q(n31[0]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n31[1]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1378), .Q(n31[2]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1335), .Q(n31[3]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n31[4]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n31[5]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n31[6]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n31[7]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n32[0]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n32[1]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n32[2]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n32[3]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n32[4]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n32[5]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1308), .Q(n32[6]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n32[7]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n33[0]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n33[1]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1303), .Q(n33[2]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n33[3]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n33[4]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1299), .Q(n33[5]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n33[6]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n33[7]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n34[0]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1294), .Q(n34[1]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n34[2]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n34[3]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n34[4]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1438), .Q(n34[5]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1439), .Q(n34[6]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1440), .Q(n34[7]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1441), .Q(n35[0]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1442), .Q(n35[1]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1443), .Q(n35[2]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1444), .Q(n35[3]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1446), .Q(n35[4]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1447), .Q(n35[5]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1449), .Q(n35[6]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1450), .Q(n35[7]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n36[0]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n36[1]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n36[2]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1454), .Q(n36[3]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1456), .Q(n36[4]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1457), .Q(n36[5]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1458), .Q(n36[6]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1459), .Q(n36[7]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1460), .Q(n37[0]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n37[1]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n37[2]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n37[3]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1398), .Q(n37[4]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n37[5]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1395), .Q(n37[6]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1394), .Q(n37[7]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1393), .Q(n38[0]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1392), .Q(n38[1]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1391), .Q(n38[2]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1390), .Q(n38[3]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1388), .Q(n38[4]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1387), .Q(n38[5]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1385), .Q(n38[6]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1384), .Q(n38[7]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1383), .Q(n39[0]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1382), .Q(n39[1]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1381), .Q(n39[2]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1380), .Q(n39[3]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1379), .Q(n39[4]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1377), .Q(n39[5]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1376), .Q(n39[6]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1375), .Q(n39[7]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1374), .Q(n40[0]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1373), .Q(n40[1]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1372), .Q(n40[2]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1371), .Q(n40[3]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1369), .Q(n40[4]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1370), .Q(n40[5]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n40[6]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n40[7]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n41[0]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n41[1]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n41[2]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n41[3]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n41[4]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n41[5]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n41[6]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n41[7]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n42[0]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n42[1]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n42[2]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n42[3]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n42[4]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n42[5]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n42[6]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1351), .Q(n42[7]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n43[0]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n43[1]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n43[2]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n43[3]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n43[4]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n43[5]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1344), .Q(n43[6]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n43[7]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n972), .Q(n44[0]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n775), .Q(n44[0]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n971), .Q(n44[1]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n774), .Q(n44[1]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n970), .Q(n44[2]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n773), .Q(n44[2]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n969), .Q(n44[3]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n772), .Q(n44[3]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n968), .Q(n44[4]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n771), .Q(n44[4]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n45[0]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n45[1]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n45[2]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n45[3]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1491), .Q(n46[0]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1490), .Q(n46[1]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1489), .Q(n46[2]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1488), .Q(n46[3]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n6));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n47[0]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n47[1]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n47[2]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n47[3]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n47[4]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n47[5]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n47[6]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n47[7]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n48[0]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n48[1]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n48[2]));
    or g295(n1876 ,n1545 ,n1868);
    or g296(n1875 ,n1546 ,n1867);
    or g297(n1874 ,n1544 ,n1869);
    or g298(n1873 ,n1541 ,n1864);
    or g299(n1872 ,n1542 ,n1863);
    or g300(n1871 ,n1543 ,n1866);
    or g301(n1870 ,n1540 ,n1865);
    or g302(n1869 ,n922 ,n1861);
    or g303(n1868 ,n926 ,n1860);
    or g304(n1867 ,n925 ,n1859);
    or g305(n1866 ,n924 ,n1858);
    or g306(n1865 ,n934 ,n1857);
    or g307(n1864 ,n921 ,n1856);
    or g308(n1863 ,n923 ,n1855);
    or g309(n1862 ,n1581 ,n1854);
    or g310(n1861 ,n1627 ,n1853);
    or g311(n1860 ,n1647 ,n1852);
    or g312(n1859 ,n1665 ,n1851);
    or g313(n1858 ,n1613 ,n1850);
    or g314(n1857 ,n1571 ,n1849);
    or g315(n1856 ,n1584 ,n1848);
    or g316(n1855 ,n1599 ,n1847);
    or g317(n1854 ,n1539 ,n1846);
    or g318(n1853 ,n1805 ,n1845);
    or g319(n1852 ,n1808 ,n1844);
    or g320(n1851 ,n1811 ,n1843);
    or g321(n1850 ,n1802 ,n1842);
    or g322(n1849 ,n1795 ,n1841);
    or g323(n1848 ,n1771 ,n1840);
    or g324(n1847 ,n1799 ,n1839);
    or g325(n1846 ,n1792 ,n1838);
    or g326(n1845 ,n1723 ,n1835);
    or g327(n1844 ,n1730 ,n1830);
    or g328(n1843 ,n1769 ,n1837);
    or g329(n1842 ,n1716 ,n1834);
    or g330(n1841 ,n1694 ,n1831);
    or g331(n1840 ,n1701 ,n1832);
    or g332(n1839 ,n1709 ,n1833);
    or g333(n1838 ,n1685 ,n1836);
    or g334(n1837 ,n1658 ,n1828);
    or g335(n1836 ,n1659 ,n1821);
    or g336(n1835 ,n1621 ,n1826);
    or g337(n1834 ,n1608 ,n1825);
    or g338(n1833 ,n1671 ,n1824);
    or g339(n1832 ,n1578 ,n1823);
    or g340(n1831 ,n1565 ,n1829);
    or g341(n1830 ,n1635 ,n1827);
    or g342(n1829 ,n1794 ,n1793);
    or g343(n1828 ,n1810 ,n1809);
    or g344(n1827 ,n1807 ,n1806);
    or g345(n1826 ,n1804 ,n1803);
    or g346(n1825 ,n1801 ,n1800);
    or g347(n1824 ,n1814 ,n1815);
    or g348(n1823 ,n1797 ,n1796);
    or g349(n1822 ,n1744 ,n1813);
    or g350(n1821 ,n1791 ,n1790);
    nor g351(n1820 ,n248 ,n1785);
    nor g352(n1819 ,n251 ,n1784);
    nor g353(n1818 ,n245 ,n1783);
    or g354(n1817 ,n1758 ,n1789);
    or g355(n1816 ,n1743 ,n1812);
    or g356(n1815 ,n1706 ,n1705);
    or g357(n1814 ,n1708 ,n1707);
    nor g358(n1813 ,n386 ,n1770);
    nor g359(n1812 ,n363 ,n1770);
    or g360(n1811 ,n1767 ,n1768);
    or g361(n1810 ,n1704 ,n1735);
    or g362(n1809 ,n1734 ,n1733);
    or g363(n1808 ,n1732 ,n1731);
    or g364(n1807 ,n1729 ,n1728);
    or g365(n1806 ,n1727 ,n1726);
    or g366(n1805 ,n1725 ,n1724);
    or g367(n1804 ,n1722 ,n1721);
    or g368(n1803 ,n1720 ,n1719);
    or g369(n1802 ,n1718 ,n1717);
    or g370(n1801 ,n1715 ,n1714);
    or g371(n1800 ,n1713 ,n1712);
    or g372(n1799 ,n1711 ,n1710);
    or g373(n1798 ,n1757 ,n1749);
    or g374(n1797 ,n1700 ,n1699);
    or g375(n1796 ,n1698 ,n1697);
    or g376(n1795 ,n1696 ,n1695);
    or g377(n1794 ,n1692 ,n1691);
    or g378(n1793 ,n1690 ,n1689);
    or g379(n1792 ,n1686 ,n1687);
    or g380(n1791 ,n1683 ,n1682);
    or g381(n1790 ,n1681 ,n1680);
    nor g382(n1789 ,n18[0] ,n1770);
    nor g383(n1788 ,n248 ,n1679);
    nor g384(n1787 ,n251 ,n1677);
    nor g385(n1786 ,n247 ,n1676);
    nor g386(n1785 ,n1759 ,n1762);
    nor g387(n1784 ,n723 ,n1761);
    nor g388(n1783 ,n1760 ,n1763);
    or g389(n1782 ,n933 ,n1764);
    or g390(n1781 ,n927 ,n1741);
    or g391(n1780 ,n931 ,n1742);
    or g392(n1779 ,n932 ,n1740);
    or g393(n1778 ,n1751 ,n1738);
    or g394(n1777 ,n1752 ,n1737);
    or g395(n1776 ,n1750 ,n1739);
    or g396(n1775 ,n1753 ,n1745);
    or g397(n1774 ,n1754 ,n1746);
    or g398(n1773 ,n1755 ,n1747);
    or g399(n1772 ,n1756 ,n1748);
    or g400(n1771 ,n1703 ,n1702);
    or g401(n1769 ,n1661 ,n1660);
    or g402(n1768 ,n1662 ,n1278);
    or g403(n1767 ,n1664 ,n1663);
    nor g404(n1766 ,n247 ,n1486);
    nor g405(n1765 ,n250 ,n1495);
    nor g406(n1764 ,n45[0] ,n1643);
    nor g407(n1763 ,n570 ,n1641);
    nor g408(n1762 ,n670 ,n1641);
    nor g409(n1761 ,n263 ,n1642);
    nor g410(n1760 ,n265 ,n1642);
    nor g411(n1759 ,n413 ,n1642);
    nor g412(n1758 ,n268 ,n1644);
    nor g413(n1757 ,n533 ,n1640);
    nor g414(n1756 ,n288 ,n1640);
    nor g415(n1755 ,n343 ,n1640);
    nor g416(n1754 ,n310 ,n1640);
    nor g417(n1753 ,n489 ,n1640);
    nor g418(n1752 ,n301 ,n1640);
    nor g419(n1751 ,n309 ,n1640);
    nor g420(n1750 ,n327 ,n1640);
    nor g421(n1749 ,n430 ,n1639);
    nor g422(n1748 ,n420 ,n1639);
    nor g423(n1747 ,n421 ,n1639);
    nor g424(n1746 ,n427 ,n1639);
    nor g425(n1745 ,n428 ,n1639);
    nor g426(n1744 ,n432 ,n1644);
    nor g427(n1743 ,n431 ,n1644);
    nor g428(n1742 ,n358 ,n1643);
    nor g429(n1741 ,n364 ,n1643);
    nor g430(n1740 ,n367 ,n1643);
    nor g431(n1739 ,n437 ,n1639);
    nor g432(n1738 ,n424 ,n1639);
    nor g433(n1737 ,n422 ,n1639);
    or g434(n1770 ,n777 ,n1518);
    or g435(n1736 ,n1530 ,n1537);
    or g436(n1735 ,n1655 ,n1654);
    or g437(n1734 ,n1653 ,n1652);
    or g438(n1733 ,n1651 ,n1649);
    or g439(n1732 ,n1646 ,n1672);
    or g440(n1731 ,n1559 ,n1277);
    or g441(n1730 ,n1637 ,n1549);
    or g442(n1729 ,n1633 ,n1634);
    or g443(n1728 ,n1555 ,n1632);
    or g444(n1727 ,n1631 ,n1630);
    or g445(n1726 ,n1629 ,n1567);
    or g446(n1725 ,n1626 ,n1625);
    or g447(n1724 ,n1624 ,n1276);
    or g448(n1723 ,n1623 ,n1622);
    or g449(n1722 ,n1620 ,n1619);
    or g450(n1721 ,n1618 ,n1628);
    or g451(n1720 ,n1615 ,n1616);
    or g452(n1719 ,n1650 ,n1614);
    or g453(n1718 ,n1611 ,n1612);
    or g454(n1717 ,n1588 ,n1275);
    or g455(n1716 ,n1610 ,n1609);
    or g456(n1715 ,n1607 ,n1606);
    or g457(n1714 ,n1605 ,n1604);
    or g458(n1713 ,n1603 ,n1563);
    or g459(n1712 ,n1602 ,n1601);
    or g460(n1711 ,n1666 ,n1597);
    or g461(n1710 ,n1595 ,n1274);
    or g462(n1709 ,n1594 ,n1670);
    or g463(n1708 ,n1591 ,n1590);
    or g464(n1707 ,n1589 ,n1598);
    or g465(n1706 ,n1587 ,n1668);
    or g466(n1705 ,n1586 ,n1585);
    or g467(n1704 ,n1657 ,n1656);
    or g468(n1703 ,n1582 ,n1617);
    or g469(n1702 ,n1583 ,n1273);
    or g470(n1701 ,n1580 ,n1579);
    or g471(n1700 ,n1577 ,n1576);
    or g472(n1699 ,n1645 ,n1575);
    or g473(n1698 ,n1574 ,n1573);
    or g474(n1697 ,n1572 ,n1638);
    or g475(n1696 ,n1570 ,n1569);
    or g476(n1695 ,n1568 ,n1279);
    or g477(n1694 ,n1566 ,n1636);
    or g478(n1693 ,n1528 ,n1536);
    or g479(n1692 ,n1564 ,n1592);
    or g480(n1691 ,n1562 ,n1667);
    or g481(n1690 ,n1560 ,n1561);
    or g482(n1689 ,n1547 ,n1558);
    or g483(n1688 ,n1524 ,n1538);
    or g484(n1687 ,n1600 ,n1272);
    or g485(n1686 ,n1557 ,n1556);
    or g486(n1685 ,n1553 ,n1554);
    or g487(n1684 ,n1527 ,n1535);
    or g488(n1683 ,n1596 ,n1552);
    or g489(n1682 ,n1551 ,n1648);
    or g490(n1681 ,n1550 ,n1593);
    or g491(n1680 ,n1548 ,n1669);
    nor g492(n1679 ,n1522 ,n1516);
    or g493(n1678 ,n1529 ,n1534);
    nor g494(n1677 ,n1521 ,n1515);
    nor g495(n1676 ,n1519 ,n1514);
    or g496(n1675 ,n1526 ,n1533);
    or g497(n1674 ,n1525 ,n1532);
    or g498(n1673 ,n1523 ,n1531);
    nor g499(n1672 ,n285 ,n1470);
    nor g500(n1671 ,n345 ,n1466);
    nor g501(n1670 ,n562 ,n1467);
    nor g502(n1669 ,n456 ,n1473);
    nor g503(n1668 ,n332 ,n1475);
    nor g504(n1667 ,n505 ,n1477);
    nor g505(n1666 ,n503 ,n1471);
    nor g506(n1665 ,n450 ,n1472);
    nor g507(n1664 ,n311 ,n1471);
    nor g508(n1663 ,n474 ,n1470);
    nor g509(n1662 ,n472 ,n1469);
    nor g510(n1661 ,n492 ,n1468);
    nor g511(n1660 ,n502 ,n1467);
    nor g512(n1659 ,n487 ,n1466);
    nor g513(n1658 ,n464 ,n1466);
    nor g514(n1657 ,n346 ,n1480);
    nor g515(n1656 ,n525 ,n1479);
    nor g516(n1655 ,n463 ,n1478);
    nor g517(n1654 ,n320 ,n1477);
    nor g518(n1653 ,n500 ,n1476);
    nor g519(n1652 ,n493 ,n1475);
    nor g520(n1651 ,n353 ,n1474);
    nor g521(n1650 ,n445 ,n1474);
    nor g522(n1649 ,n567 ,n1473);
    nor g523(n1648 ,n552 ,n1477);
    nor g524(n1647 ,n548 ,n1472);
    nor g525(n1646 ,n468 ,n1471);
    nor g526(n1645 ,n448 ,n1478);
    not g527(n1642 ,n1641);
    not g528(n1639 ,n1640);
    nor g529(n1638 ,n284 ,n1473);
    nor g530(n1637 ,n527 ,n1468);
    nor g531(n1636 ,n352 ,n1467);
    nor g532(n1635 ,n317 ,n1466);
    nor g533(n1634 ,n458 ,n1479);
    nor g534(n1633 ,n561 ,n1480);
    nor g535(n1632 ,n514 ,n1477);
    nor g536(n1631 ,n319 ,n1476);
    nor g537(n1630 ,n295 ,n1475);
    nor g538(n1629 ,n556 ,n1474);
    nor g539(n1628 ,n315 ,n1477);
    nor g540(n1627 ,n541 ,n1472);
    nor g541(n1626 ,n287 ,n1471);
    nor g542(n1625 ,n512 ,n1470);
    nor g543(n1624 ,n334 ,n1469);
    nor g544(n1623 ,n566 ,n1468);
    nor g545(n1622 ,n335 ,n1467);
    nor g546(n1621 ,n328 ,n1466);
    nor g547(n1620 ,n547 ,n1480);
    nor g548(n1619 ,n522 ,n1479);
    nor g549(n1618 ,n447 ,n1478);
    nor g550(n1617 ,n304 ,n1470);
    nor g551(n1616 ,n313 ,n1475);
    nor g552(n1615 ,n554 ,n1476);
    nor g553(n1614 ,n351 ,n1473);
    nor g554(n1613 ,n282 ,n1472);
    nor g555(n1612 ,n483 ,n1470);
    nor g556(n1611 ,n507 ,n1471);
    nor g557(n1610 ,n465 ,n1468);
    nor g558(n1609 ,n442 ,n1467);
    nor g559(n1608 ,n496 ,n1466);
    nor g560(n1607 ,n481 ,n1480);
    nor g561(n1606 ,n330 ,n1479);
    nor g562(n1605 ,n469 ,n1478);
    nor g563(n1604 ,n312 ,n1477);
    nor g564(n1603 ,n337 ,n1476);
    nor g565(n1602 ,n516 ,n1474);
    nor g566(n1601 ,n488 ,n1473);
    nor g567(n1600 ,n520 ,n1469);
    nor g568(n1599 ,n302 ,n1472);
    nor g569(n1598 ,n560 ,n1477);
    nor g570(n1597 ,n350 ,n1470);
    nor g571(n1596 ,n336 ,n1480);
    nor g572(n1595 ,n497 ,n1469);
    nor g573(n1594 ,n333 ,n1468);
    nor g574(n1593 ,n308 ,n1475);
    nor g575(n1592 ,n307 ,n1479);
    nor g576(n1591 ,n543 ,n1480);
    nor g577(n1590 ,n532 ,n1479);
    nor g578(n1589 ,n449 ,n1478);
    nor g579(n1588 ,n523 ,n1469);
    nor g580(n1587 ,n477 ,n1476);
    nor g581(n1586 ,n293 ,n1474);
    nor g582(n1585 ,n557 ,n1473);
    nor g583(n1584 ,n453 ,n1472);
    nor g584(n1583 ,n524 ,n1469);
    nor g585(n1582 ,n283 ,n1471);
    nor g586(n1581 ,n509 ,n1472);
    nor g587(n1580 ,n339 ,n1468);
    nor g588(n1579 ,n321 ,n1467);
    nor g589(n1578 ,n286 ,n1466);
    nor g590(n1577 ,n529 ,n1480);
    nor g591(n1576 ,n316 ,n1479);
    nor g592(n1575 ,n569 ,n1477);
    nor g593(n1574 ,n538 ,n1476);
    nor g594(n1573 ,n545 ,n1475);
    nor g595(n1572 ,n326 ,n1474);
    nor g596(n1571 ,n324 ,n1472);
    nor g597(n1570 ,n478 ,n1471);
    nor g598(n1569 ,n521 ,n1470);
    nor g599(n1568 ,n349 ,n1469);
    nor g600(n1567 ,n555 ,n1473);
    nor g601(n1566 ,n451 ,n1468);
    nor g602(n1565 ,n455 ,n1466);
    nor g603(n1564 ,n537 ,n1480);
    nor g604(n1563 ,n470 ,n1475);
    nor g605(n1562 ,n322 ,n1478);
    nor g606(n1561 ,n347 ,n1475);
    nor g607(n1560 ,n279 ,n1476);
    nor g608(n1559 ,n559 ,n1469);
    nor g609(n1558 ,n452 ,n1473);
    nor g610(n1557 ,n348 ,n1471);
    nor g611(n1556 ,n318 ,n1470);
    nor g612(n1555 ,n526 ,n1478);
    nor g613(n1554 ,n528 ,n1467);
    nor g614(n1553 ,n331 ,n1468);
    nor g615(n1552 ,n490 ,n1479);
    nor g616(n1551 ,n289 ,n1478);
    nor g617(n1550 ,n486 ,n1476);
    nor g618(n1549 ,n511 ,n1467);
    nor g619(n1548 ,n549 ,n1474);
    nor g620(n1547 ,n550 ,n1474);
    nor g621(n1546 ,n540 ,n1465);
    nor g622(n1545 ,n534 ,n1465);
    nor g623(n1544 ,n531 ,n1465);
    nor g624(n1543 ,n544 ,n1465);
    nor g625(n1542 ,n501 ,n1465);
    nor g626(n1541 ,n563 ,n1465);
    nor g627(n1540 ,n444 ,n1465);
    nor g628(n1539 ,n499 ,n1465);
    nor g629(n1538 ,n422 ,n1462);
    nor g630(n1537 ,n437 ,n1462);
    nor g631(n1536 ,n424 ,n1462);
    nor g632(n1535 ,n428 ,n1462);
    nor g633(n1534 ,n427 ,n1462);
    nor g634(n1533 ,n421 ,n1462);
    nor g635(n1532 ,n420 ,n1462);
    nor g636(n1531 ,n430 ,n1462);
    nor g637(n1530 ,n564 ,n1463);
    nor g638(n1529 ,n459 ,n1463);
    nor g639(n1528 ,n292 ,n1463);
    nor g640(n1527 ,n306 ,n1463);
    nor g641(n1526 ,n281 ,n1463);
    nor g642(n1525 ,n476 ,n1463);
    nor g643(n1524 ,n480 ,n1463);
    nor g644(n1523 ,n443 ,n1463);
    nor g645(n1522 ,n417 ,n1481);
    nor g646(n1521 ,n418 ,n1481);
    or g647(n1520 ,n930 ,n1414);
    nor g648(n1519 ,n412 ,n1481);
    or g649(n1518 ,n664 ,n1484);
    or g650(n1517 ,n928 ,n1415);
    nor g651(n1516 ,n661 ,n1482);
    nor g652(n1515 ,n650 ,n1482);
    nor g653(n1514 ,n605 ,n1482);
    nor g654(n1513 ,n246 ,n1410);
    or g655(n1512 ,n912 ,n1416);
    nor g656(n1511 ,n245 ,n1342);
    nor g657(n1510 ,n249 ,n1341);
    nor g658(n1509 ,n249 ,n1311);
    nor g659(n1508 ,n247 ,n1306);
    nor g660(n1507 ,n249 ,n1301);
    nor g661(n1506 ,n246 ,n1296);
    or g662(n1505 ,n918 ,n1421);
    or g663(n1504 ,n920 ,n1423);
    or g664(n1503 ,n919 ,n1422);
    or g665(n1502 ,n917 ,n1420);
    or g666(n1501 ,n1412 ,n1407);
    or g667(n1500 ,n1426 ,n1437);
    or g668(n1499 ,n915 ,n1419);
    or g669(n1498 ,n1425 ,n1436);
    or g670(n1497 ,n1424 ,n1435);
    or g671(n1496 ,n913 ,n1461);
    nor g672(n1495 ,n1434 ,n1405);
    or g673(n1494 ,n1433 ,n1283);
    or g674(n1493 ,n1413 ,n995);
    or g675(n1492 ,n1432 ,n1282);
    or g676(n1491 ,n757 ,n1431);
    or g677(n1490 ,n737 ,n1430);
    or g678(n1489 ,n735 ,n1429);
    or g679(n1488 ,n736 ,n1428);
    or g680(n1487 ,n914 ,n1418);
    nor g681(n1486 ,n1408 ,n1427);
    or g682(n1485 ,n916 ,n1402);
    or g683(n1644 ,n253 ,n1483);
    or g684(n1643 ,n812 ,n1464);
    nor g685(n1641 ,n1291 ,n1406);
    nor g686(n1640 ,n585 ,n1409);
    not g687(n1484 ,n1483);
    not g688(n1481 ,n1482);
    not g689(n1465 ,n1464);
    not g690(n1462 ,n1463);
    nor g691(n1461 ,n366 ,n1127);
    or g692(n1460 ,n1241 ,n1095);
    or g693(n1459 ,n1242 ,n1096);
    or g694(n1458 ,n1243 ,n1097);
    or g695(n1457 ,n1244 ,n1099);
    or g696(n1456 ,n1245 ,n1100);
    or g697(n1455 ,n1247 ,n1115);
    or g698(n1454 ,n1246 ,n1101);
    or g699(n1453 ,n1248 ,n1103);
    or g700(n1452 ,n1250 ,n1105);
    or g701(n1451 ,n1251 ,n1106);
    or g702(n1450 ,n1252 ,n1107);
    or g703(n1449 ,n1253 ,n1108);
    or g704(n1448 ,n1173 ,n1022);
    or g705(n1447 ,n1254 ,n1109);
    or g706(n1446 ,n1255 ,n1110);
    or g707(n1445 ,n1159 ,n1075);
    or g708(n1444 ,n1256 ,n1112);
    or g709(n1443 ,n1257 ,n1113);
    or g710(n1442 ,n1258 ,n1114);
    or g711(n1441 ,n1259 ,n1116);
    or g712(n1440 ,n1260 ,n1117);
    or g713(n1439 ,n1261 ,n1119);
    or g714(n1438 ,n1262 ,n1120);
    nor g715(n1437 ,n410 ,n1131);
    nor g716(n1436 ,n382 ,n1131);
    nor g717(n1435 ,n404 ,n1131);
    nor g718(n1434 ,n436 ,n1138);
    nor g719(n1433 ,n274 ,n1134);
    nor g720(n1432 ,n273 ,n1134);
    nor g721(n1431 ,n383 ,n1132);
    nor g722(n1430 ,n379 ,n1132);
    nor g723(n1429 ,n405 ,n1132);
    nor g724(n1428 ,n378 ,n1132);
    nor g725(n1427 ,n434 ,n1136);
    nor g726(n1426 ,n423 ,n1129);
    nor g727(n1425 ,n429 ,n1129);
    nor g728(n1424 ,n426 ,n1129);
    nor g729(n1423 ,n400 ,n1127);
    nor g730(n1422 ,n407 ,n1127);
    nor g731(n1421 ,n391 ,n1127);
    nor g732(n1420 ,n369 ,n1127);
    nor g733(n1419 ,n384 ,n1127);
    nor g734(n1418 ,n359 ,n1127);
    or g735(n1417 ,n1264 ,n1121);
    nor g736(n1416 ,n360 ,n1127);
    nor g737(n1415 ,n385 ,n1127);
    nor g738(n1414 ,n393 ,n1127);
    nor g739(n1413 ,n416 ,n1134);
    nor g740(n1412 ,n419 ,n1129);
    or g741(n1411 ,n1239 ,n1093);
    nor g742(n1410 ,n1263 ,n1271);
    or g743(n1409 ,n576 ,n992);
    nor g744(n1408 ,n265 ,n1135);
    nor g745(n1407 ,n23[0] ,n1131);
    nor g746(n1406 ,n652 ,n997);
    nor g747(n1405 ,n601 ,n1137);
    or g748(n1404 ,n1265 ,n1122);
    or g749(n1403 ,n1240 ,n1094);
    nor g750(n1402 ,n17[0] ,n1127);
    nor g751(n1401 ,n248 ,n993);
    or g752(n1400 ,n1266 ,n1123);
    nor g753(n1483 ,n720 ,n994);
    nor g754(n1482 ,n901 ,n996);
    or g755(n1480 ,n597 ,n1130);
    or g756(n1479 ,n589 ,n1130);
    or g757(n1478 ,n589 ,n1292);
    or g758(n1477 ,n596 ,n1133);
    or g759(n1476 ,n597 ,n1293);
    or g760(n1475 ,n589 ,n1293);
    or g761(n1474 ,n597 ,n1133);
    or g762(n1473 ,n589 ,n1133);
    or g763(n1472 ,n590 ,n1133);
    or g764(n1471 ,n590 ,n1293);
    or g765(n1470 ,n596 ,n1293);
    or g766(n1469 ,n597 ,n1292);
    or g767(n1468 ,n590 ,n1130);
    or g768(n1467 ,n596 ,n1130);
    or g769(n1466 ,n596 ,n1292);
    nor g770(n1464 ,n590 ,n1292);
    nor g771(n1463 ,n770 ,n1128);
    or g772(n1399 ,n1184 ,n1002);
    or g773(n1398 ,n1237 ,n1090);
    or g774(n1397 ,n1236 ,n1089);
    or g775(n1396 ,n1249 ,n1098);
    or g776(n1395 ,n1235 ,n1088);
    or g777(n1394 ,n1234 ,n1087);
    or g778(n1393 ,n1233 ,n1086);
    or g779(n1392 ,n1229 ,n1111);
    or g780(n1391 ,n1228 ,n1085);
    or g781(n1390 ,n1227 ,n1083);
    or g782(n1389 ,n1232 ,n1081);
    or g783(n1388 ,n1226 ,n1082);
    or g784(n1387 ,n1225 ,n1092);
    or g785(n1386 ,n1224 ,n1044);
    or g786(n1385 ,n1223 ,n1080);
    or g787(n1384 ,n1222 ,n1079);
    or g788(n1383 ,n1221 ,n1078);
    or g789(n1382 ,n1220 ,n1077);
    or g790(n1381 ,n1219 ,n1076);
    or g791(n1380 ,n1218 ,n1074);
    or g792(n1379 ,n1217 ,n1042);
    or g793(n1378 ,n1179 ,n1031);
    or g794(n1377 ,n1216 ,n1072);
    or g795(n1376 ,n1214 ,n1070);
    or g796(n1375 ,n1213 ,n1069);
    or g797(n1374 ,n1212 ,n1068);
    or g798(n1373 ,n1211 ,n1084);
    or g799(n1372 ,n1210 ,n1066);
    or g800(n1371 ,n1209 ,n1065);
    or g801(n1370 ,n1207 ,n1063);
    or g802(n1369 ,n1208 ,n1064);
    or g803(n1368 ,n1206 ,n1062);
    or g804(n1367 ,n1205 ,n1061);
    or g805(n1366 ,n1204 ,n1060);
    or g806(n1365 ,n1203 ,n1059);
    or g807(n1364 ,n1202 ,n1058);
    or g808(n1363 ,n1201 ,n1057);
    or g809(n1362 ,n1200 ,n1028);
    or g810(n1361 ,n1199 ,n1055);
    or g811(n1360 ,n1198 ,n1027);
    or g812(n1359 ,n1197 ,n1054);
    or g813(n1358 ,n1196 ,n1053);
    or g814(n1357 ,n1195 ,n1052);
    or g815(n1356 ,n1194 ,n1051);
    or g816(n1355 ,n1193 ,n1050);
    or g817(n1354 ,n1192 ,n1049);
    or g818(n1353 ,n1191 ,n1048);
    or g819(n1352 ,n1190 ,n1047);
    or g820(n1351 ,n1189 ,n1046);
    or g821(n1350 ,n1188 ,n1006);
    or g822(n1349 ,n1187 ,n1005);
    or g823(n1348 ,n1186 ,n1004);
    or g824(n1347 ,n1185 ,n1003);
    or g825(n1346 ,n1238 ,n1091);
    or g826(n1345 ,n1183 ,n1001);
    or g827(n1344 ,n1182 ,n1000);
    or g828(n1343 ,n1181 ,n999);
    nor g829(n1342 ,n1126 ,n1281);
    nor g830(n1341 ,n1290 ,n1280);
    or g831(n1340 ,n1230 ,n1104);
    or g832(n1339 ,n1178 ,n1056);
    or g833(n1338 ,n1176 ,n1067);
    or g834(n1337 ,n1174 ,n1033);
    or g835(n1336 ,n1175 ,n1073);
    or g836(n1335 ,n1177 ,n1045);
    or g837(n1334 ,n1172 ,n1039);
    or g838(n1333 ,n1171 ,n1038);
    or g839(n1332 ,n1163 ,n1118);
    or g840(n1331 ,n1170 ,n1036);
    or g841(n1330 ,n1166 ,n1035);
    or g842(n1329 ,n1155 ,n1034);
    or g843(n1328 ,n1168 ,n1037);
    or g844(n1327 ,n1167 ,n1032);
    or g845(n1326 ,n1215 ,n1026);
    or g846(n1325 ,n1165 ,n1102);
    or g847(n1324 ,n1164 ,n998);
    or g848(n1323 ,n1231 ,n1043);
    or g849(n1322 ,n1169 ,n1030);
    or g850(n1321 ,n1180 ,n1029);
    or g851(n1320 ,n1157 ,n1025);
    or g852(n1319 ,n1158 ,n1024);
    or g853(n1318 ,n1160 ,n1071);
    or g854(n1317 ,n1162 ,n1041);
    or g855(n1316 ,n1161 ,n1040);
    or g856(n1315 ,n1156 ,n1124);
    or g857(n1314 ,n1154 ,n1023);
    or g858(n1313 ,n1153 ,n1021);
    or g859(n1312 ,n1152 ,n1020);
    nor g860(n1311 ,n1150 ,n1270);
    or g861(n1310 ,n1151 ,n1019);
    or g862(n1309 ,n1149 ,n1018);
    or g863(n1308 ,n1148 ,n1017);
    or g864(n1307 ,n1147 ,n1016);
    nor g865(n1306 ,n1145 ,n1269);
    or g866(n1305 ,n1146 ,n1015);
    or g867(n1304 ,n1144 ,n1014);
    or g868(n1303 ,n1143 ,n1013);
    or g869(n1302 ,n1142 ,n1012);
    nor g870(n1301 ,n1140 ,n1268);
    or g871(n1300 ,n1141 ,n1011);
    or g872(n1299 ,n1139 ,n1010);
    or g873(n1298 ,n1284 ,n1009);
    or g874(n1297 ,n1285 ,n1008);
    nor g875(n1296 ,n1287 ,n1267);
    or g876(n1295 ,n1286 ,n1007);
    or g877(n1294 ,n1288 ,n1125);
    nor g878(n1291 ,n263 ,n876);
    nor g879(n1290 ,n412 ,n910);
    or g880(n1289 ,n644 ,n887);
    nor g881(n1288 ,n526 ,n950);
    nor g882(n1287 ,n446 ,n904);
    nor g883(n1286 ,n463 ,n950);
    nor g884(n1285 ,n336 ,n938);
    nor g885(n1284 ,n537 ,n938);
    nor g886(n1283 ,n354 ,n908);
    nor g887(n1282 ,n375 ,n908);
    nor g888(n1281 ,n440 ,n907);
    nor g889(n1280 ,n439 ,n911);
    nor g890(n1279 ,n539 ,n905);
    nor g891(n1278 ,n467 ,n905);
    nor g892(n1277 ,n558 ,n905);
    nor g893(n1276 ,n508 ,n905);
    nor g894(n1275 ,n338 ,n905);
    nor g895(n1274 ,n506 ,n905);
    nor g896(n1273 ,n568 ,n905);
    nor g897(n1272 ,n504 ,n905);
    nor g898(n1271 ,n399 ,n903);
    nor g899(n1270 ,n395 ,n903);
    nor g900(n1269 ,n356 ,n903);
    nor g901(n1268 ,n372 ,n903);
    nor g902(n1267 ,n380 ,n903);
    nor g903(n1266 ,n447 ,n950);
    nor g904(n1265 ,n469 ,n950);
    nor g905(n1264 ,n449 ,n950);
    nor g906(n1262 ,n448 ,n950);
    nor g907(n1261 ,n322 ,n950);
    nor g908(n1260 ,n289 ,n950);
    nor g909(n1259 ,n472 ,n966);
    nor g910(n1258 ,n559 ,n966);
    nor g911(n1257 ,n334 ,n966);
    nor g912(n1256 ,n523 ,n966);
    nor g913(n1255 ,n497 ,n966);
    nor g914(n1254 ,n524 ,n966);
    nor g915(n1253 ,n349 ,n966);
    nor g916(n1252 ,n520 ,n966);
    nor g917(n1251 ,n320 ,n964);
    nor g918(n1250 ,n514 ,n964);
    nor g919(n1249 ,n557 ,n948);
    nor g920(n1248 ,n315 ,n964);
    nor g921(n1247 ,n284 ,n948);
    nor g922(n1246 ,n312 ,n964);
    nor g923(n1245 ,n560 ,n964);
    nor g924(n1244 ,n569 ,n964);
    nor g925(n1243 ,n505 ,n964);
    nor g926(n1242 ,n552 ,n964);
    nor g927(n1241 ,n450 ,n962);
    nor g928(n1240 ,n548 ,n962);
    nor g929(n1239 ,n541 ,n962);
    nor g930(n1238 ,n282 ,n962);
    nor g931(n1237 ,n302 ,n962);
    nor g932(n1236 ,n453 ,n962);
    nor g933(n1235 ,n324 ,n962);
    nor g934(n1234 ,n509 ,n962);
    nor g935(n1233 ,n474 ,n960);
    nor g936(n1232 ,n488 ,n948);
    nor g937(n1231 ,n493 ,n940);
    nor g938(n1230 ,n295 ,n940);
    nor g939(n1229 ,n285 ,n960);
    nor g940(n1228 ,n512 ,n960);
    nor g941(n1227 ,n483 ,n960);
    nor g942(n1226 ,n350 ,n960);
    nor g943(n1225 ,n304 ,n960);
    nor g944(n1224 ,n500 ,n944);
    nor g945(n1223 ,n521 ,n960);
    nor g946(n1222 ,n318 ,n960);
    nor g947(n1221 ,n311 ,n958);
    nor g948(n1220 ,n468 ,n958);
    nor g949(n1219 ,n287 ,n958);
    nor g950(n1218 ,n507 ,n958);
    nor g951(n1217 ,n503 ,n958);
    nor g952(n1216 ,n283 ,n958);
    nor g953(n1215 ,n279 ,n944);
    nor g954(n1214 ,n478 ,n958);
    nor g955(n1213 ,n348 ,n958);
    nor g956(n1212 ,n502 ,n952);
    nor g957(n1211 ,n511 ,n952);
    nor g958(n1210 ,n335 ,n952);
    nor g959(n1209 ,n442 ,n952);
    nor g960(n1208 ,n562 ,n952);
    nor g961(n1207 ,n321 ,n952);
    nor g962(n1206 ,n352 ,n952);
    nor g963(n1205 ,n528 ,n952);
    nor g964(n1204 ,n492 ,n956);
    nor g965(n1203 ,n527 ,n956);
    nor g966(n1202 ,n566 ,n956);
    nor g967(n1201 ,n465 ,n956);
    nor g968(n1200 ,n333 ,n956);
    nor g969(n1199 ,n339 ,n956);
    nor g970(n1198 ,n451 ,n956);
    nor g971(n1197 ,n331 ,n956);
    nor g972(n1196 ,n464 ,n954);
    nor g973(n1195 ,n317 ,n954);
    nor g974(n1194 ,n328 ,n954);
    nor g975(n1193 ,n496 ,n954);
    nor g976(n1192 ,n345 ,n954);
    nor g977(n1191 ,n286 ,n954);
    nor g978(n1190 ,n455 ,n954);
    nor g979(n1189 ,n487 ,n954);
    nor g980(n1188 ,n540 ,n936);
    nor g981(n1187 ,n534 ,n936);
    nor g982(n1186 ,n531 ,n936);
    nor g983(n1185 ,n544 ,n936);
    nor g984(n1184 ,n501 ,n936);
    nor g985(n1183 ,n563 ,n936);
    nor g986(n1182 ,n444 ,n936);
    nor g987(n1181 ,n499 ,n936);
    nor g988(n1180 ,n470 ,n940);
    nor g989(n1179 ,n554 ,n944);
    nor g990(n1178 ,n567 ,n948);
    nor g991(n1177 ,n337 ,n944);
    nor g992(n1176 ,n555 ,n948);
    nor g993(n1175 ,n351 ,n948);
    nor g994(n1174 ,n293 ,n946);
    nor g995(n1173 ,n452 ,n948);
    nor g996(n1172 ,n456 ,n948);
    nor g997(n1171 ,n353 ,n946);
    nor g998(n1170 ,n556 ,n946);
    nor g999(n1169 ,n313 ,n940);
    nor g1000(n1168 ,n516 ,n946);
    nor g1001(n1167 ,n326 ,n946);
    nor g1002(n1166 ,n445 ,n946);
    nor g1003(n1165 ,n550 ,n946);
    nor g1004(n1164 ,n549 ,n946);
    nor g1005(n1163 ,n486 ,n944);
    nor g1006(n1162 ,n538 ,n944);
    nor g1007(n1161 ,n545 ,n940);
    nor g1008(n1160 ,n347 ,n940);
    nor g1009(n1159 ,n308 ,n940);
    nor g1010(n1158 ,n525 ,n942);
    nor g1011(n1157 ,n332 ,n940);
    nor g1012(n1156 ,n319 ,n944);
    nor g1013(n1155 ,n477 ,n944);
    nor g1014(n1154 ,n458 ,n942);
    nor g1015(n1153 ,n522 ,n942);
    nor g1016(n1152 ,n330 ,n942);
    nor g1017(n1151 ,n532 ,n942);
    nor g1018(n1150 ,n536 ,n904);
    nor g1019(n1149 ,n316 ,n942);
    nor g1020(n1148 ,n307 ,n942);
    nor g1021(n1147 ,n490 ,n942);
    nor g1022(n1146 ,n346 ,n938);
    nor g1023(n1145 ,n341 ,n904);
    nor g1024(n1144 ,n561 ,n938);
    nor g1025(n1143 ,n547 ,n938);
    nor g1026(n1142 ,n481 ,n938);
    nor g1027(n1141 ,n543 ,n938);
    nor g1028(n1140 ,n325 ,n904);
    nor g1029(n1139 ,n529 ,n938);
    or g1030(n1293 ,n415 ,n909);
    or g1031(n1292 ,n415 ,n967);
    not g1032(n1138 ,n1137);
    not g1033(n1136 ,n1135);
    not g1034(n1129 ,n1128);
    nor g1035(n1126 ,n48[2] ,n906);
    nor g1036(n1125 ,n261 ,n949);
    nor g1037(n1124 ,n261 ,n943);
    nor g1038(n1123 ,n260 ,n949);
    nor g1039(n1122 ,n257 ,n949);
    nor g1040(n1121 ,n262 ,n949);
    nor g1041(n1120 ,n255 ,n949);
    nor g1042(n1119 ,n258 ,n949);
    nor g1043(n1118 ,n259 ,n943);
    nor g1044(n1117 ,n259 ,n949);
    nor g1045(n1116 ,n256 ,n965);
    nor g1046(n1115 ,n255 ,n947);
    nor g1047(n1114 ,n261 ,n965);
    nor g1048(n1113 ,n260 ,n965);
    nor g1049(n1112 ,n257 ,n965);
    nor g1050(n1111 ,n261 ,n959);
    nor g1051(n1110 ,n262 ,n965);
    nor g1052(n1109 ,n255 ,n965);
    nor g1053(n1108 ,n258 ,n965);
    nor g1054(n1107 ,n259 ,n965);
    nor g1055(n1106 ,n256 ,n963);
    nor g1056(n1105 ,n261 ,n963);
    nor g1057(n1104 ,n261 ,n939);
    nor g1058(n1103 ,n260 ,n963);
    nor g1059(n1102 ,n258 ,n945);
    nor g1060(n1101 ,n257 ,n963);
    nor g1061(n1100 ,n262 ,n963);
    nor g1062(n1099 ,n255 ,n963);
    nor g1063(n1098 ,n262 ,n947);
    nor g1064(n1097 ,n258 ,n963);
    nor g1065(n1096 ,n259 ,n963);
    nor g1066(n1095 ,n256 ,n961);
    nor g1067(n1094 ,n261 ,n961);
    nor g1068(n1093 ,n260 ,n961);
    nor g1069(n1092 ,n255 ,n959);
    nor g1070(n1091 ,n257 ,n961);
    nor g1071(n1090 ,n262 ,n961);
    nor g1072(n1089 ,n255 ,n961);
    nor g1073(n1088 ,n258 ,n961);
    nor g1074(n1087 ,n259 ,n961);
    nor g1075(n1086 ,n256 ,n959);
    nor g1076(n1085 ,n260 ,n959);
    nor g1077(n1084 ,n261 ,n951);
    nor g1078(n1083 ,n257 ,n959);
    nor g1079(n1082 ,n262 ,n959);
    nor g1080(n1081 ,n257 ,n947);
    nor g1081(n1080 ,n258 ,n959);
    nor g1082(n1079 ,n259 ,n959);
    nor g1083(n1078 ,n256 ,n957);
    nor g1084(n1077 ,n261 ,n957);
    nor g1085(n1076 ,n260 ,n957);
    nor g1086(n1075 ,n259 ,n939);
    nor g1087(n1074 ,n257 ,n957);
    nor g1088(n1073 ,n260 ,n947);
    nor g1089(n1072 ,n255 ,n957);
    nor g1090(n1071 ,n258 ,n939);
    nor g1091(n1070 ,n258 ,n957);
    nor g1092(n1069 ,n259 ,n957);
    nor g1093(n1068 ,n256 ,n951);
    nor g1094(n1067 ,n261 ,n947);
    nor g1095(n1066 ,n260 ,n951);
    nor g1096(n1065 ,n257 ,n951);
    nor g1097(n1064 ,n262 ,n951);
    nor g1098(n1063 ,n255 ,n951);
    nor g1099(n1062 ,n258 ,n951);
    nor g1100(n1061 ,n259 ,n951);
    nor g1101(n1060 ,n256 ,n955);
    nor g1102(n1059 ,n261 ,n955);
    nor g1103(n1058 ,n260 ,n955);
    nor g1104(n1057 ,n257 ,n955);
    nor g1105(n1056 ,n256 ,n947);
    nor g1106(n1055 ,n255 ,n955);
    nor g1107(n1054 ,n259 ,n955);
    nor g1108(n1053 ,n256 ,n953);
    nor g1109(n1052 ,n261 ,n953);
    nor g1110(n1051 ,n260 ,n953);
    nor g1111(n1050 ,n257 ,n953);
    nor g1112(n1049 ,n262 ,n953);
    nor g1113(n1048 ,n255 ,n953);
    nor g1114(n1047 ,n258 ,n953);
    nor g1115(n1046 ,n259 ,n953);
    nor g1116(n1045 ,n257 ,n943);
    nor g1117(n1044 ,n256 ,n943);
    nor g1118(n1043 ,n256 ,n939);
    nor g1119(n1042 ,n262 ,n957);
    nor g1120(n1041 ,n255 ,n943);
    nor g1121(n1040 ,n255 ,n939);
    nor g1122(n1039 ,n259 ,n947);
    nor g1123(n1038 ,n256 ,n945);
    nor g1124(n1037 ,n257 ,n945);
    nor g1125(n1036 ,n261 ,n945);
    nor g1126(n1035 ,n260 ,n945);
    nor g1127(n1034 ,n262 ,n943);
    nor g1128(n1033 ,n262 ,n945);
    nor g1129(n1032 ,n255 ,n945);
    nor g1130(n1031 ,n260 ,n943);
    nor g1131(n1030 ,n260 ,n939);
    nor g1132(n1029 ,n257 ,n939);
    nor g1133(n1028 ,n262 ,n955);
    nor g1134(n1027 ,n258 ,n955);
    nor g1135(n1026 ,n258 ,n943);
    nor g1136(n1025 ,n262 ,n939);
    nor g1137(n1024 ,n256 ,n941);
    nor g1138(n1023 ,n261 ,n941);
    nor g1139(n1022 ,n258 ,n947);
    nor g1140(n1021 ,n260 ,n941);
    nor g1141(n1020 ,n257 ,n941);
    nor g1142(n1019 ,n262 ,n941);
    nor g1143(n1018 ,n255 ,n941);
    nor g1144(n1017 ,n258 ,n941);
    nor g1145(n1016 ,n259 ,n941);
    nor g1146(n1015 ,n256 ,n937);
    nor g1147(n1014 ,n261 ,n937);
    nor g1148(n1013 ,n260 ,n937);
    nor g1149(n1012 ,n257 ,n937);
    nor g1150(n1011 ,n262 ,n937);
    nor g1151(n1010 ,n255 ,n937);
    nor g1152(n1009 ,n258 ,n937);
    nor g1153(n1008 ,n259 ,n937);
    nor g1154(n1007 ,n256 ,n949);
    nor g1155(n1006 ,n256 ,n935);
    nor g1156(n1005 ,n261 ,n935);
    nor g1157(n1004 ,n260 ,n935);
    nor g1158(n1003 ,n257 ,n935);
    nor g1159(n1002 ,n262 ,n935);
    nor g1160(n1001 ,n255 ,n935);
    nor g1161(n1000 ,n258 ,n935);
    nor g1162(n999 ,n259 ,n935);
    nor g1163(n998 ,n259 ,n945);
    or g1164(n997 ,n25[1] ,n899);
    or g1165(n996 ,n662 ,n907);
    nor g1166(n995 ,n27[0] ,n908);
    nor g1167(n994 ,n25[1] ,n872);
    nor g1168(n993 ,n14[1] ,n929);
    or g1169(n992 ,n23[0] ,n903);
    nor g1170(n991 ,n251 ,n886);
    nor g1171(n990 ,n245 ,n878);
    nor g1172(n989 ,n250 ,n882);
    nor g1173(n988 ,n246 ,n881);
    nor g1174(n987 ,n245 ,n880);
    nor g1175(n986 ,n250 ,n902);
    nor g1176(n985 ,n249 ,n879);
    nor g1177(n984 ,n245 ,n883);
    nor g1178(n983 ,n251 ,n875);
    nor g1179(n982 ,n248 ,n885);
    nor g1180(n981 ,n246 ,n873);
    nor g1181(n980 ,n245 ,n871);
    nor g1182(n979 ,n245 ,n870);
    nor g1183(n978 ,n250 ,n869);
    nor g1184(n977 ,n249 ,n868);
    nor g1185(n976 ,n250 ,n867);
    nor g1186(n975 ,n248 ,n866);
    nor g1187(n974 ,n249 ,n865);
    nor g1188(n973 ,n251 ,n864);
    nor g1189(n972 ,n248 ,n863);
    nor g1190(n971 ,n248 ,n862);
    nor g1191(n970 ,n248 ,n861);
    nor g1192(n969 ,n250 ,n860);
    nor g1193(n968 ,n249 ,n859);
    nor g1194(n1137 ,n710 ,n892);
    nor g1195(n1135 ,n669 ,n904);
    or g1196(n1134 ,n252 ,n877);
    or g1197(n1133 ,n45[1] ,n909);
    or g1198(n1131 ,n731 ,n903);
    or g1199(n1130 ,n45[1] ,n967);
    nor g1200(n1128 ,n245 ,n904);
    or g1201(n1127 ,n793 ,n897);
    not g1202(n965 ,n966);
    not g1203(n963 ,n964);
    not g1204(n961 ,n962);
    not g1205(n959 ,n960);
    not g1206(n957 ,n958);
    not g1207(n955 ,n956);
    not g1208(n953 ,n954);
    not g1209(n951 ,n952);
    not g1210(n949 ,n950);
    not g1211(n947 ,n948);
    not g1212(n945 ,n946);
    not g1213(n943 ,n944);
    not g1214(n941 ,n942);
    not g1215(n939 ,n940);
    not g1216(n937 ,n938);
    not g1217(n935 ,n936);
    nor g1218(n934 ,n504 ,n806);
    nor g1219(n933 ,n266 ,n807);
    nor g1220(n932 ,n414 ,n807);
    nor g1221(n931 ,n415 ,n807);
    nor g1222(n930 ,n298 ,n804);
    nor g1223(n929 ,n275 ,n816);
    nor g1224(n928 ,n542 ,n804);
    nor g1225(n927 ,n425 ,n807);
    nor g1226(n926 ,n508 ,n806);
    nor g1227(n925 ,n558 ,n806);
    nor g1228(n924 ,n506 ,n806);
    nor g1229(n923 ,n568 ,n806);
    nor g1230(n922 ,n338 ,n806);
    nor g1231(n921 ,n539 ,n806);
    nor g1232(n920 ,n462 ,n804);
    nor g1233(n919 ,n329 ,n804);
    nor g1234(n918 ,n297 ,n804);
    nor g1235(n917 ,n535 ,n804);
    nor g1236(n916 ,n433 ,n804);
    nor g1237(n915 ,n303 ,n804);
    nor g1238(n914 ,n290 ,n804);
    nor g1239(n913 ,n530 ,n804);
    nor g1240(n912 ,n471 ,n804);
    or g1241(n967 ,n425 ,n812);
    nor g1242(n966 ,n598 ,n811);
    nor g1243(n964 ,n594 ,n809);
    nor g1244(n962 ,n594 ,n810);
    nor g1245(n960 ,n595 ,n809);
    nor g1246(n958 ,n595 ,n810);
    nor g1247(n956 ,n591 ,n810);
    nor g1248(n954 ,n598 ,n809);
    nor g1249(n952 ,n591 ,n809);
    nor g1250(n950 ,n598 ,n808);
    nor g1251(n948 ,n594 ,n808);
    nor g1252(n946 ,n594 ,n811);
    nor g1253(n944 ,n595 ,n811);
    nor g1254(n942 ,n591 ,n808);
    nor g1255(n940 ,n595 ,n808);
    nor g1256(n938 ,n591 ,n811);
    nor g1257(n936 ,n598 ,n810);
    not g1258(n911 ,n910);
    not g1259(n907 ,n906);
    not g1260(n903 ,n904);
    nor g1261(n902 ,n832 ,n840);
    nor g1262(n901 ,n254 ,n799);
    or g1263(n900 ,n675 ,n850);
    nor g1264(n899 ,n25[0] ,n815);
    or g1265(n898 ,n747 ,n801);
    nor g1266(n897 ,n571 ,n779);
    or g1267(n896 ,n749 ,n781);
    or g1268(n895 ,n746 ,n769);
    or g1269(n894 ,n691 ,n852);
    or g1270(n893 ,n751 ,n778);
    nor g1271(n892 ,n593 ,n814);
    or g1272(n891 ,n759 ,n798);
    or g1273(n890 ,n752 ,n800);
    or g1274(n889 ,n753 ,n767);
    or g1275(n888 ,n739 ,n802);
    or g1276(n887 ,n758 ,n849);
    nor g1277(n886 ,n830 ,n836);
    nor g1278(n885 ,n823 ,n792);
    or g1279(n884 ,n689 ,n851);
    nor g1280(n883 ,n858 ,n838);
    nor g1281(n882 ,n826 ,n837);
    nor g1282(n881 ,n834 ,n842);
    nor g1283(n880 ,n833 ,n841);
    nor g1284(n879 ,n831 ,n839);
    nor g1285(n878 ,n825 ,n843);
    nor g1286(n877 ,n254 ,n780);
    nor g1287(n876 ,n25[2] ,n821);
    nor g1288(n875 ,n857 ,n788);
    or g1289(n874 ,n686 ,n853);
    nor g1290(n873 ,n856 ,n783);
    nor g1291(n872 ,n721 ,n768);
    nor g1292(n871 ,n829 ,n785);
    nor g1293(n870 ,n828 ,n782);
    nor g1294(n869 ,n855 ,n784);
    nor g1295(n868 ,n827 ,n791);
    nor g1296(n867 ,n854 ,n786);
    nor g1297(n866 ,n835 ,n790);
    nor g1298(n865 ,n817 ,n789);
    nor g1299(n864 ,n818 ,n787);
    nor g1300(n863 ,n819 ,n844);
    nor g1301(n862 ,n820 ,n847);
    nor g1302(n861 ,n824 ,n845);
    nor g1303(n860 ,n822 ,n846);
    nor g1304(n859 ,n803 ,n848);
    nor g1305(n910 ,n660 ,n813);
    or g1306(n909 ,n45[2] ,n812);
    or g1307(n908 ,n572 ,n776);
    nor g1308(n906 ,n763 ,n813);
    or g1309(n905 ,n805 ,n807);
    nor g1310(n904 ,n21[4] ,n816);
    nor g1311(n858 ,n420 ,n761);
    nor g1312(n857 ,n438 ,n726);
    nor g1313(n856 ,n551 ,n726);
    nor g1314(n855 ,n441 ,n726);
    nor g1315(n854 ,n546 ,n726);
    nor g1316(n853 ,n371 ,n727);
    nor g1317(n852 ,n381 ,n727);
    nor g1318(n851 ,n355 ,n727);
    nor g1319(n850 ,n373 ,n727);
    nor g1320(n849 ,n467 ,n734);
    nor g1321(n848 ,n408 ,n762);
    nor g1322(n847 ,n374 ,n762);
    nor g1323(n846 ,n401 ,n762);
    nor g1324(n845 ,n388 ,n762);
    nor g1325(n844 ,n398 ,n762);
    nor g1326(n843 ,n420 ,n760);
    nor g1327(n842 ,n422 ,n760);
    nor g1328(n841 ,n428 ,n760);
    nor g1329(n840 ,n427 ,n760);
    nor g1330(n839 ,n421 ,n760);
    nor g1331(n838 ,n430 ,n760);
    nor g1332(n837 ,n424 ,n760);
    nor g1333(n836 ,n276 ,n760);
    nor g1334(n835 ,n294 ,n726);
    nor g1335(n834 ,n424 ,n761);
    nor g1336(n833 ,n422 ,n761);
    nor g1337(n832 ,n428 ,n761);
    nor g1338(n831 ,n427 ,n761);
    nor g1339(n830 ,n430 ,n761);
    nor g1340(n829 ,n466 ,n726);
    nor g1341(n828 ,n461 ,n726);
    nor g1342(n827 ,n299 ,n726);
    nor g1343(n826 ,n437 ,n761);
    nor g1344(n825 ,n421 ,n761);
    nor g1345(n824 ,n300 ,n763);
    nor g1346(n823 ,n475 ,n726);
    nor g1347(n822 ,n479 ,n763);
    nor g1348(n821 ,n272 ,n703);
    nor g1349(n820 ,n517 ,n763);
    nor g1350(n819 ,n518 ,n763);
    nor g1351(n818 ,n482 ,n726);
    nor g1352(n817 ,n305 ,n726);
    not g1353(n815 ,n814);
    not g1354(n806 ,n805);
    nor g1355(n803 ,n553 ,n763);
    or g1356(n802 ,n679 ,n750);
    or g1357(n801 ,n676 ,n741);
    or g1358(n800 ,n678 ,n743);
    nor g1359(n799 ,n48[0] ,n722);
    or g1360(n798 ,n681 ,n744);
    nor g1361(n797 ,n251 ,n712);
    nor g1362(n796 ,n246 ,n756);
    nor g1363(n795 ,n249 ,n716);
    nor g1364(n794 ,n247 ,n754);
    or g1365(n793 ,n252 ,n733);
    nor g1366(n792 ,n614 ,n725);
    nor g1367(n791 ,n617 ,n725);
    nor g1368(n790 ,n609 ,n725);
    nor g1369(n789 ,n612 ,n725);
    nor g1370(n788 ,n577 ,n725);
    nor g1371(n787 ,n574 ,n725);
    nor g1372(n786 ,n608 ,n725);
    nor g1373(n785 ,n615 ,n725);
    nor g1374(n784 ,n632 ,n725);
    nor g1375(n783 ,n627 ,n725);
    nor g1376(n782 ,n613 ,n725);
    or g1377(n781 ,n687 ,n748);
    nor g1378(n780 ,n715 ,n729);
    nor g1379(n779 ,n646 ,n718);
    or g1380(n778 ,n684 ,n738);
    or g1381(n777 ,n252 ,n745);
    nor g1382(n776 ,n713 ,n729);
    nor g1383(n775 ,n250 ,n714);
    nor g1384(n774 ,n247 ,n709);
    nor g1385(n773 ,n246 ,n704);
    nor g1386(n772 ,n247 ,n705);
    nor g1387(n771 ,n247 ,n719);
    or g1388(n770 ,n253 ,n730);
    or g1389(n769 ,n680 ,n742);
    nor g1390(n768 ,n25[0] ,n717);
    or g1391(n767 ,n677 ,n740);
    or g1392(n816 ,n593 ,n766);
    nor g1393(n814 ,n599 ,n765);
    nor g1394(n813 ,n244 ,n755);
    or g1395(n812 ,n253 ,n762);
    or g1396(n811 ,n46[3] ,n764);
    or g1397(n810 ,n267 ,n764);
    or g1398(n809 ,n267 ,n728);
    or g1399(n808 ,n46[3] ,n728);
    or g1400(n807 ,n253 ,n763);
    nor g1401(n805 ,n254 ,n734);
    or g1402(n804 ,n252 ,n732);
    not g1403(n766 ,n765);
    not g1404(n762 ,n763);
    not g1405(n760 ,n761);
    nor g1406(n759 ,n443 ,n696);
    nor g1407(n758 ,n519 ,n663);
    nor g1408(n757 ,n278 ,n659);
    or g1409(n756 ,n340 ,n668);
    or g1410(n755 ,n254 ,n674);
    or g1411(n754 ,n275 ,n667);
    nor g1412(n753 ,n480 ,n696);
    nor g1413(n752 ,n306 ,n696);
    nor g1414(n751 ,n281 ,n696);
    nor g1415(n750 ,n309 ,n658);
    nor g1416(n749 ,n564 ,n696);
    nor g1417(n748 ,n327 ,n658);
    nor g1418(n747 ,n476 ,n696);
    nor g1419(n746 ,n459 ,n696);
    nor g1420(n745 ,n263 ,n702);
    nor g1421(n744 ,n533 ,n658);
    nor g1422(n743 ,n489 ,n658);
    nor g1423(n742 ,n310 ,n658);
    nor g1424(n741 ,n288 ,n658);
    nor g1425(n740 ,n301 ,n658);
    nor g1426(n739 ,n292 ,n696);
    nor g1427(n738 ,n343 ,n658);
    nor g1428(n737 ,n269 ,n659);
    nor g1429(n736 ,n267 ,n659);
    nor g1430(n735 ,n270 ,n659);
    nor g1431(n765 ,n638 ,n672);
    or g1432(n764 ,n278 ,n666);
    nor g1433(n763 ,n1879 ,n661);
    nor g1434(n761 ,n263 ,n698);
    not g1435(n733 ,n732);
    not g1436(n731 ,n730);
    not g1437(n725 ,n726);
    nor g1438(n724 ,n251 ,n645);
    nor g1439(n723 ,n600 ,n665);
    nor g1440(n722 ,n605 ,n700);
    nor g1441(n721 ,n413 ,n694);
    nor g1442(n720 ,n263 ,n697);
    nor g1443(n719 ,n692 ,n688);
    nor g1444(n718 ,n25[0] ,n648);
    nor g1445(n717 ,n638 ,n671);
    or g1446(n716 ,n21[4] ,n667);
    nor g1447(n715 ,n48[2] ,n647);
    nor g1448(n714 ,n642 ,n682);
    or g1449(n712 ,n44[4] ,n668);
    nor g1450(n711 ,n250 ,n657);
    nor g1451(n710 ,n639 ,n665);
    nor g1452(n709 ,n693 ,n683);
    nor g1453(n708 ,n246 ,n651);
    nor g1454(n707 ,n246 ,n653);
    nor g1455(n706 ,n251 ,n643);
    nor g1456(n705 ,n695 ,n690);
    nor g1457(n704 ,n649 ,n685);
    nor g1458(n703 ,n25[0] ,n701);
    or g1459(n734 ,n252 ,n243);
    nor g1460(n732 ,n654 ,n656);
    nor g1461(n730 ,n247 ,n655);
    nor g1462(n729 ,n244 ,n673);
    or g1463(n728 ,n46[0] ,n666);
    nor g1464(n726 ,n662 ,n660);
    not g1465(n702 ,n701);
    not g1466(n700 ,n699);
    not g1467(n698 ,n697);
    nor g1468(n695 ,n498 ,n636);
    nor g1469(n694 ,n277 ,n600);
    nor g1470(n693 ,n565 ,n636);
    nor g1471(n692 ,n457 ,n636);
    nor g1472(n691 ,n323 ,n586);
    nor g1473(n690 ,n397 ,n635);
    nor g1474(n689 ,n342 ,n586);
    nor g1475(n688 ,n357 ,n635);
    nor g1476(n687 ,n495 ,n586);
    nor g1477(n686 ,n344 ,n586);
    nor g1478(n685 ,n396 ,n635);
    nor g1479(n684 ,n484 ,n586);
    nor g1480(n683 ,n394 ,n635);
    nor g1481(n682 ,n392 ,n635);
    nor g1482(n681 ,n296 ,n586);
    nor g1483(n680 ,n454 ,n586);
    nor g1484(n679 ,n513 ,n586);
    nor g1485(n678 ,n510 ,n586);
    nor g1486(n677 ,n473 ,n586);
    nor g1487(n676 ,n280 ,n586);
    nor g1488(n675 ,n271 ,n586);
    nor g1489(n701 ,n432 ,n631);
    nor g1490(n699 ,n274 ,n630);
    nor g1491(n697 ,n272 ,n601);
    or g1492(n696 ,n271 ,n604);
    not g1493(n674 ,n673);
    not g1494(n672 ,n671);
    not g1495(n670 ,n669);
    not g1496(n665 ,n664);
    not g1497(n663 ,n662);
    not g1498(n661 ,n660);
    nor g1499(n657 ,n625 ,n610);
    nor g1500(n656 ,n639 ,n593);
    nor g1501(n655 ,n629 ,n633);
    nor g1502(n654 ,n265 ,n592);
    nor g1503(n653 ,n622 ,n616);
    nor g1504(n652 ,n1916 ,n573);
    nor g1505(n651 ,n623 ,n628);
    or g1506(n650 ,n48[2] ,n607);
    nor g1507(n649 ,n485 ,n636);
    nor g1508(n648 ,n637 ,n599);
    nor g1509(n647 ,n602 ,n606);
    or g1510(n646 ,n25[1] ,n640);
    nor g1511(n645 ,n624 ,n584);
    or g1512(n644 ,n252 ,n587);
    nor g1513(n643 ,n626 ,n611);
    nor g1514(n642 ,n494 ,n636);
    nor g1515(n673 ,n27[1] ,n583);
    nor g1516(n671 ,n18[1] ,n578);
    nor g1517(n669 ,n25[1] ,n601);
    or g1518(n668 ,n581 ,n580);
    or g1519(n667 ,n579 ,n582);
    or g1520(n666 ,n253 ,n635);
    nor g1521(n664 ,n25[1] ,n641);
    nor g1522(n662 ,n412 ,n587);
    nor g1523(n660 ,n48[2] ,n588);
    or g1524(n659 ,n253 ,n636);
    or g1525(n658 ,n22[3] ,n604);
    not g1526(n641 ,n640);
    not g1527(n638 ,n637);
    not g1528(n635 ,n636);
    nor g1529(n634 ,n436 ,n252);
    or g1530(n633 ,n429 ,n426);
    or g1531(n632 ,n377 ,n1936);
    or g1532(n631 ,n268 ,n431);
    or g1533(n630 ,n416 ,n273);
    or g1534(n629 ,n419 ,n423);
    nor g1535(n628 ,n515 ,n1943);
    or g1536(n627 ,n362 ,n1936);
    nor g1537(n626 ,n264 ,n403);
    nor g1538(n625 ,n264 ,n409);
    nor g1539(n624 ,n264 ,n389);
    nor g1540(n623 ,n264 ,n370);
    nor g1541(n622 ,n264 ,n387);
    nor g1542(n621 ,n439 ,n252);
    nor g1543(n620 ,n440 ,n252);
    nor g1544(n619 ,n434 ,n252);
    nor g1545(n618 ,n435 ,n252);
    or g1546(n617 ,n361 ,n1936);
    nor g1547(n616 ,n491 ,n1943);
    or g1548(n615 ,n402 ,n1936);
    or g1549(n614 ,n406 ,n1936);
    or g1550(n613 ,n368 ,n1936);
    or g1551(n612 ,n390 ,n1936);
    nor g1552(n611 ,n460 ,n1943);
    nor g1553(n610 ,n291 ,n1943);
    or g1554(n609 ,n365 ,n1936);
    or g1555(n608 ,n411 ,n1936);
    nor g1556(n640 ,n413 ,n277);
    or g1557(n639 ,n276 ,n25[2]);
    nor g1558(n637 ,n265 ,n272);
    nor g1559(n636 ,n1877 ,n1878);
    not g1560(n607 ,n606);
    not g1561(n603 ,n602);
    not g1562(n600 ,n599);
    not g1563(n593 ,n592);
    not g1564(n588 ,n587);
    or g1565(n585 ,n252 ,n23[3]);
    nor g1566(n584 ,n314 ,n1943);
    or g1567(n583 ,n27[0] ,n27[2]);
    or g1568(n582 ,n21[3] ,n21[2]);
    or g1569(n581 ,n44[1] ,n44[0]);
    or g1570(n580 ,n44[3] ,n44[2]);
    or g1571(n579 ,n21[1] ,n21[0]);
    or g1572(n578 ,n18[0] ,n18[2]);
    or g1573(n577 ,n26[0] ,n1936);
    or g1574(n576 ,n23[1] ,n23[2]);
    or g1575(n575 ,n252 ,n1925);
    or g1576(n574 ,n376 ,n1936);
    or g1577(n573 ,n413 ,n25[2]);
    or g1578(n572 ,n253 ,n254);
    nor g1579(n571 ,n263 ,n1944);
    or g1580(n570 ,n263 ,n25[2]);
    nor g1581(n606 ,n417 ,n48[1]);
    or g1582(n605 ,n418 ,n48[2]);
    or g1583(n604 ,n253 ,n264);
    nor g1584(n602 ,n418 ,n48[0]);
    or g1585(n601 ,n25[0] ,n25[2]);
    nor g1586(n599 ,n25[2] ,n2);
    or g1587(n598 ,n270 ,n269);
    or g1588(n597 ,n266 ,n45[3]);
    or g1589(n596 ,n414 ,n45[0]);
    or g1590(n595 ,n269 ,n46[2]);
    or g1591(n594 ,n46[2] ,n46[1]);
    nor g1592(n592 ,n25[0] ,n25[1]);
    or g1593(n591 ,n270 ,n46[1]);
    or g1594(n590 ,n266 ,n414);
    or g1595(n589 ,n45[0] ,n45[3]);
    nor g1596(n587 ,n48[0] ,n48[1]);
    or g1597(n586 ,n253 ,n1943);
    not g1598(n569 ,n36[5]);
    not g1599(n568 ,n47[5]);
    not g1600(n567 ,n28[0]);
    not g1601(n566 ,n41[2]);
    not g1602(n565 ,n44[1]);
    not g1603(n564 ,n20[0]);
    not g1604(n563 ,n43[5]);
    not g1605(n562 ,n40[4]);
    not g1606(n561 ,n33[1]);
    not g1607(n560 ,n36[4]);
    not g1608(n559 ,n35[1]);
    not g1609(n558 ,n47[1]);
    not g1610(n557 ,n28[4]);
    not g1611(n556 ,n29[1]);
    not g1612(n555 ,n28[1]);
    not g1613(n554 ,n31[2]);
    not g1614(n553 ,n44[4]);
    not g1615(n552 ,n36[7]);
    not g1616(n551 ,n26[2]);
    not g1617(n550 ,n29[6]);
    not g1618(n549 ,n29[7]);
    not g1619(n548 ,n37[1]);
    not g1620(n547 ,n33[2]);
    not g1621(n546 ,n26[7]);
    not g1622(n545 ,n30[5]);
    not g1623(n544 ,n43[3]);
    not g1624(n543 ,n33[4]);
    not g1625(n542 ,n17[4]);
    not g1626(n541 ,n37[2]);
    not g1627(n540 ,n43[0]);
    not g1628(n539 ,n47[6]);
    not g1629(n538 ,n31[5]);
    not g1630(n537 ,n33[6]);
    not g1631(n536 ,n21[0]);
    not g1632(n535 ,n17[9]);
    not g1633(n534 ,n43[1]);
    not g1634(n533 ,n19[7]);
    not g1635(n532 ,n32[4]);
    not g1636(n531 ,n43[2]);
    not g1637(n530 ,n17[2]);
    not g1638(n529 ,n33[5]);
    not g1639(n528 ,n40[7]);
    not g1640(n527 ,n41[1]);
    not g1641(n526 ,n34[1]);
    not g1642(n525 ,n32[0]);
    not g1643(n524 ,n35[5]);
    not g1644(n523 ,n35[3]);
    not g1645(n522 ,n32[2]);
    not g1646(n521 ,n38[6]);
    not g1647(n520 ,n35[7]);
    not g1648(n519 ,n6);
    not g1649(n518 ,n44[0]);
    not g1650(n517 ,n44[1]);
    not g1651(n516 ,n29[3]);
    not g1652(n515 ,n21[0]);
    not g1653(n514 ,n36[1]);
    not g1654(n513 ,n12[1]);
    not g1655(n512 ,n38[2]);
    not g1656(n511 ,n40[1]);
    not g1657(n510 ,n12[3]);
    not g1658(n509 ,n37[7]);
    not g1659(n508 ,n47[2]);
    not g1660(n507 ,n39[3]);
    not g1661(n506 ,n47[4]);
    not g1662(n505 ,n36[6]);
    not g1663(n504 ,n47[7]);
    not g1664(n503 ,n39[4]);
    not g1665(n502 ,n40[0]);
    not g1666(n501 ,n43[4]);
    not g1667(n500 ,n31[0]);
    not g1668(n499 ,n43[7]);
    not g1669(n498 ,n44[3]);
    not g1670(n497 ,n35[4]);
    not g1671(n496 ,n42[3]);
    not g1672(n495 ,n12[0]);
    not g1673(n494 ,n44[0]);
    not g1674(n493 ,n30[0]);
    not g1675(n492 ,n41[0]);
    not g1676(n491 ,n21[1]);
    not g1677(n490 ,n32[7]);
    not g1678(n489 ,n19[3]);
    not g1679(n488 ,n28[3]);
    not g1680(n487 ,n42[7]);
    not g1681(n486 ,n31[7]);
    not g1682(n485 ,n44[2]);
    not g1683(n484 ,n12[5]);
    not g1684(n483 ,n38[3]);
    not g1685(n482 ,n26[10]);
    not g1686(n481 ,n33[3]);
    not g1687(n480 ,n20[2]);
    not g1688(n479 ,n44[3]);
    not g1689(n478 ,n39[6]);
    not g1690(n477 ,n31[4]);
    not g1691(n476 ,n20[6]);
    not g1692(n475 ,n26[1]);
    not g1693(n474 ,n38[0]);
    not g1694(n473 ,n12[2]);
    not g1695(n472 ,n35[0]);
    not g1696(n471 ,n17[3]);
    not g1697(n470 ,n30[3]);
    not g1698(n469 ,n34[3]);
    not g1699(n468 ,n39[1]);
    not g1700(n467 ,n47[0]);
    not g1701(n466 ,n26[3]);
    not g1702(n465 ,n41[3]);
    not g1703(n464 ,n42[0]);
    not g1704(n463 ,n34[0]);
    not g1705(n462 ,n17[6]);
    not g1706(n461 ,n26[4]);
    not g1707(n460 ,n21[3]);
    not g1708(n459 ,n20[4]);
    not g1709(n458 ,n32[1]);
    not g1710(n457 ,n44[4]);
    not g1711(n456 ,n28[7]);
    not g1712(n455 ,n42[6]);
    not g1713(n454 ,n12[4]);
    not g1714(n453 ,n37[5]);
    not g1715(n452 ,n28[6]);
    not g1716(n451 ,n41[6]);
    not g1717(n450 ,n37[0]);
    not g1718(n449 ,n34[4]);
    not g1719(n448 ,n34[5]);
    not g1720(n447 ,n34[2]);
    not g1721(n446 ,n21[3]);
    not g1722(n445 ,n29[2]);
    not g1723(n444 ,n43[6]);
    not g1724(n443 ,n20[7]);
    not g1725(n442 ,n40[3]);
    not g1726(n441 ,n26[5]);
    not g1727(n440 ,n10);
    not g1728(n439 ,n8);
    not g1729(n438 ,n26[0]);
    not g1730(n437 ,n24[0]);
    not g1731(n436 ,n11);
    not g1732(n435 ,n14[1]);
    not g1733(n434 ,n9);
    not g1734(n433 ,n17[0]);
    not g1735(n432 ,n18[1]);
    not g1736(n431 ,n18[2]);
    not g1737(n430 ,n24[7]);
    not g1738(n429 ,n23[2]);
    not g1739(n428 ,n24[3]);
    not g1740(n427 ,n24[4]);
    not g1741(n426 ,n23[3]);
    not g1742(n425 ,n45[2]);
    not g1743(n424 ,n24[1]);
    not g1744(n423 ,n23[1]);
    not g1745(n422 ,n24[2]);
    not g1746(n421 ,n24[5]);
    not g1747(n420 ,n24[6]);
    not g1748(n419 ,n23[0]);
    not g1749(n418 ,n48[1]);
    not g1750(n417 ,n48[0]);
    not g1751(n416 ,n27[0]);
    not g1752(n415 ,n45[1]);
    not g1753(n414 ,n45[3]);
    not g1754(n413 ,n25[0]);
    not g1755(n412 ,n48[2]);
    not g1756(n411 ,n1908);
    not g1757(n410 ,n1883);
    not g1758(n409 ,n1938);
    not g1759(n408 ,n1931);
    not g1760(n407 ,n1896);
    not g1761(n406 ,n1902);
    not g1762(n405 ,n1888);
    not g1763(n404 ,n1885);
    not g1764(n403 ,n1939);
    not g1765(n402 ,n1904);
    not g1766(n401 ,n1932);
    not g1767(n400 ,n1895);
    not g1768(n399 ,n1920);
    not g1769(n398 ,n1935);
    not g1770(n397 ,n1927);
    not g1771(n396 ,n1928);
    not g1772(n395 ,n1924);
    not g1773(n394 ,n1929);
    not g1774(n393 ,n1894);
    not g1775(n392 ,n1930);
    not g1776(n391 ,n1897);
    not g1777(n390 ,n1910);
    not g1778(n389 ,n1940);
    not g1779(n388 ,n1933);
    not g1780(n387 ,n1941);
    not g1781(n386 ,n1900);
    not g1782(n385 ,n1915);
    not g1783(n384 ,n1899);
    not g1784(n383 ,n1886);
    not g1785(n382 ,n1884);
    not g1786(n381 ,n1891);
    not g1787(n380 ,n1921);
    not g1788(n379 ,n1887);
    not g1789(n378 ,n1889);
    not g1790(n377 ,n1906);
    not g1791(n376 ,n1911);
    not g1792(n375 ,n1918);
    not g1793(n374 ,n1934);
    not g1794(n373 ,n1893);
    not g1795(n372 ,n1922);
    not g1796(n371 ,n1890);
    not g1797(n370 ,n1942);
    not g1798(n369 ,n1898);
    not g1799(n368 ,n1905);
    not g1800(n367 ,n1882);
    not g1801(n366 ,n1913);
    not g1802(n365 ,n1909);
    not g1803(n364 ,n1881);
    not g1804(n363 ,n1901);
    not g1805(n362 ,n1903);
    not g1806(n361 ,n1907);
    not g1807(n360 ,n1914);
    not g1808(n359 ,n1912);
    not g1809(n358 ,n1880);
    not g1810(n357 ,n1926);
    not g1811(n356 ,n1923);
    not g1812(n355 ,n1892);
    not g1813(n354 ,n1917);
    not g1814(n353 ,n29[0]);
    not g1815(n352 ,n40[6]);
    not g1816(n351 ,n28[2]);
    not g1817(n350 ,n38[4]);
    not g1818(n349 ,n35[6]);
    not g1819(n348 ,n39[7]);
    not g1820(n347 ,n30[6]);
    not g1821(n346 ,n33[0]);
    not g1822(n345 ,n42[4]);
    not g1823(n344 ,n22[0]);
    not g1824(n343 ,n19[5]);
    not g1825(n342 ,n22[2]);
    not g1826(n341 ,n21[1]);
    not g1827(n340 ,n44[4]);
    not g1828(n339 ,n41[5]);
    not g1829(n338 ,n47[3]);
    not g1830(n337 ,n31[3]);
    not g1831(n336 ,n33[7]);
    not g1832(n335 ,n40[2]);
    not g1833(n334 ,n35[2]);
    not g1834(n333 ,n41[4]);
    not g1835(n332 ,n30[4]);
    not g1836(n331 ,n41[7]);
    not g1837(n330 ,n32[3]);
    not g1838(n329 ,n17[7]);
    not g1839(n328 ,n42[2]);
    not g1840(n327 ,n19[0]);
    not g1841(n326 ,n29[5]);
    not g1842(n325 ,n21[2]);
    not g1843(n324 ,n37[6]);
    not g1844(n323 ,n22[1]);
    not g1845(n322 ,n34[6]);
    not g1846(n321 ,n40[5]);
    not g1847(n320 ,n36[0]);
    not g1848(n319 ,n31[1]);
    not g1849(n318 ,n38[7]);
    not g1850(n317 ,n42[1]);
    not g1851(n316 ,n32[5]);
    not g1852(n315 ,n36[2]);
    not g1853(n314 ,n21[2]);
    not g1854(n313 ,n30[2]);
    not g1855(n312 ,n36[3]);
    not g1856(n311 ,n39[0]);
    not g1857(n310 ,n19[4]);
    not g1858(n309 ,n19[1]);
    not g1859(n308 ,n30[7]);
    not g1860(n307 ,n32[6]);
    not g1861(n306 ,n20[3]);
    not g1862(n305 ,n26[9]);
    not g1863(n304 ,n38[5]);
    not g1864(n303 ,n17[10]);
    not g1865(n302 ,n37[4]);
    not g1866(n301 ,n19[2]);
    not g1867(n300 ,n44[2]);
    not g1868(n299 ,n26[6]);
    not g1869(n298 ,n17[5]);
    not g1870(n297 ,n17[8]);
    not g1871(n296 ,n12[7]);
    not g1872(n295 ,n30[1]);
    not g1873(n294 ,n26[8]);
    not g1874(n293 ,n29[4]);
    not g1875(n292 ,n20[1]);
    not g1876(n291 ,n21[4]);
    not g1877(n290 ,n17[1]);
    not g1878(n289 ,n34[7]);
    not g1879(n288 ,n19[6]);
    not g1880(n287 ,n39[2]);
    not g1881(n286 ,n42[5]);
    not g1882(n285 ,n38[1]);
    not g1883(n284 ,n28[5]);
    not g1884(n283 ,n39[5]);
    not g1885(n282 ,n37[3]);
    not g1886(n281 ,n20[5]);
    not g1887(n280 ,n12[6]);
    not g1888(n279 ,n31[6]);
    not g1889(n278 ,n46[0]);
    not g1890(n277 ,n1916);
    not g1891(n276 ,n2);
    not g1892(n275 ,n21[4]);
    not g1893(n274 ,n27[1]);
    not g1894(n273 ,n27[2]);
    not g1895(n272 ,n1944);
    not g1896(n271 ,n22[3]);
    not g1897(n270 ,n46[2]);
    not g1898(n269 ,n46[1]);
    not g1899(n268 ,n18[0]);
    not g1900(n267 ,n46[3]);
    not g1901(n266 ,n45[0]);
    not g1902(n265 ,n25[2]);
    not g1903(n264 ,n1943);
    not g1904(n263 ,n25[1]);
    not g1905(n262 ,n5[4]);
    not g1906(n261 ,n5[1]);
    not g1907(n260 ,n5[2]);
    not g1908(n259 ,n5[7]);
    not g1909(n258 ,n5[6]);
    not g1910(n257 ,n5[3]);
    not g1911(n256 ,n5[0]);
    not g1912(n255 ,n5[5]);
    not g1913(n254 ,n1936);
    not g1914(n253 ,n1);
    not g1915(n252 ,n1);
    not g1916(n251 ,n1);
    not g1917(n250 ,n1);
    not g1918(n249 ,n1);
    not g1919(n248 ,n1);
    not g1920(n247 ,n1);
    not g1921(n246 ,n1);
    not g1922(n245 ,n1);
    or g1923(n244 ,n412 ,n588);
    or g1924(n243 ,n48[2] ,n603);
    xor g1925(n1931 ,n44[4] ,n53);
    xor g1926(n1932 ,n44[3] ,n51);
    nor g1927(n53 ,n44[3] ,n52);
    xor g1928(n1933 ,n44[2] ,n49);
    not g1929(n52 ,n51);
    nor g1930(n51 ,n44[2] ,n50);
    xnor g1931(n1934 ,n44[1] ,n44[0]);
    not g1932(n50 ,n49);
    nor g1933(n49 ,n44[1] ,n44[0]);
    not g1934(n1935 ,n44[0]);
    xor g1935(n1938 ,n21[4] ,n58);
    xor g1936(n1939 ,n21[3] ,n56);
    nor g1937(n58 ,n21[3] ,n57);
    xor g1938(n1940 ,n21[2] ,n54);
    not g1939(n57 ,n56);
    nor g1940(n56 ,n21[2] ,n55);
    xnor g1941(n1941 ,n21[1] ,n21[0]);
    not g1942(n55 ,n54);
    nor g1943(n54 ,n21[1] ,n21[0]);
    not g1944(n1942 ,n21[0]);
    or g1945(n1937 ,n60 ,n61);
    or g1946(n61 ,n44[3] ,n59);
    or g1947(n60 ,n44[2] ,n44[0]);
    or g1948(n59 ,n44[4] ,n44[1]);
    or g1949(n1943 ,n63 ,n64);
    or g1950(n64 ,n21[3] ,n62);
    or g1951(n63 ,n21[2] ,n21[0]);
    or g1952(n62 ,n21[4] ,n21[1]);
    or g1953(n1936 ,n26[10] ,n79);
    nor g1954(n79 ,n73 ,n78);
    nor g1955(n78 ,n26[7] ,n77);
    nor g1956(n77 ,n67 ,n76);
    or g1957(n76 ,n69 ,n75);
    nor g1958(n75 ,n71 ,n74);
    or g1959(n74 ,n26[2] ,n72);
    or g1960(n73 ,n70 ,n68);
    nor g1961(n72 ,n65 ,n66);
    or g1962(n71 ,n26[4] ,n26[3]);
    not g1963(n70 ,n26[9]);
    not g1964(n69 ,n26[6]);
    not g1965(n68 ,n26[8]);
    not g1966(n67 ,n26[5]);
    not g1967(n66 ,n26[0]);
    not g1968(n65 ,n26[1]);
    or g1969(n1916 ,n84 ,n92);
    nor g1970(n92 ,n83 ,n91);
    or g1971(n91 ,n81 ,n90);
    nor g1972(n90 ,n17[6] ,n89);
    nor g1973(n89 ,n87 ,n88);
    nor g1974(n88 ,n86 ,n85);
    or g1975(n87 ,n82 ,n80);
    or g1976(n86 ,n17[3] ,n17[2]);
    or g1977(n85 ,n17[1] ,n17[0]);
    or g1978(n84 ,n17[10] ,n17[9]);
    not g1979(n83 ,n17[7]);
    not g1980(n82 ,n17[5]);
    not g1981(n81 ,n17[8]);
    not g1982(n80 ,n17[4]);
    or g1983(n1944 ,n17[10] ,n107);
    nor g1984(n107 ,n101 ,n106);
    nor g1985(n106 ,n17[7] ,n105);
    nor g1986(n105 ,n95 ,n104);
    or g1987(n104 ,n97 ,n103);
    nor g1988(n103 ,n99 ,n102);
    or g1989(n102 ,n17[2] ,n100);
    or g1990(n101 ,n98 ,n96);
    nor g1991(n100 ,n93 ,n94);
    or g1992(n99 ,n17[4] ,n17[3]);
    not g1993(n98 ,n17[9]);
    not g1994(n97 ,n17[6]);
    not g1995(n96 ,n17[8]);
    not g1996(n95 ,n17[5]);
    not g1997(n94 ,n17[0]);
    not g1998(n93 ,n17[1]);
    xor g1999(n1882 ,n45[3] ,n115);
    nor g2000(n1881 ,n114 ,n115);
    nor g2001(n115 ,n110 ,n113);
    nor g2002(n114 ,n45[2] ,n112);
    nor g2003(n1880 ,n112 ,n111);
    not g2004(n113 ,n112);
    nor g2005(n112 ,n108 ,n109);
    nor g2006(n111 ,n45[1] ,n45[0]);
    not g2007(n110 ,n45[2]);
    not g2008(n109 ,n45[0]);
    not g2009(n108 ,n45[1]);
    nor g2010(n1910 ,n150 ,n151);
    nor g2011(n151 ,n116 ,n149);
    nor g2012(n150 ,n26[9] ,n148);
    nor g2013(n1909 ,n147 ,n148);
    not g2014(n149 ,n148);
    nor g2015(n148 ,n118 ,n146);
    nor g2016(n147 ,n26[8] ,n145);
    nor g2017(n1908 ,n144 ,n145);
    not g2018(n146 ,n145);
    nor g2019(n145 ,n124 ,n143);
    nor g2020(n144 ,n26[7] ,n142);
    nor g2021(n1907 ,n141 ,n142);
    not g2022(n143 ,n142);
    nor g2023(n142 ,n119 ,n140);
    nor g2024(n141 ,n26[6] ,n139);
    nor g2025(n1906 ,n138 ,n139);
    not g2026(n140 ,n139);
    nor g2027(n139 ,n120 ,n137);
    nor g2028(n138 ,n26[5] ,n136);
    nor g2029(n1905 ,n135 ,n136);
    not g2030(n137 ,n136);
    nor g2031(n136 ,n117 ,n134);
    nor g2032(n135 ,n26[4] ,n133);
    nor g2033(n1904 ,n132 ,n133);
    not g2034(n134 ,n133);
    nor g2035(n133 ,n123 ,n131);
    nor g2036(n132 ,n26[3] ,n130);
    nor g2037(n1903 ,n129 ,n130);
    not g2038(n131 ,n130);
    nor g2039(n130 ,n121 ,n128);
    nor g2040(n129 ,n26[2] ,n127);
    nor g2041(n1902 ,n127 ,n126);
    not g2042(n128 ,n127);
    nor g2043(n127 ,n122 ,n125);
    nor g2044(n126 ,n26[1] ,n26[0]);
    not g2045(n125 ,n26[0]);
    not g2046(n124 ,n26[7]);
    not g2047(n123 ,n26[3]);
    not g2048(n122 ,n26[1]);
    not g2049(n121 ,n26[2]);
    not g2050(n120 ,n26[5]);
    not g2051(n119 ,n26[6]);
    not g2052(n118 ,n26[8]);
    not g2053(n117 ,n26[4]);
    not g2054(n116 ,n26[9]);
    xor g2055(n1918 ,n27[2] ,n155);
    nor g2056(n1917 ,n155 ,n154);
    nor g2057(n155 ,n153 ,n152);
    nor g2058(n154 ,n27[1] ,n27[0]);
    not g2059(n153 ,n27[1]);
    not g2060(n152 ,n27[0]);
    xor g2061(n1899 ,n17[10] ,n191);
    nor g2062(n1898 ,n190 ,n191);
    nor g2063(n191 ,n156 ,n189);
    nor g2064(n190 ,n17[9] ,n188);
    nor g2065(n1897 ,n187 ,n188);
    not g2066(n189 ,n188);
    nor g2067(n188 ,n158 ,n186);
    nor g2068(n187 ,n17[8] ,n185);
    nor g2069(n1896 ,n184 ,n185);
    not g2070(n186 ,n185);
    nor g2071(n185 ,n164 ,n183);
    nor g2072(n184 ,n17[7] ,n182);
    nor g2073(n1895 ,n181 ,n182);
    not g2074(n183 ,n182);
    nor g2075(n182 ,n159 ,n180);
    nor g2076(n181 ,n17[6] ,n179);
    nor g2077(n1894 ,n178 ,n179);
    not g2078(n180 ,n179);
    nor g2079(n179 ,n160 ,n177);
    nor g2080(n178 ,n17[5] ,n176);
    nor g2081(n1915 ,n175 ,n176);
    not g2082(n177 ,n176);
    nor g2083(n176 ,n157 ,n174);
    nor g2084(n175 ,n17[4] ,n173);
    nor g2085(n1914 ,n172 ,n173);
    not g2086(n174 ,n173);
    nor g2087(n173 ,n163 ,n171);
    nor g2088(n172 ,n17[3] ,n170);
    nor g2089(n1913 ,n169 ,n170);
    not g2090(n171 ,n170);
    nor g2091(n170 ,n161 ,n168);
    nor g2092(n169 ,n17[2] ,n167);
    nor g2093(n1912 ,n167 ,n166);
    not g2094(n168 ,n167);
    nor g2095(n167 ,n162 ,n165);
    nor g2096(n166 ,n17[1] ,n17[0]);
    not g2097(n165 ,n17[0]);
    not g2098(n164 ,n17[7]);
    not g2099(n163 ,n17[3]);
    not g2100(n162 ,n17[1]);
    not g2101(n161 ,n17[2]);
    not g2102(n160 ,n17[5]);
    not g2103(n159 ,n17[6]);
    not g2104(n158 ,n17[8]);
    not g2105(n157 ,n17[4]);
    not g2106(n156 ,n17[9]);
    xor g2107(n1901 ,n18[2] ,n195);
    nor g2108(n1900 ,n195 ,n194);
    nor g2109(n195 ,n193 ,n192);
    nor g2110(n194 ,n18[1] ,n18[0]);
    not g2111(n193 ,n18[1]);
    not g2112(n192 ,n18[0]);
    xor g2113(n1885 ,n23[3] ,n203);
    nor g2114(n1884 ,n202 ,n203);
    nor g2115(n203 ,n198 ,n201);
    nor g2116(n202 ,n23[2] ,n200);
    nor g2117(n1883 ,n200 ,n199);
    not g2118(n201 ,n200);
    nor g2119(n200 ,n196 ,n197);
    nor g2120(n199 ,n23[1] ,n23[0]);
    not g2121(n198 ,n23[2]);
    not g2122(n197 ,n23[0]);
    not g2123(n196 ,n23[1]);
    nor g2124(n1921 ,n213 ,n214);
    nor g2125(n214 ,n205 ,n212);
    nor g2126(n213 ,n21[3] ,n211);
    nor g2127(n1922 ,n210 ,n211);
    not g2128(n212 ,n211);
    nor g2129(n211 ,n206 ,n209);
    nor g2130(n210 ,n21[2] ,n208);
    nor g2131(n1923 ,n208 ,n207);
    not g2132(n209 ,n208);
    nor g2133(n208 ,n204 ,n1924);
    nor g2134(n207 ,n21[1] ,n21[0]);
    not g2135(n206 ,n21[2]);
    not g2136(n1924 ,n21[0]);
    not g2137(n205 ,n21[3]);
    not g2138(n204 ,n21[1]);
    xor g2139(n1889 ,n221 ,n46[3]);
    nor g2140(n1888 ,n220 ,n221);
    nor g2141(n221 ,n216 ,n219);
    nor g2142(n220 ,n46[2] ,n218);
    nor g2143(n1887 ,n218 ,n217);
    not g2144(n219 ,n218);
    nor g2145(n218 ,n215 ,n1886);
    nor g2146(n217 ,n46[1] ,n46[0]);
    not g2147(n216 ,n46[2]);
    not g2148(n1886 ,n46[0]);
    not g2149(n215 ,n46[1]);
    xor g2150(n1926 ,n44[4] ,n232);
    nor g2151(n1927 ,n231 ,n232);
    nor g2152(n232 ,n223 ,n230);
    nor g2153(n231 ,n44[3] ,n229);
    nor g2154(n1928 ,n228 ,n229);
    not g2155(n230 ,n229);
    nor g2156(n229 ,n224 ,n227);
    nor g2157(n228 ,n44[2] ,n226);
    nor g2158(n1929 ,n226 ,n225);
    not g2159(n227 ,n226);
    nor g2160(n226 ,n222 ,n1930);
    nor g2161(n225 ,n44[1] ,n44[0]);
    not g2162(n224 ,n44[2]);
    not g2163(n1930 ,n44[0]);
    not g2164(n223 ,n44[3]);
    not g2165(n222 ,n44[1]);
    xor g2166(n1893 ,n239 ,n22[3]);
    nor g2167(n1892 ,n238 ,n239);
    nor g2168(n239 ,n234 ,n237);
    nor g2169(n238 ,n22[2] ,n236);
    nor g2170(n1891 ,n236 ,n235);
    not g2171(n237 ,n236);
    nor g2172(n236 ,n233 ,n1890);
    nor g2173(n235 ,n22[1] ,n22[0]);
    not g2174(n234 ,n22[2]);
    not g2175(n1890 ,n22[0]);
    not g2176(n233 ,n22[1]);
    not g2177(n1919 ,n44[4]);
    nor g2178(n1925 ,n21[4] ,n242);
    nor g2179(n242 ,n240 ,n241);
    not g2180(n241 ,n21[2]);
    not g2181(n240 ,n21[3]);
    buf g2182(n1263 ,n21[4]);
    not g2183(n713 ,n243);
    buf g2184(n1132 ,n666);
    buf g2185(n727 ,n604);
    buf g2186(n1920 ,n214);
    buf g2187(n1911 ,n151);
endmodule
