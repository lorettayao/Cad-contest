module top(n0, n1, n4, n5, n2, n3, n6, n7, n12, n14, n15, n8, n9, n10, n11, n13);
    input n0, n1, n2, n3;
    input [7:0] n4, n5;
    output [2:0] n6, n7, n8, n9, n10, n11;
    output [7:0] n12, n13;
    output n14, n15;
    wire n0, n1, n2, n3;
    wire [7:0] n4, n5;
    wire [2:0] n6, n7, n8, n9, n10, n11;
    wire [7:0] n12, n13;
    wire n14, n15;
    wire [31:0] n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259;
    buf g0(n13[6], n8[0]);
    buf g1(n13[7], n8[1]);
    buf g2(n12[7], 1'b0);
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n249), .Q(n7[0]));
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n248), .Q(n7[1]));
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n247), .Q(n7[2]));
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n244), .Q(n6[1]));
    dff g7(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n246), .Q(n6[2]));
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n245), .Q(n6[0]));
    or g9(n249 ,n117 ,n245);
    or g10(n248 ,n115 ,n244);
    or g11(n247 ,n116 ,n246);
    nor g12(n246 ,n65 ,n242);
    nor g13(n245 ,n65 ,n241);
    nor g14(n244 ,n65 ,n243);
    nor g15(n243 ,n186 ,n238);
    nor g16(n242 ,n236 ,n240);
    nor g17(n241 ,n237 ,n239);
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n234), .Q(n15));
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n233), .Q(n14));
    nor g20(n240 ,n196 ,n59);
    nor g21(n239 ,n194 ,n59);
    or g22(n238 ,n167 ,n235);
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n224), .Q(n16[4]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n229), .Q(n16[1]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n230), .Q(n16[2]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n226), .Q(n16[3]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n219), .Q(n16[7]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n223), .Q(n16[5]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n222), .Q(n16[6]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n227), .Q(n16[0]));
    nor g31(n237 ,n92 ,n232);
    nor g32(n236 ,n90 ,n232);
    nor g33(n235 ,n91 ,n232);
    nor g34(n234 ,n65 ,n228);
    nor g35(n233 ,n65 ,n225);
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n221), .Q(n16[8]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n220), .Q(n16[9]));
    not g38(n231 ,n232);
    or g39(n230 ,n211 ,n210);
    or g40(n229 ,n213 ,n212);
    nor g41(n228 ,n192 ,n217);
    or g42(n227 ,n215 ,n193);
    or g43(n226 ,n209 ,n208);
    nor g44(n232 ,n195 ,n197);
    nor g45(n225 ,n205 ,n204);
    or g46(n224 ,n207 ,n198);
    or g47(n223 ,n218 ,n191);
    or g48(n222 ,n203 ,n214);
    or g49(n221 ,n201 ,n206);
    or g50(n220 ,n199 ,n216);
    or g51(n219 ,n202 ,n200);
    nor g52(n218 ,n78 ,n189);
    nor g53(n217 ,n94 ,n185);
    nor g54(n216 ,n84 ,n190);
    nor g55(n215 ,n93 ,n189);
    nor g56(n214 ,n88 ,n190);
    nor g57(n213 ,n101 ,n189);
    nor g58(n212 ,n87 ,n190);
    nor g59(n211 ,n111 ,n189);
    nor g60(n210 ,n83 ,n190);
    nor g61(n209 ,n110 ,n189);
    nor g62(n208 ,n89 ,n190);
    nor g63(n207 ,n102 ,n189);
    nor g64(n206 ,n86 ,n190);
    nor g65(n205 ,n95 ,n183);
    nor g66(n204 ,n154 ,n182);
    nor g67(n203 ,n109 ,n189);
    nor g68(n202 ,n70 ,n189);
    nor g69(n201 ,n99 ,n189);
    nor g70(n200 ,n85 ,n190);
    nor g71(n199 ,n79 ,n189);
    nor g72(n198 ,n81 ,n190);
    or g73(n197 ,n181 ,n180);
    or g74(n196 ,n139 ,n187);
    or g75(n195 ,n176 ,n179);
    or g76(n194 ,n139 ,n188);
    nor g77(n193 ,n16[0] ,n190);
    nor g78(n192 ,n3 ,n184);
    nor g79(n191 ,n82 ,n190);
    or g80(n188 ,n169 ,n170);
    or g81(n187 ,n171 ,n60);
    or g82(n186 ,n60 ,n168);
    or g83(n190 ,n259 ,n175);
    or g84(n189 ,n66 ,n175);
    not g85(n185 ,n184);
    not g86(n183 ,n182);
    or g87(n181 ,n147 ,n174);
    or g88(n180 ,n173 ,n172);
    or g89(n179 ,n149 ,n177);
    nor g90(n184 ,n3 ,n178);
    nor g91(n182 ,n154 ,n178);
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n159), .Q(n12[1]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n161), .Q(n12[2]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n151), .Q(n12[3]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n157), .Q(n12[5]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n158), .Q(n12[0]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n148), .Q(n12[4]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n152), .Q(n12[6]));
    nor g99(n177 ,n5[3] ,n153);
    nor g100(n176 ,n4[4] ,n150);
    nor g101(n178 ,n66 ,n154);
    nor g102(n174 ,n5[0] ,n146);
    nor g103(n173 ,n5[2] ,n145);
    nor g104(n172 ,n4[2] ,n156);
    or g105(n171 ,n143 ,n164);
    or g106(n170 ,n162 ,n155);
    or g107(n169 ,n167 ,n163);
    or g108(n168 ,n160 ,n164);
    or g109(n175 ,n65 ,n154);
    nor g110(n162 ,n68 ,n140);
    nor g111(n161 ,n65 ,n140);
    nor g112(n160 ,n76 ,n133);
    nor g113(n159 ,n65 ,n141);
    nor g114(n158 ,n65 ,n137);
    nor g115(n157 ,n65 ,n135);
    nor g116(n167 ,n67 ,n142);
    nor g117(n166 ,n75 ,n135);
    nor g118(n165 ,n69 ,n141);
    nor g119(n164 ,n72 ,n133);
    nor g120(n163 ,n80 ,n137);
    not g121(n156 ,n155);
    or g122(n153 ,n5[4] ,n135);
    nor g123(n152 ,n65 ,n138);
    nor g124(n151 ,n65 ,n133);
    or g125(n150 ,n4[5] ,n133);
    nor g126(n149 ,n5[5] ,n138);
    nor g127(n148 ,n65 ,n142);
    nor g128(n147 ,n4[0] ,n144);
    or g129(n146 ,n5[1] ,n137);
    or g130(n145 ,n4[3] ,n140);
    nor g131(n155 ,n4[1] ,n141);
    nor g132(n154 ,n134 ,n136);
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n131), .Q(n13[0]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n130), .Q(n13[1]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n129), .Q(n13[2]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n128), .Q(n13[3]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n127), .Q(n13[4]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n126), .Q(n13[5]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n114), .Q(n8[0]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n112), .Q(n8[2]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n123), .Q(n9[0]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n124), .Q(n9[1]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n125), .Q(n9[2]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n122), .Q(n10[0]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n118), .Q(n8[1]));
    not g146(n144 ,n143);
    not g147(n138 ,n139);
    not g148(n137 ,n136);
    not g149(n135 ,n134);
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n113), .Q(n11[0]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n132), .Q(n11[1]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n120), .Q(n11[2]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n121), .Q(n10[2]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n119), .Q(n10[1]));
    nor g155(n143 ,n6[2] ,n64);
    or g156(n142 ,n90 ,n61);
    or g157(n141 ,n6[2] ,n62);
    or g158(n140 ,n6[2] ,n63);
    nor g159(n139 ,n90 ,n63);
    nor g160(n136 ,n6[2] ,n61);
    nor g161(n134 ,n90 ,n62);
    or g162(n133 ,n90 ,n64);
    nor g163(n132 ,n100 ,n65);
    nor g164(n131 ,n65 ,n77);
    nor g165(n130 ,n65 ,n69);
    nor g166(n129 ,n65 ,n73);
    nor g167(n128 ,n65 ,n68);
    nor g168(n127 ,n95 ,n65);
    nor g169(n126 ,n94 ,n65);
    nor g170(n125 ,n96 ,n65);
    nor g171(n124 ,n74 ,n65);
    nor g172(n123 ,n103 ,n65);
    nor g173(n122 ,n107 ,n65);
    nor g174(n121 ,n104 ,n65);
    nor g175(n120 ,n71 ,n65);
    nor g176(n119 ,n98 ,n65);
    nor g177(n118 ,n91 ,n65);
    nor g178(n117 ,n105 ,n1);
    nor g179(n116 ,n108 ,n1);
    nor g180(n115 ,n97 ,n1);
    nor g181(n114 ,n92 ,n65);
    nor g182(n113 ,n106 ,n65);
    nor g183(n112 ,n90 ,n65);
    not g184(n111 ,n16[2]);
    not g185(n110 ,n16[3]);
    not g186(n109 ,n16[6]);
    not g187(n108 ,n7[2]);
    not g188(n107 ,n9[0]);
    not g189(n106 ,n10[0]);
    not g190(n105 ,n7[0]);
    not g191(n104 ,n9[2]);
    not g192(n103 ,n8[0]);
    not g193(n102 ,n16[4]);
    not g194(n101 ,n16[1]);
    not g195(n100 ,n10[1]);
    not g196(n99 ,n16[8]);
    not g197(n98 ,n9[1]);
    not g198(n97 ,n7[1]);
    not g199(n96 ,n8[2]);
    not g200(n95 ,n14);
    not g201(n94 ,n15);
    not g202(n93 ,n16[0]);
    not g203(n92 ,n6[0]);
    not g204(n91 ,n6[1]);
    not g205(n90 ,n6[2]);
    not g206(n89 ,n252);
    not g207(n88 ,n255);
    not g208(n87 ,n250);
    not g209(n86 ,n257);
    not g210(n85 ,n256);
    not g211(n84 ,n258);
    not g212(n83 ,n251);
    not g213(n82 ,n254);
    not g214(n81 ,n253);
    not g215(n80 ,n5[0]);
    not g216(n79 ,n16[9]);
    not g217(n78 ,n16[5]);
    not g218(n77 ,n4[0]);
    not g219(n76 ,n4[5]);
    not g220(n75 ,n5[3]);
    not g221(n74 ,n8[1]);
    not g222(n73 ,n4[2]);
    not g223(n72 ,n4[4]);
    not g224(n71 ,n10[2]);
    not g225(n70 ,n16[7]);
    not g226(n69 ,n4[1]);
    not g227(n68 ,n4[3]);
    not g228(n67 ,n3);
    not g229(n66 ,n259);
    not g230(n65 ,n1);
    or g231(n64 ,n6[0] ,n6[1]);
    or g232(n63 ,n92 ,n91);
    or g233(n62 ,n91 ,n6[0]);
    or g234(n61 ,n92 ,n6[1]);
    or g235(n60 ,n165 ,n163);
    or g236(n59 ,n166 ,n231);
    nor g237(n259 ,n23 ,n26);
    or g238(n26 ,n18 ,n25);
    or g239(n25 ,n24 ,n22);
    or g240(n24 ,n21 ,n17);
    or g241(n23 ,n19 ,n20);
    nor g242(n22 ,n16[4] ,n16[3]);
    not g243(n21 ,n16[9]);
    not g244(n20 ,n16[5]);
    not g245(n19 ,n16[6]);
    not g246(n18 ,n16[7]);
    not g247(n17 ,n16[8]);
    xor g248(n258 ,n16[9] ,n58);
    nor g249(n257 ,n57 ,n58);
    nor g250(n58 ,n33 ,n56);
    nor g251(n57 ,n16[8] ,n55);
    nor g252(n256 ,n54 ,n55);
    not g253(n56 ,n55);
    nor g254(n55 ,n29 ,n53);
    nor g255(n54 ,n16[7] ,n52);
    nor g256(n255 ,n51 ,n52);
    not g257(n53 ,n52);
    nor g258(n52 ,n30 ,n50);
    nor g259(n51 ,n16[6] ,n49);
    nor g260(n254 ,n48 ,n49);
    not g261(n50 ,n49);
    nor g262(n49 ,n27 ,n47);
    nor g263(n48 ,n16[5] ,n46);
    nor g264(n253 ,n45 ,n46);
    not g265(n47 ,n46);
    nor g266(n46 ,n34 ,n44);
    nor g267(n45 ,n16[4] ,n43);
    nor g268(n252 ,n42 ,n43);
    not g269(n44 ,n43);
    nor g270(n43 ,n35 ,n41);
    nor g271(n42 ,n16[3] ,n40);
    nor g272(n251 ,n39 ,n40);
    not g273(n41 ,n40);
    nor g274(n40 ,n28 ,n38);
    nor g275(n39 ,n16[2] ,n37);
    nor g276(n250 ,n37 ,n36);
    not g277(n38 ,n37);
    nor g278(n37 ,n31 ,n32);
    nor g279(n36 ,n16[1] ,n16[0]);
    not g280(n35 ,n16[3]);
    not g281(n34 ,n16[4]);
    not g282(n33 ,n16[8]);
    not g283(n32 ,n16[0]);
    not g284(n31 ,n16[1]);
    not g285(n30 ,n16[6]);
    not g286(n29 ,n16[7]);
    not g287(n28 ,n16[2]);
    not g288(n27 ,n16[5]);
endmodule
