module top(n0, n1, n2, n3, n5, n8, n6, n9, n4, n7, n10, n11, n12, n13);
    input n0, n1;
    input [15:0] n2;
    input [7:0] n3, n4;
    input [3:0] n5, n6, n7;
    input [5:0] n8;
    input [1:0] n9;
    output [7:0] n10;
    output [3:0] n11;
    output [1:0] n12;
    output n13;
    wire n0, n1;
    wire [15:0] n2;
    wire [7:0] n3, n4;
    wire [3:0] n5, n6, n7;
    wire [5:0] n8;
    wire [1:0] n9;
    wire [7:0] n10;
    wire [3:0] n11;
    wire [1:0] n12;
    wire n13;
    wire [7:0] n14;
    wire [7:0] n15;
    wire [15:0] n16;
    wire [7:0] n17;
    wire [7:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [15:0] n22;
    wire [15:0] n23;
    wire [7:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [2:0] n37;
    wire [2:0] n38;
    wire [7:0] n39;
    wire [7:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [7:0] n43;
    wire [7:0] n44;
    wire [7:0] n45;
    wire [7:0] n46;
    wire [7:0] n47;
    wire n48, n49, n50, n51, n52, n53, n54, n55;
    wire n56, n57, n58, n59, n60, n61, n62, n63;
    wire n64, n65, n66, n67, n68, n69, n70, n71;
    wire n72, n73, n74, n75, n76, n77, n78, n79;
    wire n80, n81, n82, n83, n84, n85, n86, n87;
    wire n88, n89, n90, n91, n92, n93, n94, n95;
    wire n96, n97, n98, n99, n100, n101, n102, n103;
    wire n104, n105, n106, n107, n108, n109, n110, n111;
    wire n112, n113, n114, n115, n116, n117, n118, n119;
    wire n120, n121, n122, n123, n124, n125, n126, n127;
    wire n128, n129, n130, n131, n132, n133, n134, n135;
    wire n136, n137, n138, n139, n140, n141, n142, n143;
    wire n144, n145, n146, n147, n148, n149, n150, n151;
    wire n152, n153, n154, n155, n156, n157, n158, n159;
    wire n160, n161, n162, n163, n164, n165, n166, n167;
    wire n168, n169, n170, n171, n172, n173, n174, n175;
    wire n176, n177, n178, n179, n180, n181, n182, n183;
    wire n184, n185, n186, n187, n188, n189, n190, n191;
    wire n192, n193, n194, n195, n196, n197, n198, n199;
    wire n200, n201, n202, n203, n204, n205, n206, n207;
    wire n208, n209, n210, n211, n212, n213, n214, n215;
    wire n216, n217, n218, n219, n220, n221, n222, n223;
    wire n224, n225, n226, n227, n228, n229, n230, n231;
    wire n232, n233, n234, n235, n236, n237, n238, n239;
    wire n240, n241, n242, n243, n244, n245, n246, n247;
    wire n248, n249, n250, n251, n252, n253, n254, n255;
    wire n256, n257, n258, n259, n260, n261, n262, n263;
    wire n264, n265, n266, n267, n268, n269, n270, n271;
    wire n272, n273, n274, n275, n276, n277, n278, n279;
    wire n280, n281, n282, n283, n284, n285, n286, n287;
    wire n288, n289, n290, n291, n292, n293, n294, n295;
    wire n296, n297, n298, n299, n300, n301, n302, n303;
    wire n304, n305, n306, n307, n308, n309, n310, n311;
    wire n312, n313, n314, n315, n316, n317, n318, n319;
    wire n320, n321, n322, n323, n324, n325, n326, n327;
    wire n328, n329, n330, n331, n332, n333, n334, n335;
    wire n336, n337, n338, n339, n340, n341, n342, n343;
    wire n344, n345, n346, n347, n348, n349, n350, n351;
    wire n352, n353, n354, n355, n356, n357, n358, n359;
    wire n360, n361, n362, n363, n364, n365, n366, n367;
    wire n368, n369, n370, n371, n372, n373, n374, n375;
    wire n376, n377, n378, n379, n380, n381, n382, n383;
    wire n384, n385, n386, n387, n388, n389, n390, n391;
    wire n392, n393, n394, n395, n396, n397, n398, n399;
    wire n400, n401, n402, n403, n404, n405, n406, n407;
    wire n408, n409, n410, n411, n412, n413, n414, n415;
    wire n416, n417, n418, n419, n420, n421, n422, n423;
    wire n424, n425, n426, n427, n428, n429, n430, n431;
    wire n432, n433, n434, n435, n436, n437, n438, n439;
    wire n440, n441, n442, n443, n444, n445, n446, n447;
    wire n448, n449, n450, n451, n452, n453, n454, n455;
    wire n456, n457, n458, n459, n460, n461, n462, n463;
    wire n464, n465, n466, n467, n468, n469, n470, n471;
    wire n472, n473, n474, n475, n476, n477, n478, n479;
    wire n480, n481, n482, n483, n484, n485, n486, n487;
    wire n488, n489, n490, n491, n492, n493, n494, n495;
    wire n496, n497, n498, n499, n500, n501, n502, n503;
    wire n504, n505, n506, n507, n508, n509, n510, n511;
    wire n512, n513, n514, n515, n516, n517, n518, n519;
    wire n520, n521, n522, n523, n524, n525, n526, n527;
    wire n528, n529, n530, n531, n532, n533, n534, n535;
    dff g0(.RN(n1), .SN(1'b1), .CK(n0), .D(n109), .Q(n21[2]));
    dff g1(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[5]), .Q(n30[13]));
    or g2(n416 ,n239 ,n410);
    not g3(n60 ,n30[14]);
    dff g4(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[7]), .Q(n17[7]));
    not g5(n485 ,n18[2]);
    not g6(n186 ,n31[2]);
    xnor g7(n113 ,n2[2] ,n3[2]);
    dff g8(.RN(n1), .SN(1'b1), .CK(n0), .D(n96), .Q(n39[2]));
    xor g9(n138 ,n2[5] ,n3[5]);
    dff g10(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[0]), .Q(n30[8]));
    nor g11(n239 ,n181 ,n214);
    dff g12(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[1]), .Q(n29[3]));
    or g13(n65 ,n53 ,n30[11]);
    dff g14(.RN(n1), .SN(1'b1), .CK(n0), .D(n93), .Q(n40[0]));
    or g15(n529 ,n525 ,n524);
    nor g16(n351 ,n347 ,n343);
    nor g17(n252 ,n194 ,n212);
    nor g18(n259 ,n434 ,n216);
    nor g19(n350 ,n338 ,n336);
    xnor g20(n391 ,n30[0] ,n380);
    xnor g21(n170 ,n121 ,n32[3]);
    not g22(n439 ,n19[3]);
    nor g23(n233 ,n463 ,n212);
    or g24(n68 ,n55 ,n30[0]);
    not g25(n467 ,n22[2]);
    not g26(n474 ,n22[7]);
    nor g27(n227 ,n466 ,n212);
    or g28(n533 ,n530 ,n531);
    dff g29(.RN(n1), .SN(1'b1), .CK(n0), .D(n137), .Q(n15[3]));
    dff g30(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[6]), .Q(n21[6]));
    dff g31(.RN(n1), .SN(1'b1), .CK(n0), .D(n85), .Q(n42[2]));
    nor g32(n242 ,n460 ,n213);
    dff g33(.RN(n1), .SN(1'b1), .CK(n0), .D(n84), .Q(n42[3]));
    dff g34(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[1]), .Q(n25[3]));
    nor g35(n366 ,n356 ,n364);
    xor g36(n131 ,n16[1] ,n39[1]);
    xor g37(n83 ,n43[2] ,n7[0]);
    nor g38(n206 ,n37[0] ,n204);
    not g39(n466 ,n23[7]);
    not g40(n182 ,n32[2]);
    nor g41(n408 ,n209 ,n404);
    dff g42(.RN(n512), .SN(1'b1), .CK(n0), .D(n504), .Q(n47[4]));
    or g43(n201 ,n179 ,n37[1]);
    nor g44(n223 ,n492 ,n208);
    dff g45(.RN(n512), .SN(1'b1), .CK(n0), .D(n506), .Q(n47[2]));
    not g46(n446 ,n15[7]);
    dff g47(.RN(n1), .SN(1'b1), .CK(n0), .D(n142), .Q(n30[7]));
    or g48(n210 ,n37[0] ,n201);
    xor g49(n132 ,n16[0] ,n39[0]);
    not g50(n196 ,n34[4]);
    dff g51(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[5]), .Q(n29[7]));
    nor g52(n229 ,n443 ,n213);
    dff g53(.RN(n1), .SN(1'b1), .CK(n0), .D(n134), .Q(n15[2]));
    not g54(n58 ,n30[7]);
    xnor g55(n370 ,n362 ,n35[1]);
    dff g56(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[7]), .Q(n18[7]));
    dff g57(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[0]), .Q(n28[2]));
    xor g58(n94 ,n34[4] ,n8[4]);
    nor g59(n423 ,n420 ,n421);
    or g60(n323 ,n232 ,n286);
    dff g61(.RN(n1), .SN(1'b1), .CK(n0), .D(n148), .Q(n20[3]));
    not g62(n454 ,n26[3]);
    xnor g63(n381 ,n376 ,n33[3]);
    not g64(n205 ,n204);
    xor g65(n140 ,n2[6] ,n3[6]);
    not g66(n200 ,n199);
    nor g67(n398 ,n25[1] ,n389);
    xor g68(n139 ,n28[1] ,n41[1]);
    xor g69(n361 ,n500 ,n36[3]);
    dff g70(.RN(n1), .SN(1'b1), .CK(n0), .D(n126), .Q(n15[1]));
    dff g71(.RN(n1), .SN(1'b1), .CK(n0), .D(n494), .Q(n10[5]));
    or g72(n405 ,n213 ,n397);
    nor g73(n284 ,n465 ,n215);
    dff g74(.RN(n1), .SN(1'b1), .CK(n0), .D(n99), .Q(n39[0]));
    dff g75(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[2]), .Q(n26[4]));
    dff g76(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[3]), .Q(n22[5]));
    nor g77(n167 ,n63 ,n155);
    xnor g78(n74 ,n8[2] ,n34[2]);
    dff g79(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[3]), .Q(n29[5]));
    or g80(n319 ,n275 ,n223);
    xnor g81(n116 ,n5[1] ,n8[1]);
    not g82(n447 ,n27[3]);
    dff g83(.RN(n1), .SN(1'b1), .CK(n0), .D(n496), .Q(n10[7]));
    buf g84(n11[0], 1'b0);
    xor g85(n126 ,n29[1] ,n40[1]);
    xor g86(n360 ,n497 ,n36[0]);
    nor g87(n357 ,n196 ,n349);
    or g88(n425 ,n407 ,n424);
    or g89(n62 ,n56 ,n30[2]);
    or g90(n399 ,n241 ,n396);
    nor g91(n289 ,n480 ,n215);
    dff g92(.RN(n1), .SN(1'b1), .CK(n0), .D(n92), .Q(n40[1]));
    or g93(n523 ,n501 ,n507);
    nor g94(n402 ,n197 ,n390);
    xnor g95(n163 ,n5[1] ,n125);
    dff g96(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[4]), .Q(n22[6]));
    or g97(n415 ,n251 ,n409);
    dff g98(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[6]), .Q(n30[14]));
    or g99(n154 ,n67 ,n152);
    xnor g100(n117 ,n2[2] ,n3[1]);
    nor g101(n263 ,n487 ,n210);
    xnor g102(n387 ,n32[2] ,n379);
    dff g103(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[0]), .Q(n25[2]));
    xor g104(n171 ,n115 ,n111);
    not g105(n431 ,n29[7]);
    dff g106(.RN(n1), .SN(1'b1), .CK(n0), .D(n105), .Q(n19[3]));
    not g107(n489 ,n17[6]);
    nor g108(n248 ,n474 ,n214);
    not g109(n468 ,n20[1]);
    nor g110(n353 ,n208 ,n351);
    dff g111(.RN(n1), .SN(1'b1), .CK(n0), .D(n98), .Q(n39[1]));
    not g112(n185 ,n31[3]);
    not g113(n469 ,n22[3]);
    xor g114(n85 ,n42[2] ,n4[3]);
    not g115(n519 ,n47[5]);
    xor g116(n105 ,n23[3] ,n45[3]);
    nor g117(n385 ,n255 ,n380);
    or g118(n303 ,n293 ,n273);
    xor g119(n172 ,n122 ,n123);
    xor g120(n96 ,n39[2] ,n9[0]);
    xor g121(n146 ,n25[2] ,n42[2]);
    nor g122(n288 ,n454 ,n215);
    xor g123(n95 ,n39[3] ,n6[0]);
    dff g124(.RN(n1), .SN(1'b1), .CK(n0), .D(n106), .Q(n19[2]));
    not g125(n433 ,n28[2]);
    or g126(n327 ,n247 ,n249);
    not g127(n511 ,n1);
    not g128(n188 ,n34[5]);
    or g129(n531 ,n528 ,n523);
    or g130(n203 ,n178 ,n179);
    dff g131(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[3]), .Q(n16[5]));
    dff g132(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[0]), .Q(n26[2]));
    or g133(n364 ,n211 ,n358);
    dff g134(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[1]), .Q(n16[3]));
    dff g135(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[7]), .Q(n24[7]));
    not g136(n481 ,n14[3]);
    dff g137(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[5]), .Q(n16[7]));
    xor g138(n91 ,n40[2] ,n9[1]);
    xnor g139(n69 ,n6[1] ,n33[1]);
    dff g140(.RN(n1), .SN(1'b1), .CK(n0), .D(n144), .Q(n24[3]));
    xnor g141(n367 ,n359 ,n35[2]);
    not g142(n183 ,n36[2]);
    xnor g143(n389 ,n30[1] ,n382);
    dff g144(.RN(n1), .SN(1'b1), .CK(n0), .D(n135), .Q(n36[1]));
    xor g145(n129 ,n16[3] ,n39[3]);
    dff g146(.RN(n1), .SN(1'b1), .CK(n0), .D(n76), .Q(n35[0]));
    nor g147(n224 ,n486 ,n208);
    dff g148(.RN(n1), .SN(1'b1), .CK(n0), .D(n510), .Q(n38[1]));
    or g149(n530 ,n522 ,n521);
    or g150(n363 ,n211 ,n355);
    xor g151(n133 ,n2[4] ,n3[4]);
    or g152(n428 ,n394 ,n426);
    not g153(n490 ,n16[6]);
    or g154(n318 ,n284 ,n283);
    xor g155(n143 ,n35[1] ,n3[1]);
    xnor g156(n403 ,n387 ,n31[2]);
    dff g157(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[0]), .Q(n23[2]));
    dff g158(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[7]), .Q(n20[7]));
    nor g159(n287 ,n447 ,n210);
    dff g160(.RN(n1), .SN(1'b1), .CK(n0), .D(n139), .Q(n24[1]));
    nor g161(n356 ,n188 ,n351);
    or g162(n209 ,n37[0] ,n205);
    dff g163(.RN(n1), .SN(1'b1), .CK(n0), .D(n110), .Q(n41[1]));
    not g164(n392 ,n391);
    not g165(n192 ,n35[3]);
    nor g166(n218 ,n481 ,n208);
    or g167(n526 ,n513 ,n514);
    or g168(n212 ,n180 ,n202);
    nor g169(n198 ,n178 ,n37[2]);
    dff g170(.RN(n1), .SN(1'b1), .CK(n0), .D(n493), .Q(n10[4]));
    or g171(n215 ,n178 ,n201);
    dff g172(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[2]), .Q(n30[10]));
    or g173(n336 ,n302 ,n296);
    dff g174(.RN(n1), .SN(1'b1), .CK(n0), .D(n500), .Q(n10[3]));
    not g175(n450 ,n17[7]);
    xnor g176(n112 ,n5[3] ,n36[3]);
    or g177(n317 ,n225 ,n280);
    dff g178(.RN(n1), .SN(1'b1), .CK(n0), .D(n79), .Q(n45[3]));
    not g179(n514 ,n508);
    nor g180(n262 ,n453 ,n209);
    or g181(n310 ,n271 ,n268);
    dff g182(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[2]), .Q(n22[4]));
    dff g183(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[5]), .Q(n23[7]));
    xnor g184(n160 ,n5[0] ,n111);
    xnor g185(n175 ,n120 ,n32[2]);
    dff g186(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[6]), .Q(n20[6]));
    dff g187(.RN(n1), .SN(1'b1), .CK(n0), .D(n80), .Q(n45[2]));
    xor g188(n127 ,n46[3] ,n4[7]);
    nor g189(n374 ,n208 ,n369);
    dff g190(.RN(n1), .SN(1'b1), .CK(n0), .D(n145), .Q(n20[1]));
    xor g191(n106 ,n23[2] ,n45[2]);
    xnor g192(n380 ,n378 ,n33[0]);
    not g193(n515 ,n504);
    dff g194(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[3]), .Q(n23[5]));
    dff g195(.RN(n1), .SN(1'b1), .CK(n0), .D(n108), .Q(n21[3]));
    nor g196(n204 ,n180 ,n37[2]);
    or g197(n527 ,n516 ,n515);
    xor g198(n107 ,n34[0] ,n8[0]);
    dff g199(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[6]), .Q(n24[6]));
    not g200(n470 ,n22[6]);
    xor g201(n87 ,n41[3] ,n6[2]);
    or g202(n326 ,n291 ,n224);
    dff g203(.RN(n1), .SN(1'b1), .CK(n0), .D(n175), .Q(n35[2]));
    nor g204(n220 ,n484 ,n208);
    buf g205(n11[1], 1'b0);
    or g206(n208 ,n37[0] ,n200);
    not g207(n55 ,n30[1]);
    xor g208(n92 ,n40[1] ,n4[1]);
    not g209(n478 ,n14[2]);
    dff g210(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[6]), .Q(n18[6]));
    dff g211(.RN(n1), .SN(1'b1), .CK(n0), .D(n101), .Q(n43[3]));
    xnor g212(n368 ,n360 ,n35[0]);
    dff g213(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[2]), .Q(n27[4]));
    nor g214(n354 ,n208 ,n349);
    or g215(n340 ,n328 ,n325);
    nor g216(n244 ,n439 ,n212);
    nor g217(n397 ,n25[0] ,n391);
    nor g218(n228 ,n471 ,n213);
    not g219(n435 ,n16[7]);
    dff g220(.RN(n1), .SN(1'b1), .CK(n0), .D(n130), .Q(n14[2]));
    not g221(n189 ,n25[0]);
    or g222(n329 ,n235 ,n240);
    xnor g223(n118 ,n5[2] ,n8[2]);
    nor g224(n226 ,n477 ,n214);
    xor g225(n142 ,n2[7] ,n3[7]);
    nor g226(n250 ,n193 ,n212);
    or g227(n498 ,n348 ,n346);
    dff g228(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[1]), .Q(n27[3]));
    xnor g229(n157 ,n8[4] ,n73);
    or g230(n300 ,n229 ,n261);
    nor g231(n290 ,n195 ,n210);
    nor g232(n234 ,n470 ,n214);
    nor g233(n247 ,n469 ,n214);
    not g234(n465 ,n21[3]);
    not g235(n434 ,n15[2]);
    or g236(n312 ,n245 ,n230);
    dff g237(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[2]), .Q(n37[2]));
    xnor g238(n114 ,n2[3] ,n3[3]);
    nor g239(n293 ,n440 ,n213);
    not g240(n178 ,n37[0]);
    dff g241(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[11]), .Q(n26[1]));
    xor g242(n88 ,n41[2] ,n4[2]);
    or g243(n315 ,n274 ,n282);
    nor g244(n258 ,n429 ,n216);
    or g245(n499 ,n333 ,n332);
    dff g246(.RN(n1), .SN(1'b1), .CK(n0), .D(n165), .Q(n36[2]));
    not g247(n443 ,n25[6]);
    nor g248(n199 ,n37[2] ,n37[1]);
    buf g249(n12[1], 1'b0);
    not g250(n464 ,n24[7]);
    nor g251(n253 ,n192 ,n214);
    or g252(n155 ,n64 ,n149);
    xor g253(n110 ,n41[1] ,n7[2]);
    or g254(n63 ,n59 ,n30[15]);
    dff g255(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[3]), .Q(n29[1]));
    dff g256(.RN(n1), .SN(1'b1), .CK(n0), .D(n90), .Q(n34[5]));
    nor g257(n249 ,n462 ,n212);
    not g258(n59 ,n30[10]);
    dff g259(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[13]), .Q(n23[1]));
    dff g260(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[2]), .Q(n29[4]));
    xnor g261(n121 ,n3[3] ,n35[3]);
    xor g262(n77 ,n33[2] ,n6[2]);
    not g263(n49 ,n38[1]);
    not g264(n451 ,n27[7]);
    dff g265(.RN(n1), .SN(1'b1), .CK(n0), .D(n138), .Q(n30[5]));
    or g266(n214 ,n180 ,n203);
    dff g267(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[3]), .Q(n25[5]));
    xnor g268(n411 ,n30[3] ,n404);
    not g269(n461 ,n24[6]);
    dff g270(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[1]), .Q(n28[3]));
    dff g271(.RN(n1), .SN(1'b1), .CK(n0), .D(n104), .Q(n18[2]));
    dff g272(.RN(n1), .SN(1'b1), .CK(n0), .D(n497), .Q(n10[0]));
    dff g273(.RN(n1), .SN(1'b1), .CK(n0), .D(n78), .Q(n46[2]));
    or g274(n308 ,n234 ,n233);
    not g275(n492 ,n14[1]);
    xnor g276(n156 ,n8[5] ,n72);
    dff g277(.RN(n1), .SN(1'b1), .CK(n0), .D(n89), .Q(n17[3]));
    xor g278(n150 ,n32[3] ,n31[3]);
    nor g279(n417 ,n25[3] ,n411);
    nor g280(n271 ,n472 ,n215);
    or g281(n213 ,n178 ,n205);
    not g282(n294 ,n293);
    xor g283(n144 ,n28[3] ,n41[3]);
    nor g284(n273 ,n433 ,n209);
    xor g285(n86 ,n42[1] ,n7[3]);
    or g286(n528 ,n503 ,n505);
    or g287(n534 ,n529 ,n532);
    not g288(n484 ,n14[6]);
    not g289(n460 ,n25[7]);
    or g290(n321 ,n289 ,n272);
    xor g291(n141 ,n28[2] ,n41[2]);
    nor g292(n286 ,n449 ,n209);
    dff g293(.RN(n1), .SN(1'b1), .CK(n0), .D(n156), .Q(n26[0]));
    not g294(n455 ,n26[6]);
    xnor g295(n164 ,n112 ,n31[3]);
    nor g296(n222 ,n478 ,n208);
    dff g297(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[5]), .Q(n28[7]));
    dff g298(.RN(n1), .SN(1'b1), .CK(n0), .D(n168), .Q(n34[2]));
    nor g299(n243 ,n488 ,n214);
    xor g300(n82 ,n44[2] ,n7[1]);
    xor g301(n147 ,n40[3] ,n6[1]);
    dff g302(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[7]), .Q(n30[15]));
    xor g303(n90 ,n34[5] ,n8[5]);
    not g304(n52 ,n30[5]);
    xnor g305(n71 ,n6[0] ,n33[0]);
    nor g306(n279 ,n438 ,n216);
    nor g307(n237 ,n187 ,n214);
    not g308(n462 ,n23[3]);
    or g309(n497 ,n341 ,n331);
    dff g310(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[6]), .Q(n17[6]));
    not g311(n480 ,n21[7]);
    not g312(n452 ,n26[2]);
    xor g313(n362 ,n498 ,n36[1]);
    or g314(n325 ,n292 ,n290);
    xor g315(n98 ,n39[1] ,n4[0]);
    nor g316(n352 ,n342 ,n337);
    not g317(n482 ,n20[7]);
    nor g318(n257 ,n441 ,n216);
    nor g319(n230 ,n483 ,n212);
    not g320(n436 ,n28[6]);
    nor g321(n410 ,n402 ,n406);
    not g322(n437 ,n28[7]);
    not g323(n432 ,n17[3]);
    or g324(n522 ,n47[0] ,n47[2]);
    nor g325(n386 ,n255 ,n382);
    not g326(n179 ,n37[2]);
    nor g327(n372 ,n208 ,n368);
    dff g328(.RN(n1), .SN(1'b1), .CK(n0), .D(n169), .Q(n34[3]));
    xnor g329(n413 ,n30[2] ,n403);
    not g330(n412 ,n411);
    dff g331(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[4]), .Q(n25[6]));
    dff g332(.RN(n1), .SN(1'b1), .CK(n0), .D(n509), .Q(n38[2]));
    or g333(n504 ,n354 ,n365);
    xor g334(n174 ,n116 ,n117);
    dff g335(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[15]), .Q(n22[1]));
    not g336(n190 ,n25[3]);
    dff g337(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[1]), .Q(n30[9]));
    xor g338(n76 ,n35[0] ,n3[0]);
    dff g339(.RN(n1), .SN(1'b1), .CK(n0), .D(n159), .Q(n33[0]));
    or g340(n316 ,n242 ,n278);
    nor g341(n277 ,n431 ,n216);
    not g342(n57 ,n38[0]);
    nor g343(n232 ,n468 ,n213);
    nor g344(n283 ,n432 ,n210);
    dff g345(.RN(n1), .SN(1'b1), .CK(n0), .D(n164), .Q(n36[3]));
    nor g346(n407 ,n209 ,n403);
    nor g347(n535 ,n534 ,n533);
    dff g348(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[6]), .Q(n19[6]));
    or g349(n66 ,n58 ,n30[6]);
    nor g350(n240 ,n444 ,n212);
    nor g351(n383 ,n216 ,n379);
    dff g352(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[3]), .Q(n27[5]));
    xnor g353(n73 ,n2[8] ,n3[4]);
    or g354(n216 ,n178 ,n200);
    xor g355(n99 ,n39[0] ,n7[0]);
    or g356(n343 ,n316 ,n313);
    nor g357(n50 ,n38[1] ,n38[0]);
    nor g358(n236 ,n183 ,n212);
    xnor g359(n379 ,n375 ,n33[2]);
    or g360(n427 ,n393 ,n425);
    dff g361(.RN(n512), .SN(1'b1), .CK(n0), .D(n535), .Q(n13));
    or g362(n328 ,n253 ,n252);
    xor g363(n104 ,n22[2] ,n46[2]);
    or g364(n320 ,n246 ,n244);
    dff g365(.RN(n1), .SN(1'b1), .CK(n0), .D(n32[2]), .Q(n11[2]));
    dff g366(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[0]), .Q(n16[2]));
    nor g367(n265 ,n464 ,n209);
    nor g368(n349 ,n334 ,n339);
    not g369(n457 ,n21[2]);
    nor g370(n373 ,n208 ,n370);
    dff g371(.RN(n1), .SN(1'b1), .CK(n0), .D(n495), .Q(n10[6]));
    nor g372(n502 ,n37[2] ,n350);
    nor g373(n280 ,n456 ,n209);
    dff g374(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[4]), .Q(n29[6]));
    dff g375(.RN(n1), .SN(1'b1), .CK(n0), .D(n147), .Q(n40[3]));
    dff g376(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[0]), .Q(n37[0]));
    dff g377(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[2]), .Q(n28[4]));
    or g378(n507 ,n400 ,n416);
    dff g379(.RN(n1), .SN(1'b1), .CK(n0), .D(n97), .Q(n23[0]));
    nor g380(n245 ,n485 ,n214);
    dff g381(.RN(n1), .SN(1'b1), .CK(n0), .D(n160), .Q(n30[0]));
    xor g382(n97 ,n2[12] ,n3[6]);
    xor g383(n78 ,n46[2] ,n7[3]);
    or g384(n302 ,n256 ,n260);
    xnor g385(n375 ,n34[2] ,n367);
    dff g386(.RN(n1), .SN(1'b1), .CK(n0), .D(n94), .Q(n34[4]));
    nor g387(n251 ,n184 ,n212);
    dff g388(.RN(n1), .SN(1'b1), .CK(n0), .D(n170), .Q(n35[3]));
    or g389(n345 ,n320 ,n318);
    xor g390(n134 ,n29[2] ,n40[2]);
    xnor g391(n115 ,n5[0] ,n8[0]);
    not g392(n184 ,n36[0]);
    not g393(n491 ,n15[0]);
    dff g394(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[7]), .Q(n25[1]));
    xor g395(n153 ,n27[2] ,n43[2]);
    or g396(n524 ,n519 ,n518);
    or g397(n67 ,n52 ,n30[4]);
    not g398(n195 ,n32[3]);
    or g399(n505 ,n340 ,n428);
    dff g400(.RN(n1), .SN(1'b1), .CK(n0), .D(n498), .Q(n10[1]));
    dff g401(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[3]), .Q(n26[5]));
    not g402(n516 ,n502);
    or g403(n346 ,n323 ,n319);
    dff g404(.RN(n1), .SN(1'b1), .CK(n0), .D(n129), .Q(n14[3]));
    or g405(n306 ,n226 ,n254);
    or g406(n532 ,n527 ,n526);
    dff g407(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[2]), .Q(n23[4]));
    or g408(n506 ,n335 ,n427);
    xor g409(n84 ,n42[3] ,n6[3]);
    xnor g410(n404 ,n388 ,n31[3]);
    dff g411(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[6]), .Q(n15[6]));
    nor g412(n246 ,n442 ,n214);
    or g413(n149 ,n65 ,n61);
    dff g414(.RN(n1), .SN(1'b1), .CK(n0), .D(n153), .Q(n17[2]));
    not g415(n471 ,n20[2]);
    nor g416(n282 ,n445 ,n210);
    not g417(n517 ,n47[1]);
    dff g418(.RN(n1), .SN(1'b1), .CK(n0), .D(n136), .Q(n36[0]));
    not g419(n496 ,n352);
    xor g420(n93 ,n40[0] ,n7[1]);
    xor g421(n109 ,n26[2] ,n44[2]);
    dff g422(.RN(n512), .SN(1'b1), .CK(n0), .D(n507), .Q(n47[1]));
    nor g423(n256 ,n479 ,n213);
    xnor g424(n122 ,n5[3] ,n8[3]);
    not g425(n187 ,n35[2]);
    nor g426(n501 ,n37[2] ,n352);
    dff g427(.RN(n1), .SN(1'b1), .CK(n0), .D(n57), .Q(n38[0]));
    xnor g428(n165 ,n124 ,n31[2]);
    dff g429(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[7]), .Q(n15[7]));
    not g430(n430 ,n15[1]);
    dff g431(.RN(n1), .SN(1'b1), .CK(n0), .D(n75), .Q(n33[3]));
    nor g432(n358 ,n34[5] ,n494);
    or g433(n152 ,n68 ,n62);
    dff g434(.RN(n1), .SN(1'b1), .CK(n0), .D(n177), .Q(n32[2]));
    dff g435(.RN(n1), .SN(1'b1), .CK(n0), .D(n174), .Q(n29[0]));
    nor g436(n285 ,n459 ,n215);
    xnor g437(n70 ,n8[3] ,n34[3]);
    not g438(n54 ,n30[8]);
    dff g439(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[0]), .Q(n27[2]));
    not g440(n180 ,n37[1]);
    nor g441(n235 ,n467 ,n214);
    xnor g442(n377 ,n34[1] ,n370);
    not g443(n477 ,n18[7]);
    dff g444(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[4]), .Q(n30[12]));
    nor g445(n275 ,n430 ,n216);
    not g446(n191 ,n35[0]);
    nor g447(n238 ,n458 ,n212);
    xnor g448(n72 ,n2[10] ,n3[5]);
    nor g449(n384 ,n216 ,n381);
    dff g450(.RN(n1), .SN(1'b1), .CK(n0), .D(n95), .Q(n39[3]));
    xor g451(n176 ,n32[3] ,n166);
    dff g452(.RN(n1), .SN(1'b1), .CK(n0), .D(n172), .Q(n25[0]));
    dff g453(.RN(n1), .SN(1'b1), .CK(n0), .D(n162), .Q(n30[2]));
    dff g454(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[5]), .Q(n22[7]));
    xnor g455(n376 ,n34[3] ,n369);
    dff g456(.RN(n1), .SN(1'b1), .CK(n0), .D(n158), .Q(n33[1]));
    or g457(n400 ,n250 ,n395);
    nor g458(n267 ,n455 ,n215);
    or g459(n307 ,n270 ,n269);
    not g460(n197 ,n25[1]);
    or g461(n334 ,n308 ,n305);
    nor g462(n221 ,n475 ,n208);
    dff g463(.RN(n512), .SN(1'b1), .CK(n0), .D(n508), .Q(n47[0]));
    not g464(n453 ,n24[2]);
    not g465(n448 ,n27[6]);
    xor g466(n137 ,n29[3] ,n40[3]);
    not g467(n512 ,n511);
    or g468(n344 ,n317 ,n314);
    nor g469(n409 ,n401 ,n405);
    nor g470(n274 ,n452 ,n215);
    nor g471(n211 ,n198 ,n204);
    not g472(n438 ,n15[3]);
    xor g473(n130 ,n16[2] ,n39[2]);
    xnor g474(n158 ,n9[1] ,n69);
    xnor g475(n162 ,n5[2] ,n113);
    xor g476(n89 ,n27[3] ,n43[3]);
    not g477(n193 ,n36[1]);
    nor g478(n424 ,n418 ,n422);
    dff g479(.RN(n1), .SN(1'b1), .CK(n0), .D(n157), .Q(n27[0]));
    not g480(n459 ,n26[7]);
    dff g481(.RN(n1), .SN(1'b1), .CK(n0), .D(n30[3]), .Q(n30[11]));
    xor g482(n509 ,n38[2] ,n51);
    nor g483(n419 ,n294 ,n414);
    not g484(n463 ,n23[6]);
    not g485(n494 ,n351);
    or g486(n314 ,n279 ,n218);
    xor g487(n81 ,n44[3] ,n4[5]);
    or g488(n296 ,n257 ,n220);
    xor g489(n108 ,n26[3] ,n44[3]);
    dff g490(.RN(n1), .SN(1'b1), .CK(n0), .D(n140), .Q(n30[6]));
    not g491(n53 ,n30[12]);
    not g492(n429 ,n29[6]);
    nor g493(n281 ,n451 ,n210);
    nor g494(n219 ,n435 ,n208);
    or g495(n503 ,n353 ,n366);
    or g496(n298 ,n258 ,n217);
    nor g497(n401 ,n189 ,n392);
    or g498(n421 ,n213 ,n417);
    dff g499(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[5]), .Q(n26[7]));
    not g500(n472 ,n21[6]);
    or g501(n330 ,n285 ,n281);
    nor g502(n207 ,n178 ,n199);
    dff g503(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[5]), .Q(n28[1]));
    dff g504(.RN(n1), .SN(1'b1), .CK(n0), .D(n81), .Q(n44[3]));
    dff g505(.RN(n1), .SN(1'b1), .CK(n0), .D(n173), .Q(n28[0]));
    dff g506(.RN(n1), .SN(1'b1), .CK(n0), .D(n132), .Q(n14[0]));
    dff g507(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[4]), .Q(n16[6]));
    dff g508(.RN(n1), .SN(1'b1), .CK(n0), .D(n499), .Q(n10[2]));
    xnor g509(n123 ,n2[6] ,n3[3]);
    or g510(n295 ,n243 ,n238);
    dff g511(.RN(n1), .SN(1'b1), .CK(n0), .D(n100), .Q(n22[0]));
    buf g512(n13, 1'b0);
    or g513(n508 ,n399 ,n415);
    not g514(n456 ,n24[3]);
    not g515(n479 ,n20[6]);
    or g516(n525 ,n517 ,n520);
    or g517(n332 ,n299 ,n297);
    dff g518(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[4]), .Q(n28[6]));
    not g519(n48 ,n38[0]);
    or g520(n396 ,n372 ,n385);
    not g521(n513 ,n506);
    not g522(n475 ,n14[0]);
    dff g523(.RN(n1), .SN(1'b1), .CK(n0), .D(n146), .Q(n20[2]));
    nor g524(n260 ,n461 ,n209);
    not g525(n56 ,n30[3]);
    buf g526(n12[0], 1'b0);
    nor g527(n270 ,n186 ,n215);
    not g528(n487 ,n17[2]);
    nor g529(n51 ,n49 ,n48);
    not g530(n445 ,n27[2]);
    xor g531(n79 ,n45[3] ,n4[6]);
    dff g532(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[5]), .Q(n25[7]));
    not g533(n414 ,n413);
    xnor g534(n159 ,n9[0] ,n71);
    or g535(n339 ,n300 ,n298);
    not g536(n495 ,n350);
    xnor g537(n388 ,n32[3] ,n381);
    xnor g538(n382 ,n377 ,n33[1]);
    nor g539(n225 ,n476 ,n213);
    xor g540(n173 ,n118 ,n119);
    dff g541(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[6]), .Q(n14[6]));
    nor g542(n266 ,n448 ,n210);
    not g543(n483 ,n19[2]);
    dff g544(.RN(n512), .SN(1'b1), .CK(n0), .D(n502), .Q(n47[6]));
    not g545(n440 ,n25[2]);
    nor g546(n292 ,n185 ,n215);
    nor g547(n217 ,n490 ,n208);
    nor g548(n264 ,n457 ,n215);
    or g549(n304 ,n231 ,n265);
    xnor g550(n124 ,n5[2] ,n36[2]);
    nor g551(n231 ,n482 ,n213);
    dff g552(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[7]), .Q(n19[7]));
    nor g553(n365 ,n357 ,n363);
    dff g554(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[4]), .Q(n27[6]));
    dff g555(.RN(n1), .SN(1'b1), .CK(n0), .D(n107), .Q(n34[0]));
    xnor g556(n119 ,n2[4] ,n3[2]);
    dff g557(.RN(n1), .SN(1'b1), .CK(n0), .D(n127), .Q(n46[3]));
    dff g558(.RN(n1), .SN(1'b1), .CK(n0), .D(n171), .Q(n16[0]));
    not g559(n486 ,n14[7]);
    xnor g560(n168 ,n74 ,n31[2]);
    xor g561(n135 ,n36[1] ,n5[1]);
    or g562(n426 ,n408 ,n423);
    nor g563(n510 ,n51 ,n50);
    not g564(n473 ,n19[7]);
    or g565(n64 ,n54 ,n30[9]);
    or g566(n331 ,n303 ,n311);
    not g567(n449 ,n24[1]);
    or g568(n311 ,n276 ,n221);
    dff g569(.RN(n1), .SN(1'b1), .CK(n0), .D(n163), .Q(n30[1]));
    xnor g570(n125 ,n2[1] ,n3[1]);
    dff g571(.RN(n1), .SN(1'b1), .CK(n0), .D(n161), .Q(n30[3]));
    nor g572(n254 ,n473 ,n212);
    nor g573(n241 ,n191 ,n214);
    xnor g574(n161 ,n5[3] ,n114);
    nor g575(n268 ,n489 ,n210);
    xor g576(n359 ,n499 ,n36[2]);
    or g577(n422 ,n213 ,n419);
    dff g578(.RN(n512), .SN(1'b1), .CK(n0), .D(n505), .Q(n47[3]));
    dff g579(.RN(n1), .SN(1'b1), .CK(n0), .D(n32[3]), .Q(n11[3]));
    or g580(n299 ,n228 ,n262);
    nor g581(n166 ,n66 ,n154);
    xor g582(n177 ,n32[2] ,n167);
    or g583(n338 ,n295 ,n310);
    or g584(n348 ,n327 ,n322);
    dff g585(.RN(n512), .SN(1'b1), .CK(n0), .D(n503), .Q(n47[5]));
    dff g586(.RN(n1), .SN(1'b1), .CK(n0), .D(n83), .Q(n43[2]));
    or g587(n342 ,n306 ,n321);
    nor g588(n261 ,n436 ,n209);
    xor g589(n80 ,n45[2] ,n7[2]);
    dff g590(.RN(n1), .SN(1'b1), .CK(n0), .D(n176), .Q(n32[3]));
    xnor g591(n378 ,n34[0] ,n368);
    dff g592(.RN(n1), .SN(1'b1), .CK(n0), .D(n86), .Q(n42[1]));
    or g593(n337 ,n304 ,n326);
    dff g594(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[1]), .Q(n16[1]));
    xor g595(n102 ,n22[3] ,n46[3]);
    or g596(n322 ,n288 ,n287);
    dff g597(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[4]), .Q(n23[6]));
    dff g598(.RN(n1), .SN(1'b1), .CK(n0), .D(n150), .Q(n31[3]));
    not g599(n493 ,n349);
    xor g600(n145 ,n25[1] ,n42[1]);
    or g601(n333 ,n312 ,n301);
    nor g602(n418 ,n293 ,n413);
    dff g603(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[7]), .Q(n14[7]));
    or g604(n335 ,n309 ,n307);
    dff g605(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[7]), .Q(n21[7]));
    or g606(n313 ,n277 ,n219);
    dff g607(.RN(n1), .SN(1'b1), .CK(n0), .D(n2[9]), .Q(n27[1]));
    nor g608(n269 ,n182 ,n210);
    not g609(n520 ,n47[3]);
    or g610(n61 ,n60 ,n30[13]);
    not g611(n181 ,n35[1]);
    dff g612(.RN(n1), .SN(1'b1), .CK(n0), .D(n131), .Q(n14[1]));
    dff g613(.RN(n1), .SN(1'b1), .CK(n0), .D(n128), .Q(n15[0]));
    nor g614(n420 ,n190 ,n412);
    dff g615(.RN(n1), .SN(1'b1), .CK(n0), .D(n151), .Q(n31[2]));
    or g616(n305 ,n267 ,n266);
    dff g617(.RN(n1), .SN(1'b1), .CK(n0), .D(n133), .Q(n30[4]));
    dff g618(.RN(n1), .SN(1'b1), .CK(n0), .D(n29[0]), .Q(n29[2]));
    dff g619(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[1]), .Q(n26[3]));
    dff g620(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[0]), .Q(n22[2]));
    not g621(n444 ,n23[2]);
    or g622(n500 ,n345 ,n344);
    nor g623(n276 ,n491 ,n216);
    not g624(n476 ,n20[3]);
    dff g625(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[2]), .Q(n25[4]));
    or g626(n521 ,n47[4] ,n47[6]);
    dff g627(.RN(n1), .SN(1'b1), .CK(n0), .D(n77), .Q(n33[2]));
    not g628(n390 ,n389);
    dff g629(.RN(n1), .SN(1'b1), .CK(n0), .D(n16[2]), .Q(n16[4]));
    nor g630(n291 ,n446 ,n216);
    not g631(n488 ,n18[6]);
    or g632(n394 ,n374 ,n384);
    nor g633(n272 ,n450 ,n210);
    or g634(n324 ,n248 ,n227);
    dff g635(.RN(n1), .SN(1'b1), .CK(n0), .D(n38[1]), .Q(n37[1]));
    dff g636(.RN(n1), .SN(1'b1), .CK(n0), .D(n28[3]), .Q(n28[5]));
    xor g637(n101 ,n43[3] ,n4[4]);
    or g638(n395 ,n373 ,n386);
    nor g639(n278 ,n437 ,n209);
    xor g640(n151 ,n32[2] ,n31[2]);
    not g641(n194 ,n36[3]);
    or g642(n202 ,n179 ,n37[0]);
    xor g643(n148 ,n25[3] ,n42[3]);
    dff g644(.RN(n512), .SN(1'b1), .CK(n0), .D(n501), .Q(n47[7]));
    or g645(n347 ,n324 ,n330);
    nor g646(n371 ,n208 ,n367);
    nor g647(n355 ,n34[4] ,n493);
    dff g648(.RN(n1), .SN(1'b1), .CK(n0), .D(n82), .Q(n44[2]));
    dff g649(.RN(n1), .SN(1'b1), .CK(n0), .D(n26[4]), .Q(n26[6]));
    xnor g650(n369 ,n361 ,n35[3]);
    dff g651(.RN(n1), .SN(1'b1), .CK(n0), .D(n102), .Q(n18[3]));
    or g652(n301 ,n264 ,n263);
    dff g653(.RN(n1), .SN(1'b1), .CK(n0), .D(n23[1]), .Q(n23[3]));
    xor g654(n103 ,n34[1] ,n8[1]);
    dff g655(.RN(n1), .SN(1'b1), .CK(n0), .D(n22[1]), .Q(n22[3]));
    not g656(n442 ,n18[3]);
    dff g657(.RN(n1), .SN(1'b1), .CK(n0), .D(n143), .Q(n35[1]));
    or g658(n297 ,n259 ,n222);
    or g659(n393 ,n371 ,n383);
    not g660(n441 ,n15[6]);
    xnor g661(n169 ,n70 ,n31[3]);
    or g662(n406 ,n213 ,n398);
    or g663(n341 ,n329 ,n315);
    dff g664(.RN(n1), .SN(1'b1), .CK(n0), .D(n91), .Q(n40[2]));
    dff g665(.RN(n1), .SN(1'b1), .CK(n0), .D(n88), .Q(n41[2]));
    xnor g666(n111 ,n2[0] ,n3[0]);
    xor g667(n75 ,n33[3] ,n6[3]);
    dff g668(.RN(n1), .SN(1'b1), .CK(n0), .D(n87), .Q(n41[3]));
    dff g669(.RN(n1), .SN(1'b1), .CK(n0), .D(n27[5]), .Q(n27[7]));
    not g670(n458 ,n19[6]);
    dff g671(.RN(n1), .SN(1'b1), .CK(n0), .D(n103), .Q(n34[1]));
    xnor g672(n120 ,n3[2] ,n35[2]);
    xor g673(n128 ,n29[0] ,n40[0]);
    or g674(n309 ,n237 ,n236);
    not g675(n518 ,n47[7]);
    dff g676(.RN(n1), .SN(1'b1), .CK(n0), .D(n141), .Q(n24[2]));
    or g677(n255 ,n206 ,n207);
    xor g678(n100 ,n2[14] ,n3[7]);
    xor g679(n136 ,n36[0] ,n5[0]);
endmodule
