module top (n0, n1, n4, n5, n2, n3, n9, n6, n7, n8, n15, n16, n10, n11, n12, n13, n14, n17, n18);
    input n0, n1, n2, n3;
    input [31:0] n4, n5;
    input [3:0] n6;
    input [1:0] n7;
    input [7:0] n8;
    output [31:0] n9, n10, n11, n12, n13, n14;
    output [7:0] n15;
    output [3:0] n16;
    output [15:0] n17, n18;
    wire n0, n1, n2, n3;
    wire [31:0] n4, n5;
    wire [3:0] n6;
    wire [1:0] n7;
    wire [7:0] n8;
    wire [31:0] n9, n10, n11, n12, n13, n14;
    wire [7:0] n15;
    wire [3:0] n16;
    wire [15:0] n17, n18;
    wire [31:0] n19;
    wire [31:0] n20;
    wire [7:0] n21;
    wire [31:0] n22;
    wire [3:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [3:0] n26;
    wire [7:0] n27;
    wire [31:0] n28;
    wire [7:0] n29;
    wire [31:0] n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119;
    or g0(n1553 ,n1462 ,n1461);
    nor g1(n1393 ,n353 ,n1369);
    nor g2(n677 ,n97 ,n610);
    nor g3(n587 ,n433 ,n3);
    nor g4(n919 ,n322 ,n103);
    or g5(n1192 ,n1097 ,n680);
    not g6(n281 ,n5[13]);
    nor g7(n795 ,n402 ,n99);
    or g8(n541 ,n4[9] ,n4[8]);
    nor g9(n1817 ,n193 ,n1446);
    or g10(n535 ,n4[3] ,n4[2]);
    not g11(n214 ,n5[2]);
    or g12(n1275 ,n798 ,n721);
    nor g13(n1667 ,n1107 ,n1445);
    nor g14(n1733 ,n452 ,n1440);
    not g15(n332 ,n20[23]);
    not g16(n304 ,n24[7]);
    or g17(n1301 ,n1099 ,n995);
    or g18(n1963 ,n567 ,n1516);
    nor g19(n957 ,n409 ,n102);
    dff g20(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1882), .Q(n22[15]));
    nor g21(n1769 ,n468 ,n1444);
    nor g22(n709 ,n559 ,n642);
    not g23(n218 ,n28[3]);
    or g24(n876 ,n171 ,n640);
    or g25(n1176 ,n736 ,n1085);
    not g26(n431 ,n9[17]);
    nor g27(n680 ,n2061 ,n106);
    nor g28(n803 ,n519 ,n99);
    not g29(n105 ,n104);
    or g30(n1854 ,n1675 ,n1594);
    dff g31(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1134), .Q(n24[11]));
    nor g32(n986 ,n355 ,n101);
    nor g33(n1337 ,n860 ,n1315);
    not g34(n196 ,n5[25]);
    nor g35(n963 ,n330 ,n103);
    nor g36(n1616 ,n1117 ,n1443);
    or g37(n1252 ,n940 ,n778);
    dff g38(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1222), .Q(n13[20]));
    or g39(n1920 ,n1728 ,n1641);
    not g40(n258 ,n28[11]);
    or g41(n1271 ,n949 ,n1004);
    nor g42(n2065 ,n61 ,n62);
    or g43(n2115 ,n2110 ,n2112);
    or g44(n1892 ,n1699 ,n1621);
    or g45(n1554 ,n1464 ,n1463);
    nor g46(n2072 ,n85 ,n86);
    not g47(n369 ,n25[30]);
    nor g48(n938 ,n219 ,n99);
    or g49(n879 ,n239 ,n640);
    not g50(n251 ,n28[24]);
    nor g51(n1067 ,n159 ,n106);
    dff g52(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1901), .Q(n30[28]));
    or g53(n1996 ,n1775 ,n1836);
    not g54(n490 ,n30[7]);
    or g55(n1322 ,n533 ,n712);
    nor g56(n1604 ,n878 ,n1443);
    dff g57(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1884), .Q(n22[13]));
    nor g58(n1061 ,n163 ,n105);
    or g59(n1869 ,n1338 ,n1828);
    nor g60(n1603 ,n879 ,n1443);
    nor g61(n1477 ,n498 ,n1370);
    nor g62(n1032 ,n363 ,n105);
    not g63(n176 ,n9[9]);
    dff g64(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1905), .Q(n30[24]));
    nor g65(n1612 ,n1108 ,n1443);
    or g66(n1960 ,n1768 ,n1669);
    or g67(n1857 ,n701 ,n1811);
    buf g68(n11[21], n10[21]);
    nor g69(n1397 ,n347 ,n1369);
    buf g70(n12[5], n10[5]);
    or g71(n1446 ,n554 ,n1373);
    or g72(n1331 ,n1269 ,n1267);
    not g73(n141 ,n25[18]);
    not g74(n166 ,n25[11]);
    dff g75(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1261), .Q(n18[2]));
    or g76(n1279 ,n958 ,n1012);
    nor g77(n822 ,n473 ,n102);
    nor g78(n701 ,n638 ,n619);
    or g79(n2010 ,n1803 ,n1850);
    nor g80(n760 ,n300 ,n100);
    nor g81(n907 ,n381 ,n643);
    dff g82(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1176), .Q(n24[6]));
    or g83(n1178 ,n809 ,n1087);
    buf g84(n12[13], n10[13]);
    not g85(n98 ,n97);
    or g86(n2109 ,n2090 ,n2093);
    dff g87(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1939), .Q(n28[22]));
    not g88(n519 ,n10[3]);
    nor g89(n582 ,n204 ,n3);
    not g90(n360 ,n25[8]);
    or g91(n2006 ,n1795 ,n1846);
    or g92(n2118 ,n2111 ,n2117);
    nor g93(n1784 ,n272 ,n1446);
    not g94(n1444 ,n1445);
    dff g95(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1203), .Q(n15[5]));
    or g96(n1190 ,n832 ,n984);
    not g97(n478 ,n9[12]);
    nor g98(n1480 ,n360 ,n1368);
    nor g99(n1613 ,n1118 ,n1443);
    not g100(n456 ,n11[12]);
    or g101(n1316 ,n638 ,n717);
    nor g102(n92 ,n69 ,n90);
    dff g103(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2057), .Q(n25[0]));
    or g104(n885 ,n194 ,n640);
    not g105(n423 ,n9[23]);
    buf g106(n11[28], n10[28]);
    dff g107(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1290), .Q(n10[25]));
    nor g108(n933 ,n501 ,n102);
    not g109(n392 ,n28[30]);
    nor g110(n43 ,n38 ,n42);
    nor g111(n1441 ,n640 ,n1374);
    nor g112(n1692 ,n161 ,n1442);
    dff g113(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1182), .Q(n24[1]));
    nor g114(n1724 ,n463 ,n1440);
    or g115(n875 ,n242 ,n640);
    not g116(n316 ,n24[17]);
    or g117(n1954 ,n1762 ,n1663);
    dff g118(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2013), .Q(n25[12]));
    nor g119(n1685 ,n353 ,n1442);
    dff g120(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1854), .Q(n22[30]));
    not g121(n135 ,n8[1]);
    or g122(n1198 ,n924 ,n771);
    nor g123(n1424 ,n146 ,n1368);
    nor g124(n1456 ,n357 ,n1369);
    nor g125(n837 ,n220 ,n102);
    not g126(n2084 ,n24[19]);
    dff g127(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2038), .Q(n9[12]));
    or g128(n1834 ,n685 ,n1770);
    nor g129(n1503 ,n487 ,n1371);
    nor g130(n661 ,n97 ,n622);
    nor g131(n1681 ,n376 ,n1442);
    or g132(n1530 ,n1408 ,n1409);
    not g133(n252 ,n10[7]);
    nor g134(n846 ,n393 ,n99);
    buf g135(n12[11], n10[11]);
    dff g136(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1201), .Q(n20[11]));
    or g137(n1357 ,n1330 ,n1348);
    nor g138(n1449 ,n514 ,n1370);
    nor g139(n1766 ,n218 ,n1444);
    nor g140(n1455 ,n152 ,n1368);
    not g141(n338 ,n20[20]);
    nor g142(n832 ,n437 ,n102);
    or g143(n1887 ,n1695 ,n1616);
    or g144(n1879 ,n1688 ,n1608);
    dff g145(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1960), .Q(n28[1]));
    not g146(n148 ,n20[1]);
    xnor g147(n595 ,n20[28] ,n24[28]);
    dff g148(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1334), .Q(n15[2]));
    or g149(n1533 ,n1415 ,n1414);
    dff g150(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1133), .Q(n11[2]));
    nor g151(n2068 ,n53 ,n52);
    or g152(n1195 ,n827 ,n1062);
    nor g153(n1344 ,n528 ,n1321);
    or g154(n1937 ,n1745 ,n1591);
    not g155(n469 ,n9[29]);
    or g156(n1157 ,n731 ,n1058);
    nor g157(n703 ,n638 ,n623);
    or g158(n1164 ,n808 ,n1043);
    not g159(n372 ,n22[1]);
    dff g160(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1137), .Q(n10[13]));
    not g161(n306 ,n24[28]);
    or g162(n1171 ,n975 ,n1093);
    not g163(n397 ,n30[1]);
    nor g164(n1693 ,n138 ,n1442);
    dff g165(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1166), .Q(n20[22]));
    dff g166(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1331), .Q(n15[0]));
    or g167(n1175 ,n861 ,n1096);
    nor g168(n1665 ,n1111 ,n1445);
    or g169(n1268 ,n931 ,n1017);
    or g170(n1299 ,n929 ,n1013);
    nor g171(n1501 ,n156 ,n1369);
    not g172(n481 ,n18[3]);
    buf g173(n17[10], n10[2]);
    not g174(n382 ,n22[30]);
    or g175(n2018 ,n1819 ,n1861);
    nor g176(n896 ,n480 ,n99);
    or g177(n552 ,n4[17] ,n4[16]);
    dff g178(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1366), .Q(n23[1]));
    dff g179(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1138), .Q(n20[31]));
    or g180(n2112 ,n2098 ,n2091);
    nor g181(n1660 ,n1116 ,n1445);
    not g182(n122 ,n20[28]);
    nor g183(n1375 ,n137 ,n1365);
    not g184(n267 ,n9[11]);
    not g185(n261 ,n28[22]);
    dff g186(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1305), .Q(n27[6]));
    or g187(n1956 ,n1764 ,n1665);
    nor g188(n1671 ,n885 ,n1441);
    nor g189(n1482 ,n500 ,n1371);
    not g190(n475 ,n30[6]);
    or g191(n2028 ,n1518 ,n1964);
    nor g192(n1006 ,n320 ,n101);
    nor g193(n1661 ,n1105 ,n1441);
    not g194(n472 ,n30[30]);
    or g195(n542 ,n4[11] ,n4[10]);
    or g196(n534 ,n8[1] ,n8[0]);
    xnor g197(n622 ,n20[12] ,n24[12]);
    nor g198(n990 ,n132 ,n96);
    not g199(n601 ,n600);
    not g200(n352 ,n25[5]);
    or g201(n2052 ,n1567 ,n1988);
    xnor g202(n618 ,n20[27] ,n24[27]);
    not g203(n31 ,n29[4]);
    or g204(n1282 ,n817 ,n981);
    dff g205(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1165), .Q(n24[10]));
    dff g206(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1168), .Q(n24[9]));
    not g207(n390 ,n25[9]);
    nor g208(n1422 ,n170 ,n1370);
    or g209(n1110 ,n207 ,n640);
    or g210(n1928 ,n1735 ,n1637);
    dff g211(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1350), .Q(n16[3]));
    nor g212(n1064 ,n149 ,n106);
    dff g213(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1157), .Q(n24[16]));
    nor g214(n947 ,n521 ,n99);
    buf g215(n14[12], n10[8]);
    nor g216(n1037 ,n141 ,n106);
    nor g217(n1495 ,n260 ,n1371);
    nor g218(n974 ,n366 ,n643);
    nor g219(n555 ,n295 ,n109);
    nor g220(n754 ,n312 ,n103);
    dff g221(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2047), .Q(n9[3]));
    or g222(n1125 ,n840 ,n1066);
    or g223(n1130 ,n801 ,n672);
    buf g224(n14[22], n10[18]);
    or g225(n1840 ,n682 ,n1782);
    nor g226(n769 ,n303 ,n101);
    or g227(n1896 ,n1705 ,n1626);
    or g228(n1241 ,n910 ,n1076);
    not g229(n418 ,n30[2]);
    dff g230(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1881), .Q(n22[16]));
    nor g231(n691 ,n638 ,n621);
    or g232(n878 ,n212 ,n640);
    or g233(n1258 ,n954 ,n1083);
    or g234(n2000 ,n1783 ,n1840);
    or g235(n1116 ,n197 ,n640);
    nor g236(n659 ,n97 ,n655);
    or g237(n2007 ,n1797 ,n1847);
    or g238(n1976 ,n582 ,n1542);
    nor g239(n784 ,n304 ,n101);
    nor g240(n972 ,n126 ,n103);
    nor g241(n1803 ,n389 ,n1447);
    nor g242(n954 ,n318 ,n104);
    nor g243(n1019 ,n155 ,n105);
    nor g244(n1448 ,n147 ,n1369);
    not g245(n120 ,n24[30]);
    or g246(n625 ,n564 ,n95);
    or g247(n1167 ,n973 ,n1090);
    or g248(n1835 ,n688 ,n1772);
    or g249(n1837 ,n689 ,n1776);
    or g250(n1184 ,n720 ,n1057);
    nor g251(n1799 ,n183 ,n1446);
    nor g252(n1609 ,n873 ,n1443);
    nor g253(n576 ,n488 ,n3);
    xnor g254(n635 ,n294 ,n148);
    dff g255(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1124), .Q(n11[7]));
    dff g256(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1198), .Q(n12[17]));
    dff g257(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2053), .Q(n9[29]));
    not g258(n117 ,n24[13]);
    nor g259(n674 ,n96 ,n612);
    dff g260(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1912), .Q(n30[17]));
    nor g261(n839 ,n96 ,n595);
    nor g262(n1734 ,n515 ,n1440);
    nor g263(n1731 ,n475 ,n1440);
    nor g264(n785 ,n115 ,n101);
    or g265(n1980 ,n569 ,n1551);
    nor g266(n1605 ,n877 ,n1443);
    dff g267(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2009), .Q(n25[16]));
    not g268(n168 ,n9[18]);
    or g269(n2057 ,n1754 ,n1875);
    or g270(n2054 ,n1571 ,n1990);
    not g271(n230 ,n12[28]);
    nor g272(n1414 ,n240 ,n1370);
    or g273(n631 ,n537 ,n552);
    dff g274(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1903), .Q(n30[26]));
    or g275(n1845 ,n694 ,n1792);
    or g276(n1914 ,n1721 ,n1585);
    or g277(n718 ,n632 ,n631);
    nor g278(n939 ,n396 ,n99);
    dff g279(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1224), .Q(n20[4]));
    nor g280(n1407 ,n263 ,n1371);
    nor g281(n658 ,n97 ,n608);
    or g282(n1147 ,n739 ,n1053);
    not g283(n437 ,n10[6]);
    buf g284(n17[7], 1'b0);
    not g285(n558 ,n557);
    not g286(n313 ,n24[29]);
    nor g287(n1683 ,n363 ,n1442);
    nor g288(n854 ,n208 ,n102);
    nor g289(n1757 ,n202 ,n1444);
    nor g290(n1719 ,n391 ,n1440);
    nor g291(n1017 ,n334 ,n96);
    buf g292(n17[5], 1'b0);
    not g293(n277 ,n5[15]);
    not g294(n136 ,n20[4]);
    nor g295(n849 ,n283 ,n99);
    dff g296(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1216), .Q(n20[7]));
    nor g297(n920 ,n188 ,n102);
    or g298(n1905 ,n1713 ,n1589);
    dff g299(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1194), .Q(n20[15]));
    or g300(n1850 ,n697 ,n1801);
    nor g301(n824 ,n334 ,n103);
    or g302(n1964 ,n566 ,n1519);
    or g303(n589 ,n129 ,n127);
    nor g304(n684 ,n638 ,n603);
    not g305(n383 ,n16[0]);
    nor g306(n1402 ,n391 ,n1371);
    nor g307(n1658 ,n1113 ,n1445);
    or g308(n1133 ,n956 ,n757);
    dff g309(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1308), .Q(n21[3]));
    nor g310(n1419 ,n432 ,n1370);
    nor g311(n1831 ,n349 ,n1447);
    or g312(n1131 ,n794 ,n762);
    or g313(n1186 ,n823 ,n1059);
    nor g314(n1654 ,n1118 ,n1441);
    or g315(n2104 ,n2079 ,n24[6]);
    nor g316(n916 ,n221 ,n98);
    or g317(n1923 ,n1731 ,n1634);
    nor g318(n1702 ,n356 ,n1442);
    not g319(n169 ,n5[29]);
    buf g320(n11[16], n10[16]);
    xnor g321(n623 ,n20[7] ,n24[7]);
    or g322(n1194 ,n824 ,n1061);
    dff g323(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1906), .Q(n30[23]));
    nor g324(n1413 ,n389 ,n1368);
    nor g325(n1730 ,n490 ,n1440);
    not g326(n438 ,n9[3]);
    not g327(n111 ,n24[11]);
    not g328(n268 ,n9[8]);
    nor g329(n1597 ,n1100 ,n1443);
    nor g330(n1650 ,n1113 ,n1441);
    or g331(n1321 ,n523 ,n710);
    nor g332(n695 ,n638 ,n653);
    dff g333(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1120), .Q(n11[10]));
    nor g334(n1680 ,n361 ,n1442);
    nor g335(n1824 ,n368 ,n1447);
    or g336(n34 ,n29[6] ,n29[5]);
    or g337(n1974 ,n574 ,n1538);
    or g338(n1946 ,n1833 ,n1655);
    not g339(n331 ,n21[1]);
    nor g340(n1065 ,n138 ,n105);
    nor g341(n943 ,n513 ,n99);
    dff g342(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1207), .Q(n20[9]));
    or g343(n2049 ,n1561 ,n1985);
    dff g344(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1908), .Q(n30[21]));
    nor g345(n1452 ,n140 ,n1368);
    nor g346(n792 ,n476 ,n99);
    or g347(n1572 ,n1501 ,n1500);
    not g348(n355 ,n16[2]);
    or g349(n1912 ,n1720 ,n1578);
    nor g350(n688 ,n638 ,n597);
    dff g351(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1910), .Q(n30[19]));
    or g352(n1526 ,n1401 ,n1400);
    not g353(n279 ,n13[10]);
    dff g354(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2021), .Q(n25[4]));
    not g355(n216 ,n6[3]);
    nor g356(n726 ,n121 ,n103);
    not g357(n280 ,n13[22]);
    nor g358(n731 ,n315 ,n103);
    not g359(n482 ,n27[5]);
    nor g360(n1723 ,n209 ,n1440);
    nor g361(n1744 ,n249 ,n1444);
    not g362(n248 ,n13[19]);
    nor g363(n1010 ,n328 ,n101);
    or g364(n2114 ,n2107 ,n2109);
    nor g365(n717 ,n649 ,n600);
    nor g366(n1727 ,n445 ,n1440);
    not g367(n476 ,n10[12]);
    nor g368(n1087 ,n353 ,n106);
    or g369(n2025 ,n1577 ,n1993);
    buf g370(n11[29], n10[29]);
    buf g371(n12[4], n10[4]);
    or g372(n522 ,n4[5] ,n4[4]);
    buf g373(n12[0], n10[0]);
    or g374(n1203 ,n899 ,n709);
    nor g375(n683 ,n638 ,n618);
    dff g376(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1855), .Q(n22[31]));
    nor g377(n1493 ,n144 ,n1368);
    or g378(n624 ,n15[1] ,n543);
    dff g379(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1867), .Q(n22[26]));
    or g380(n1163 ,n735 ,n1044);
    dff g381(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1147), .Q(n24[2]));
    or g382(n1847 ,n696 ,n1796);
    nor g383(n1475 ,n372 ,n1369);
    nor g384(n767 ,n315 ,n101);
    nor g385(n1632 ,n1117 ,n1441);
    buf g386(n12[6], n10[6]);
    buf g387(n17[11], n10[3]);
    or g388(n1542 ,n1433 ,n1432);
    nor g389(n1765 ,n416 ,n1444);
    nor g390(n1752 ,n222 ,n1444);
    nor g391(n565 ,n415 ,n3);
    nor g392(n2070 ,n91 ,n92);
    nor g393(n1464 ,n145 ,n1369);
    buf g394(n14[17], n10[13]);
    or g395(n1529 ,n1407 ,n1406);
    or g396(n1319 ,n1060 ,n870);
    nor g397(n1676 ,n139 ,n1442);
    nor g398(n1458 ,n475 ,n1371);
    nor g399(n1806 ,n281 ,n1446);
    dff g400(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1186), .Q(n20[16]));
    or g401(n1998 ,n1777 ,n1837);
    or g402(n1267 ,n788 ,n1003);
    or g403(n1910 ,n1718 ,n1582);
    nor g404(n1339 ,n848 ,n1313);
    nor g405(n662 ,n96 ,n620);
    or g406(n1101 ,n253 ,n640);
    or g407(n1565 ,n1487 ,n1486);
    or g408(n1129 ,n963 ,n1055);
    or g409(n1945 ,n1753 ,n1579);
    or g410(n2032 ,n1527 ,n1968);
    dff g411(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1258), .Q(n20[27]));
    not g412(n134 ,n20[10]);
    dff g413(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2005), .Q(n25[20]));
    or g414(n2021 ,n1825 ,n1866);
    not g415(n312 ,n24[8]);
    dff g416(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2011), .Q(n25[14]));
    nor g417(n1641 ,n1116 ,n1441);
    nor g418(n823 ,n324 ,n103);
    or g419(n1545 ,n1436 ,n1437);
    nor g420(n787 ,n111 ,n96);
    dff g421(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2012), .Q(n25[13]));
    or g422(n2095 ,n2084 ,n24[18]);
    not g423(n292 ,n2065);
    dff g424(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1930), .Q(n28[31]));
    nor g425(n640 ,n293 ,n553);
    nor g426(n863 ,n131 ,n103);
    dff g427(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1945), .Q(n28[16]));
    or g428(n1541 ,n1431 ,n1430);
    nor g429(n805 ,n328 ,n103);
    or g430(n1948 ,n1756 ,n1657);
    not g431(n236 ,n11[3]);
    or g432(n1531 ,n1411 ,n1410);
    not g433(n272 ,n5[24]);
    nor g434(n1819 ,n184 ,n1446);
    nor g435(n1400 ,n141 ,n1368);
    dff g436(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1195), .Q(n20[13]));
    not g437(n219 ,n10[22]);
    dff g438(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2023), .Q(n25[2]));
    not g439(n96 ,n99);
    not g440(n363 ,n22[22]);
    nor g441(n1583 ,n877 ,n1441);
    or g442(n1360 ,n711 ,n1352);
    nor g443(n1325 ,n640 ,n864);
    nor g444(n1403 ,n227 ,n1370);
    nor g445(n681 ,n638 ,n605);
    nor g446(n995 ,n325 ,n101);
    not g447(n298 ,n24[2]);
    dff g448(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1298), .Q(n10[21]));
    or g449(n1280 ,n816 ,n980);
    nor g450(n1601 ,n880 ,n1443);
    not g451(n513 ,n10[19]);
    nor g452(n971 ,n276 ,n99);
    nor g453(n1081 ,n162 ,n106);
    nor g454(n1633 ,n1114 ,n1441);
    nor g455(n1596 ,n883 ,n1441);
    or g456(n543 ,n15[2] ,n15[3]);
    not g457(n509 ,n14[0]);
    or g458(n1232 ,n900 ,n674);
    dff g459(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2041), .Q(n9[9]));
    or g460(n1883 ,n1691 ,n1612);
    nor g461(n1735 ,n418 ,n1440);
    nor g462(n1417 ,n149 ,n1369);
    not g463(n127 ,n4[2]);
    or g464(n2046 ,n1555 ,n1983);
    or g465(n1970 ,n580 ,n1530);
    buf g466(n14[18], n10[14]);
    nor g467(n88 ,n29[5] ,n86);
    or g468(n712 ,n15[0] ,n624);
    nor g469(n918 ,n413 ,n102);
    not g470(n424 ,n13[20]);
    or g471(n1159 ,n727 ,n1034);
    nor g472(n1487 ,n495 ,n1371);
    nor g473(n771 ,n316 ,n96);
    not g474(n435 ,n12[17]);
    or g475(n1539 ,n1427 ,n1426);
    not g476(n48 ,n27[3]);
    or g477(n1873 ,n1682 ,n1603);
    nor g478(n819 ,n333 ,n104);
    or g479(n1255 ,n919 ,n1078);
    nor g480(n566 ,n504 ,n3);
    not g481(n479 ,n27[7]);
    nor g482(n801 ,n510 ,n102);
    or g483(n647 ,n539 ,n522);
    nor g484(n1753 ,n430 ,n1444);
    dff g485(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2033), .Q(n9[17]));
    not g486(n324 ,n20[16]);
    not g487(n320 ,n20[13]);
    or g488(n1153 ,n923 ,n1030);
    or g489(n1852 ,n699 ,n1806);
    or g490(n1283 ,n888 ,n983);
    not g491(n393 ,n11[11]);
    nor g492(n1647 ,n1109 ,n1441);
    nor g493(n851 ,n101 ,n602);
    buf g494(n18[11], 1'b0);
    not g495(n374 ,n22[0]);
    or g496(n1952 ,n1760 ,n1660);
    nor g497(n1645 ,n882 ,n1445);
    nor g498(n730 ,n118 ,n103);
    not g499(n108 ,n24[0]);
    nor g500(n82 ,n29[3] ,n80);
    nor g501(n1773 ,n178 ,n1446);
    or g502(n2016 ,n1815 ,n1858);
    nor g503(n1690 ,n163 ,n1442);
    or g504(n1306 ,n828 ,n985);
    not g505(n368 ,n25[4]);
    dff g506(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2070), .Q(n29[6]));
    or g507(n44 ,n27[7] ,n43);
    nor g508(n1406 ,n222 ,n1370);
    or g509(n1281 ,n935 ,n979);
    nor g510(n794 ,n516 ,n99);
    not g511(n188 ,n13[27]);
    nor g512(n780 ,n121 ,n100);
    dff g513(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1244), .Q(n12[20]));
    nor g514(n1461 ,n231 ,n1370);
    nor g515(n741 ,n296 ,n103);
    or g516(n1274 ,n792 ,n976);
    or g517(n1135 ,n797 ,n722);
    nor g518(n1093 ,n292 ,n638);
    dff g519(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2056), .Q(n9[26]));
    not g520(n241 ,n11[7]);
    dff g521(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1359), .Q(n23[2]));
    not g522(n132 ,n20[29]);
    nor g523(n912 ,n245 ,n98);
    dff g524(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1131), .Q(n11[4]));
    or g525(n2100 ,n2076 ,n2077);
    xnor g526(n653 ,n20[19] ,n24[19]);
    not g527(n2085 ,n24[12]);
    dff g528(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1141), .Q(n24[28]));
    nor g529(n1054 ,n349 ,n106);
    nor g530(n1459 ,n351 ,n1369);
    not g531(n174 ,n12[18]);
    nor g532(n900 ,n455 ,n102);
    nor g533(n835 ,n517 ,n102);
    or g534(n1560 ,n1475 ,n1476);
    dff g535(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1193), .Q(n11[8]));
    nor g536(n838 ,n128 ,n103);
    or g537(n529 ,n4[29] ,n4[28]);
    or g538(n2013 ,n1809 ,n1853);
    dff g539(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1171), .Q(n27[4]));
    or g540(n1361 ,n1353 ,n1352);
    nor g541(n2064 ,n64 ,n65);
    nor g542(n1779 ,n253 ,n1446);
    nor g543(n1091 ,n287 ,n638);
    dff g544(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2054), .Q(n9[28]));
    or g545(n1247 ,n950 ,n772);
    or g546(n1971 ,n577 ,n1532);
    dff g547(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2015), .Q(n25[10]));
    or g548(n1842 ,n691 ,n1786);
    or g549(n1304 ,n854 ,n1016);
    not g550(n333 ,n20[17]);
    or g551(n1270 ,n947 ,n992);
    nor g552(n1051 ,n368 ,n106);
    xnor g553(n619 ,n20[10] ,n24[10]);
    not g554(n299 ,n24[19]);
    nor g555(n1711 ,n425 ,n1440);
    not g556(n353 ,n22[20]);
    not g557(n351 ,n22[5]);
    nor g558(n797 ,n250 ,n102);
    dff g559(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1220), .Q(n13[21]));
    not g560(n167 ,n6[2]);
    nor g561(n906 ,n429 ,n102);
    not g562(n253 ,n5[26]);
    or g563(n2105 ,n2089 ,n2096);
    nor g564(n568 ,n168 ,n3);
    nor g565(n62 ,n47 ,n60);
    nor g566(n1405 ,n274 ,n1371);
    buf g567(n17[15], n10[7]);
    or g568(n1292 ,n951 ,n1007);
    nor g569(n585 ,n422 ,n3);
    or g570(n1922 ,n1730 ,n1633);
    dff g571(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1864), .Q(n22[27]));
    not g572(n231 ,n28[5]);
    not g573(n470 ,n12[23]);
    not g574(n1440 ,n1441);
    or g575(n867 ,n641 ,n102);
    not g576(n2078 ,n24[3]);
    nor g577(n810 ,n205 ,n99);
    nor g578(n1751 ,n227 ,n1444);
    nor g579(n1762 ,n175 ,n1444);
    nor g580(n1756 ,n170 ,n1444);
    or g581(n1251 ,n748 ,n1082);
    not g582(n645 ,n644);
    not g583(n206 ,n6[1]);
    not g584(n270 ,n9[24]);
    nor g585(n670 ,n96 ,n594);
    dff g586(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2027), .Q(n9[23]));
    nor g587(n1433 ,n378 ,n1369);
    or g588(n1257 ,n641 ,n891);
    dff g589(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1877), .Q(n22[20]));
    nor g590(n2066 ,n58 ,n59);
    nor g591(n940 ,n470 ,n102);
    nor g592(n755 ,n312 ,n101);
    dff g593(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2039), .Q(n9[11]));
    nor g594(n1338 ,n850 ,n1314);
    not g595(n151 ,n25[24]);
    dff g596(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1286), .Q(n12[26]));
    nor g597(n1418 ,n209 ,n1371);
    not g598(n516 ,n11[4]);
    nor g599(n1821 ,n211 ,n1446);
    nor g600(n1640 ,n1103 ,n1441);
    or g601(n634 ,n8[1] ,n527);
    or g602(n1309 ,n852 ,n994);
    or g603(n1260 ,n641 ,n855);
    not g604(n430 ,n28[16]);
    or g605(n1917 ,n1725 ,n1650);
    not g606(n370 ,n16[1]);
    nor g607(n1659 ,n1117 ,n1445);
    not g608(n276 ,n11[13]);
    nor g609(n1708 ,n260 ,n1440);
    not g610(n263 ,n30[17]);
    not g611(n518 ,n10[24]);
    not g612(n594 ,n593);
    or g613(n1872 ,n1337 ,n1830);
    nor g614(n1030 ,n377 ,n105);
    or g615(n1907 ,n1715 ,n1629);
    not g616(n289 ,n7[1]);
    not g617(n226 ,n10[18]);
    nor g618(n913 ,n339 ,n103);
    not g619(n394 ,n13[24]);
    nor g620(n1497 ,n387 ,n1369);
    or g621(n1226 ,n964 ,n677);
    nor g622(n815 ,n426 ,n99);
    or g623(n1535 ,n1418 ,n1419);
    dff g624(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1208), .Q(n13[31]));
    nor g625(n1342 ,n641 ,n1317);
    not g626(n428 ,n13[31]);
    dff g627(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1127), .Q(n21[1]));
    or g628(n1189 ,n926 ,n671);
    not g629(n389 ,n25[15]);
    dff g630(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1311), .Q(n11[12]));
    or g631(n1859 ,n702 ,n1816);
    nor g632(n776 ,n110 ,n96);
    nor g633(n1506 ,n425 ,n1371);
    or g634(n1204 ,n745 ,n1035);
    dff g635(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1129), .Q(n21[0]));
    not g636(n239 ,n5[23]);
    or g637(n2107 ,n2095 ,n2101);
    dff g638(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2004), .Q(n25[21]));
    not g639(n309 ,n24[23]);
    or g640(n1961 ,n1769 ,n1670);
    nor g641(n685 ,n638 ,n602);
    dff g642(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1199), .Q(n11[15]));
    or g643(n1273 ,n799 ,n1005);
    dff g644(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1128), .Q(n11[5]));
    or g645(n1527 ,n1402 ,n1403);
    or g646(n1844 ,n693 ,n1791);
    or g647(n1183 ,n814 ,n1052);
    not g648(n308 ,n24[31]);
    buf g649(n18[7], n14[7]);
    dff g650(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1123), .Q(n10[28]));
    or g651(n1944 ,n1752 ,n1584);
    dff g652(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2019), .Q(n25[6]));
    nor g653(n86 ,n71 ,n84);
    or g654(n1856 ,n686 ,n1810);
    or g655(n39 ,n27[4] ,n27[3]);
    nor g656(n764 ,n307 ,n101);
    nor g657(n2119 ,n2114 ,n2118);
    or g658(n2037 ,n1537 ,n1973);
    dff g659(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1994), .Q(n25[31]));
    or g660(n1240 ,n921 ,n668);
    not g661(n184 ,n5[7]);
    nor g662(n1691 ,n149 ,n1442);
    or g663(n1915 ,n1722 ,n1661);
    dff g664(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1179), .Q(n26[0]));
    nor g665(n1062 ,n161 ,n106);
    nor g666(n790 ,n110 ,n645);
    nor g667(n1642 ,n884 ,n1445);
    not g668(n380 ,n25[26]);
    nor g669(n679 ,n96 ,n654);
    dff g670(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1938), .Q(n28[23]));
    or g671(n2113 ,n2106 ,n2105);
    or g672(n1523 ,n1395 ,n1394);
    nor g673(n762 ,n118 ,n100);
    or g674(n1172 ,n750 ,n1084);
    or g675(n1154 ,n741 ,n1037);
    nor g676(n549 ,n270 ,n3);
    or g677(n633 ,n544 ,n531);
    nor g678(n721 ,n108 ,n100);
    nor g679(n1426 ,n202 ,n1370);
    dff g680(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1942), .Q(n28[19]));
    or g681(n637 ,n589 ,n95);
    or g682(n2031 ,n1525 ,n1967);
    not g683(n295 ,n23[0]);
    nor g684(n1386 ,n261 ,n1370);
    not g685(n2080 ,n24[23]);
    or g686(n1933 ,n1743 ,n1646);
    nor g687(n36 ,n31 ,n35);
    nor g688(n1581 ,n876 ,n1441);
    nor g689(n1060 ,n172 ,n105);
    nor g690(n1755 ,n432 ,n1444);
    or g691(n1269 ,n641 ,n907);
    dff g692(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2050), .Q(n9[0]));
    dff g693(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2001), .Q(n25[24]));
    nor g694(n910 ,n323 ,n103);
    or g695(n1969 ,n586 ,n1528);
    nor g696(n1578 ,n873 ,n1441);
    not g697(n395 ,n12[22]);
    nor g698(n1389 ,n162 ,n1368);
    or g699(n2099 ,n2080 ,n24[22]);
    nor g700(n1678 ,n156 ,n1442);
    or g701(n1546 ,n1448 ,n1480);
    dff g702(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1219), .Q(n13[22]));
    nor g703(n56 ,n51 ,n54);
    nor g704(n1018 ,n136 ,n96);
    or g705(n1358 ,n1328 ,n1346);
    dff g706(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1243), .Q(n13[3]));
    or g707(n2019 ,n1821 ,n1863);
    not g708(n278 ,n12[19]);
    dff g709(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1289), .Q(n10[26]));
    nor g710(n1630 ,n874 ,n1441);
    nor g711(n765 ,n120 ,n101);
    nor g712(n1602 ,n1100 ,n1441);
    nor g713(n1069 ,n342 ,n105);
    or g714(n2117 ,n2108 ,n2116);
    nor g715(n902 ,n400 ,n102);
    not g716(n514 ,n28[8]);
    buf g717(n18[13], n10[1]);
    or g718(n1213 ,n920 ,n836);
    dff g719(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2000), .Q(n25[25]));
    or g720(n531 ,n4[25] ,n4[24]);
    or g721(n1561 ,n1478 ,n1477);
    nor g722(n808 ,n332 ,n103);
    dff g723(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1281), .Q(n10[31]));
    or g724(n1160 ,n753 ,n1086);
    dff g725(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1284), .Q(n10[29]));
    nor g726(n1826 ,n348 ,n1447);
    xnor g727(n620 ,n20[11] ,n24[11]);
    nor g728(n671 ,n97 ,n592);
    dff g729(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1302), .Q(n14[6]));
    or g730(n1298 ,n933 ,n999);
    not g731(n192 ,n6[0]);
    nor g732(n1745 ,n251 ,n1444);
    nor g733(n1384 ,n154 ,n1368);
    buf g734(n17[3], n14[7]);
    not g735(n133 ,n20[26]);
    dff g736(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1892), .Q(n22[5]));
    dff g737(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1119), .Q(n27[0]));
    not g738(n398 ,n9[27]);
    nor g739(n1471 ,n143 ,n1368);
    or g740(n2004 ,n1790 ,n1844);
    nor g741(n1649 ,n878 ,n1445);
    not g742(n447 ,n30[28]);
    or g743(n20[0] ,n19[0] ,n2119);
    not g744(n100 ,n102);
    not g745(n377 ,n22[26]);
    dff g746(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1911), .Q(n30[18]));
    nor g747(n1002 ,n164 ,n96);
    dff g748(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1246), .Q(n12[31]));
    nor g749(n1411 ,n265 ,n1371);
    nor g750(n789 ,n300 ,n638);
    not g751(n408 ,n30[8]);
    xnor g752(n605 ,n20[24] ,n24[24]);
    nor g753(n548 ,n474 ,n3);
    dff g754(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1142), .Q(n24[27]));
    nor g755(n65 ,n50 ,n63);
    not g756(n450 ,n9[7]);
    or g757(n1263 ,n641 ,n986);
    not g758(n434 ,n9[1]);
    nor g759(n1028 ,n153 ,n105);
    nor g760(n752 ,n303 ,n104);
    not g761(n142 ,n22[7]);
    dff g762(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1292), .Q(n10[24]));
    or g763(n2102 ,n2088 ,n24[24]);
    nor g764(n953 ,n271 ,n102);
    xnor g765(n603 ,n20[29] ,n24[29]);
    nor g766(n796 ,n336 ,n104);
    dff g767(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1934), .Q(n28[28]));
    or g768(n1205 ,n862 ,n760);
    nor g769(n1599 ,n1101 ,n1443);
    not g770(n362 ,n22[23]);
    not g771(n442 ,n11[9]);
    buf g772(n17[2], n14[6]);
    or g773(n1307 ,n849 ,n988);
    or g774(n2002 ,n1787 ,n1842);
    or g775(n630 ,n540 ,n529);
    or g776(n1256 ,n897 ,n775);
    or g777(n2094 ,n2087 ,n24[26]);
    or g778(n544 ,n4[27] ,n4[26]);
    nor g779(n1673 ,n1115 ,n1441);
    dff g780(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1926), .Q(n30[4]));
    nor g781(n917 ,n512 ,n102);
    or g782(n881 ,n196 ,n640);
    nor g783(n905 ,n327 ,n103);
    not g784(n480 ,n13[14]);
    not g785(n254 ,n5[11]);
    not g786(n2079 ,n24[7]);
    nor g787(n1825 ,n207 ,n1446);
    or g788(n1140 ,n724 ,n1022);
    or g789(n1522 ,n1393 ,n1392);
    or g790(n1145 ,n829 ,n1024);
    or g791(n1886 ,n1694 ,n1615);
    or g792(n1246 ,n835 ,n761);
    or g793(n1836 ,n684 ,n1774);
    nor g794(n1582 ,n875 ,n1441);
    or g795(n1867 ,n1679 ,n1599);
    dff g796(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1318), .Q(n13[19]));
    not g797(n113 ,n24[9]);
    or g798(n1550 ,n1458 ,n1457);
    not g799(n325 ,n20[18]);
    nor g800(n719 ,n294 ,n103);
    nor g801(n734 ,n114 ,n104);
    or g802(n1199 ,n969 ,n768);
    or g803(n1318 ,n887 ,n678);
    or g804(n1102 ,n200 ,n640);
    dff g805(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1909), .Q(n30[20]));
    or g806(n1959 ,n1767 ,n1668);
    nor g807(n687 ,n638 ,n610);
    not g808(n401 ,n10[4]);
    nor g809(n728 ,n117 ,n103);
    dff g810(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2006), .Q(n25[19]));
    or g811(n1132 ,n961 ,n785);
    nor g812(n1392 ,n346 ,n1368);
    dff g813(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1260), .Q(n15[4]));
    nor g814(n723 ,n314 ,n104);
    not g815(n144 ,n25[29]);
    nor g816(n949 ,n403 ,n102);
    buf g817(n18[5], n14[5]);
    not g818(n407 ,n10[1]);
    not g819(n403 ,n10[14]);
    not g820(n294 ,n24[1]);
    dff g821(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1303), .Q(n27[5]));
    dff g822(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1919), .Q(n30[10]));
    not g823(n650 ,n649);
    dff g824(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1122), .Q(n11[9]));
    not g825(n2081 ,n24[14]);
    nor g826(n1634 ,n1112 ,n1441);
    dff g827(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1173), .Q(n20[19]));
    or g828(n1868 ,n1339 ,n1826);
    not g829(n162 ,n25[21]);
    or g830(n1235 ,n908 ,n663);
    dff g831(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1920), .Q(n30[9]));
    dff g832(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1214), .Q(n13[26]));
    or g833(n1155 ,n807 ,n1039);
    or g834(n2014 ,n1812 ,n1856);
    not g835(n410 ,n14[5]);
    dff g836(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2007), .Q(n25[18]));
    dff g837(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1125), .Q(n21[2]));
    nor g838(n682 ,n638 ,n604);
    nor g839(n1380 ,n362 ,n1369);
    nor g840(n639 ,n23[2] ,n553);
    dff g841(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1256), .Q(n12[19]));
    or g842(n1231 ,n896 ,n660);
    nor g843(n667 ,n97 ,n613);
    or g844(n1897 ,n1707 ,n1627);
    nor g845(n976 ,n326 ,n100);
    nor g846(n1770 ,n194 ,n1446);
    not g847(n381 ,n15[0]);
    nor g848(n1080 ,n359 ,n106);
    not g849(n436 ,n13[12]);
    nor g850(n774 ,n296 ,n101);
    not g851(n224 ,n27[6]);
    buf g852(n12[14], n10[14]);
    nor g853(n1688 ,n384 ,n1442);
    or g854(n1927 ,n1734 ,n1636);
    nor g855(n975 ,n266 ,n639);
    not g856(n1345 ,n1344);
    nor g857(n1425 ,n138 ,n1369);
    or g858(n1543 ,n1434 ,n1435);
    or g859(n1999 ,n1781 ,n1839);
    or g860(n1984 ,n563 ,n1558);
    or g861(n1294 ,n952 ,n1009);
    nor g862(n915 ,n484 ,n98);
    nor g863(n58 ,n27[3] ,n56);
    nor g864(n1008 ,n318 ,n96);
    or g865(n1557 ,n1470 ,n1469);
    or g866(n1211 ,n872 ,n843);
    nor g867(n1009 ,n148 ,n101);
    not g868(n73 ,n29[1]);
    nor g869(n844 ,n326 ,n103);
    not g870(n346 ,n25[20]);
    not g871(n433 ,n9[13]);
    not g872(n409 ,n10[26]);
    not g873(n211 ,n5[6]);
    nor g874(n1056 ,n365 ,n106);
    nor g875(n783 ,n311 ,n97);
    nor g876(n1092 ,n291 ,n638);
    dff g877(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1184), .Q(n24[0]));
    or g878(n1564 ,n1484 ,n1485);
    not g879(n256 ,n10[2]);
    or g880(n2091 ,n24[1] ,n24[0]);
    not g881(n454 ,n11[14]);
    or g882(n1121 ,n960 ,n769);
    nor g883(n55 ,n27[2] ,n53);
    nor g884(n961 ,n236 ,n102);
    or g885(n1978 ,n579 ,n1546);
    nor g886(n816 ,n180 ,n99);
    nor g887(n1709 ,n447 ,n1440);
    or g888(n2008 ,n1799 ,n1848);
    dff g889(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1297), .Q(n27[3]));
    not g890(n109 ,n23[1]);
    nor g891(n1070 ,n147 ,n105);
    not g892(n356 ,n22[3]);
    nor g893(n590 ,n434 ,n3);
    dff g894(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1202), .Q(n20[10]));
    nor g895(n1026 ,n344 ,n106);
    buf g896(n12[8], n10[8]);
    or g897(n1367 ,n1192 ,n1360);
    buf g898(n18[6], n14[6]);
    nor g899(n672 ,n97 ,n636);
    buf g900(n17[14], n10[6]);
    xnor g901(n649 ,n108 ,n19[0]);
    nor g902(n1794 ,n242 ,n1446);
    not g903(n152 ,n25[6]);
    xnor g904(n606 ,n20[6] ,n24[6]);
    buf g905(n11[17], n10[17]);
    xnor g906(n596 ,n20[22] ,n24[22]);
    nor g907(n751 ,n310 ,n104);
    dff g908(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1873), .Q(n22[23]));
    not g909(n97 ,n99);
    nor g910(n770 ,n314 ,n101);
    not g911(n426 ,n11[5]);
    dff g912(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1299), .Q(n14[7]));
    nor g913(n1000 ,n133 ,n101);
    or g914(n2089 ,n24[11] ,n24[10]);
    or g915(n1875 ,n1336 ,n1832);
    or g916(n1979 ,n572 ,n1548);
    nor g917(n1813 ,n354 ,n1447);
    not g918(n121 ,n24[22]);
    dff g919(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1300), .Q(n10[19]));
    or g920(n2015 ,n1813 ,n1857);
    not g921(n237 ,n28[10]);
    nor g922(n91 ,n29[6] ,n89);
    or g923(n1314 ,n638 ,n713);
    not g924(n319 ,n20[11]);
    not g925(n326 ,n20[12]);
    or g926(n1935 ,n1742 ,n1645);
    nor g927(n904 ,n436 ,n99);
    not g928(n2083 ,n24[21]);
    nor g929(n1372 ,n137 ,n1363);
    nor g930(n1614 ,n1113 ,n1443);
    or g931(n530 ,n15[4] ,n15[5]);
    nor g932(n1488 ,n369 ,n1368);
    or g933(n1180 ,n734 ,n1041);
    not g934(n66 ,n65);
    dff g935(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1234), .Q(n13[11]));
    nor g936(n748 ,n308 ,n104);
    or g937(n1851 ,n698 ,n1804);
    nor g938(n750 ,n304 ,n103);
    dff g939(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1358), .Q(n16[1]));
    or g940(n1254 ,n930 ,n998);
    not g941(n386 ,n25[16]);
    buf g942(n12[10], n10[10]);
    nor g943(n79 ,n29[2] ,n77);
    or g944(n1215 ,n915 ,n856);
    not g945(n90 ,n89);
    or g946(n1908 ,n1716 ,n1583);
    not g947(n343 ,n22[21]);
    buf g948(n14[14], n10[10]);
    nor g949(n1491 ,n472 ,n1371);
    nor g950(n743 ,n316 ,n104);
    not g951(n161 ,n22[13]);
    not g952(n190 ,n13[9]);
    not g953(n384 ,n22[18]);
    dff g954(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1190), .Q(n10[6]));
    dff g955(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1944), .Q(n28[17]));
    dff g956(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1940), .Q(n28[21]));
    nor g957(n1592 ,n882 ,n1441);
    not g958(n232 ,n13[18]);
    or g959(n1158 ,n805 ,n1033);
    nor g960(n998 ,n210 ,n101);
    nor g961(n1039 ,n376 ,n105);
    or g962(n2022 ,n1827 ,n1868);
    dff g963(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1891), .Q(n22[6]));
    or g964(n1182 ,n719 ,n1054);
    buf g965(n18[15], n10[3]);
    nor g966(n775 ,n299 ,n96);
    nor g967(n834 ,n401 ,n102);
    nor g968(n1084 ,n140 ,n105);
    not g969(n60 ,n59);
    nor g970(n950 ,n506 ,n99);
    or g971(n1202 ,n871 ,n1068);
    not g972(n63 ,n62);
    not g973(n225 ,n5[5]);
    or g974(n2005 ,n1793 ,n1845);
    not g975(n477 ,n10[29]);
    or g976(n1558 ,n1472 ,n1471);
    dff g977(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1146), .Q(n24[24]));
    nor g978(n1695 ,n378 ,n1442);
    or g979(n95 ,n4[1] ,n4[0]);
    dff g980(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1239), .Q(n13[6]));
    nor g981(n1754 ,n247 ,n1446);
    nor g982(n956 ,n483 ,n99);
    dff g983(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1189), .Q(n13[2]));
    dff g984(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1235), .Q(n13[10]));
    not g985(n471 ,n13[5]);
    dff g986(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1164), .Q(n20[23]));
    nor g987(n1721 ,n265 ,n1440);
    nor g988(n583 ,n421 ,n3);
    nor g989(n1589 ,n880 ,n1441);
    or g990(n2061 ,n34 ,n37);
    nor g991(n665 ,n97 ,n623);
    or g992(n1149 ,n726 ,n1029);
    not g993(n70 ,n29[0]);
    dff g994(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1152), .Q(n24[20]));
    not g995(n459 ,n10[30]);
    not g996(n2059 ,n2060);
    not g997(n118 ,n24[4]);
    dff g998(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1273), .Q(n10[7]));
    or g999(n1841 ,n681 ,n1784);
    nor g1000(n1759 ,n237 ,n1444);
    or g1001(n1987 ,n578 ,n1564);
    dff g1002(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1205), .Q(n14[1]));
    nor g1003(n1481 ,n468 ,n1370);
    nor g1004(n1057 ,n367 ,n106);
    buf g1005(n12[1], n10[1]);
    nor g1006(n889 ,n243 ,n99);
    nor g1007(n871 ,n134 ,n104);
    buf g1008(n12[2], n10[2]);
    or g1009(n628 ,n23[1] ,n525);
    or g1010(n1893 ,n1701 ,n1622);
    or g1011(n2045 ,n1553 ,n1981);
    nor g1012(n1462 ,n414 ,n1371);
    nor g1013(n77 ,n73 ,n70);
    nor g1014(n1348 ,n1325 ,n1343);
    not g1015(n342 ,n22[9]);
    or g1016(n2051 ,n1565 ,n1987);
    not g1017(n191 ,n28[2]);
    nor g1018(n67 ,n27[6] ,n65);
    nor g1019(n1376 ,n137 ,n1362);
    not g1020(n255 ,n5[27]);
    nor g1021(n80 ,n75 ,n78);
    nor g1022(n946 ,n174 ,n99);
    dff g1023(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1253), .Q(n12[21]));
    not g1024(n521 ,n18[1]);
    nor g1025(n984 ,n327 ,n101);
    not g1026(n307 ,n24[6]);
    not g1027(n314 ,n24[10]);
    nor g1028(n892 ,n136 ,n103);
    not g1029(n293 ,n23[2]);
    nor g1030(n994 ,n331 ,n101);
    dff g1031(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1918), .Q(n30[11]));
    buf g1032(n14[8], 1'b0);
    nor g1033(n1416 ,n388 ,n1368);
    dff g1034(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2075), .Q(n29[1]));
    nor g1035(n666 ,n97 ,n606);
    or g1036(n1924 ,n1732 ,n1638);
    not g1037(n228 ,n10[15]);
    not g1038(n327 ,n20[6]);
    nor g1039(n68 ,n45 ,n66);
    nor g1040(n1430 ,n258 ,n1370);
    not g1041(n427 ,n10[28]);
    or g1042(n1118 ,n281 ,n640);
    nor g1043(n1712 ,n417 ,n1440);
    nor g1044(n806 ,n505 ,n99);
    not g1045(n391 ,n30[18]);
    or g1046(n1962 ,n549 ,n1674);
    not g1047(n322 ,n19[1]);
    nor g1048(n550 ,n419 ,n3);
    nor g1049(n1651 ,n1115 ,n1445);
    or g1050(n1239 ,n918 ,n666);
    or g1051(n532 ,n4[23] ,n4[22]);
    dff g1052(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1213), .Q(n13[27]));
    nor g1053(n1617 ,n1116 ,n1443);
    nor g1054(n1822 ,n352 ,n1447);
    not g1055(n465 ,n9[2]);
    nor g1056(n756 ,n114 ,n96);
    or g1057(n1898 ,n1706 ,n1671);
    nor g1058(n83 ,n72 ,n81);
    dff g1059(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1295), .Q(n12[25]));
    nor g1060(n563 ,n465 ,n3);
    or g1061(n1972 ,n576 ,n1534);
    or g1062(n1369 ,n107 ,n1365);
    or g1063(n1312 ,n846 ,n787);
    nor g1064(n807 ,n340 ,n103);
    or g1065(n1122 ,n811 ,n782);
    dff g1066(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1895), .Q(n22[2]));
    nor g1067(n1083 ,n156 ,n106);
    or g1068(n1238 ,n916 ,n665);
    not g1069(n396 ,n12[27]);
    not g1070(n288 ,n2066);
    nor g1071(n1374 ,n137 ,n1364);
    nor g1072(n827 ,n320 ,n103);
    or g1073(n2111 ,n2099 ,n2097);
    dff g1074(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1893), .Q(n22[4]));
    nor g1075(n1786 ,n239 ,n1446);
    buf g1076(n17[0], n14[4]);
    not g1077(n155 ,n22[31]);
    dff g1078(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2040), .Q(n9[10]));
    or g1079(n877 ,n233 ,n640);
    nor g1080(n61 ,n27[4] ,n59);
    nor g1081(n1451 ,n142 ,n1369);
    xnor g1082(n616 ,n20[4] ,n24[4]);
    nor g1083(n856 ,n97 ,n604);
    nor g1084(n1789 ,n154 ,n1447);
    dff g1085(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1223), .Q(n13[18]));
    nor g1086(n1795 ,n350 ,n1447);
    or g1087(n1228 ,n893 ,n659);
    dff g1088(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2008), .Q(n25[17]));
    or g1089(n2009 ,n1802 ,n1849);
    nor g1090(n1044 ,n146 ,n106);
    not g1091(n512 ,n13[26]);
    nor g1092(n840 ,n335 ,n104);
    or g1093(n1520 ,n1388 ,n1389);
    or g1094(n1165 ,n723 ,n1047);
    not g1095(n156 ,n22[27]);
    or g1096(n1207 ,n859 ,n1069);
    nor g1097(n1090 ,n290 ,n638);
    nor g1098(n1588 ,n879 ,n1441);
    or g1099(n1234 ,n906 ,n662);
    buf g1100(n14[23], n10[19]);
    or g1101(n2101 ,n2082 ,n24[17]);
    not g1102(n266 ,n27[4]);
    dff g1103(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2010), .Q(n25[15]));
    nor g1104(n826 ,n230 ,n98);
    or g1105(n1224 ,n892 ,n1075);
    nor g1106(n1780 ,n364 ,n1447);
    nor g1107(n793 ,n130 ,n104);
    nor g1108(n584 ,n406 ,n3);
    not g1109(n257 ,n30[19]);
    xnor g1110(n597 ,n20[30] ,n24[30]);
    dff g1111(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2032), .Q(n9[18]));
    nor g1112(n1736 ,n397 ,n1440);
    not g1113(n340 ,n20[24]);
    dff g1114(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1283), .Q(n10[30]));
    or g1115(n1289 ,n957 ,n1000);
    or g1116(n1107 ,n186 ,n640);
    not g1117(n467 ,n9[5]);
    nor g1118(n1791 ,n162 ,n1447);
    not g1119(n638 ,n639);
    or g1120(n1366 ,n1319 ,n1361);
    nor g1121(n711 ,n628 ,n629);
    nor g1122(n1675 ,n382 ,n1442);
    dff g1123(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1257), .Q(n15[6]));
    dff g1124(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1276), .Q(n10[11]));
    xnor g1125(n651 ,n294 ,n19[1]);
    or g1126(n1909 ,n1717 ,n1581);
    or g1127(n2033 ,n1529 ,n1969);
    nor g1128(n656 ,n97 ,n605);
    nor g1129(n2073 ,n82 ,n83);
    or g1130(n2090 ,n24[31] ,n24[30]);
    nor g1131(n1474 ,n191 ,n1370);
    or g1132(n2096 ,n24[9] ,n24[8]);
    dff g1133(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2046), .Q(n9[4]));
    nor g1134(n1763 ,n217 ,n1444);
    or g1135(n646 ,n547 ,n526);
    not g1136(n129 ,n4[3]);
    nor g1137(n1445 ,n640 ,n1376);
    nor g1138(n1021 ,n369 ,n106);
    or g1139(n1347 ,n625 ,n93);
    nor g1140(n1747 ,n261 ,n1444);
    or g1141(n1217 ,n813 ,n656);
    dff g1142(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1915), .Q(n30[15]));
    or g1143(n2001 ,n1785 ,n1841);
    dff g1144(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1158), .Q(n20[25]));
    dff g1145(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1285), .Q(n10[4]));
    nor g1146(n1063 ,n206 ,n105);
    or g1147(n525 ,n23[0] ,n23[2]);
    nor g1148(n1095 ,n285 ,n638);
    or g1149(n1941 ,n1749 ,n1586);
    or g1150(n1310 ,n971 ,n766);
    nor g1151(n1082 ,n150 ,n105);
    not g1152(n483 ,n11[2]);
    nor g1153(n1774 ,n144 ,n1447);
    or g1154(n1142 ,n744 ,n1073);
    or g1155(n1882 ,n1690 ,n1611);
    nor g1156(n1788 ,n212 ,n1446);
    not g1157(n75 ,n29[2]);
    dff g1158(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1948), .Q(n28[13]));
    nor g1159(n836 ,n97 ,n618);
    nor g1160(n1635 ,n1110 ,n1441);
    not g1161(n318 ,n20[27]);
    dff g1162(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1904), .Q(n30[25]));
    or g1163(n527 ,n8[3] ,n8[2]);
    or g1164(n864 ,n644 ,n641);
    or g1165(n1973 ,n587 ,n1536);
    or g1166(n1930 ,n1738 ,n1580);
    nor g1167(n1470 ,n515 ,n1371);
    nor g1168(n1420 ,n161 ,n1369);
    not g1169(n399 ,n30[21]);
    or g1170(n1957 ,n1765 ,n1666);
    or g1171(n1447 ,n554 ,n1372);
    not g1172(n107 ,n3);
    nor g1173(n799 ,n252 ,n99);
    not g1174(n198 ,n5[28]);
    not g1175(n183 ,n5[17]);
    nor g1176(n1014 ,n338 ,n101);
    dff g1177(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1225), .Q(n13[1]));
    nor g1178(n1606 ,n876 ,n1443);
    nor g1179(n700 ,n638 ,n622);
    or g1180(n1114 ,n184 ,n640);
    nor g1181(n663 ,n97 ,n619);
    nor g1182(n1594 ,n884 ,n1443);
    nor g1183(n1805 ,n388 ,n1447);
    not g1184(n420 ,n30[20]);
    or g1185(n1152 ,n746 ,n1031);
    nor g1186(n845 ,n319 ,n103);
    not g1187(n78 ,n77);
    not g1188(n341 ,n15[3]);
    or g1189(n524 ,n6[1] ,n6[0]);
    or g1190(n1244 ,n942 ,n777);
    not g1191(n416 ,n28[4]);
    or g1192(n1350 ,n1329 ,n1340);
    nor g1193(n937 ,n395 ,n98);
    or g1194(n1123 ,n934 ,n977);
    not g1195(n388 ,n25[14]);
    or g1196(n1551 ,n1456 ,n1455);
    not g1197(n2077 ,n24[4]);
    nor g1198(n749 ,n309 ,n104);
    nor g1199(n833 ,n460 ,n102);
    nor g1200(n578 ,n269 ,n3);
    or g1201(n2039 ,n1541 ,n1975);
    nor g1202(n732 ,n300 ,n104);
    nor g1203(n772 ,n313 ,n101);
    nor g1204(n1443 ,n640 ,n1375);
    nor g1205(n861 ,n489 ,n639);
    not g1206(n215 ,n9[6]);
    or g1207(n1311 ,n818 ,n759);
    dff g1208(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2028), .Q(n9[22]));
    not g1209(n171 ,n5[20]);
    or g1210(n546 ,n6[3] ,n6[2]);
    or g1211(n2042 ,n1547 ,n1978);
    nor g1212(n872 ,n464 ,n99);
    not g1213(n285 ,n2067);
    nor g1214(n781 ,n302 ,n101);
    dff g1215(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2003), .Q(n25[22]));
    nor g1216(n865 ,n509 ,n99);
    nor g1217(n739 ,n298 ,n103);
    nor g1218(n925 ,n440 ,n99);
    nor g1219(n1020 ,n382 ,n105);
    or g1220(n1943 ,n1751 ,n1653);
    not g1221(n297 ,n26[0]);
    or g1222(n1938 ,n1746 ,n1648);
    nor g1223(n1465 ,n356 ,n1369);
    nor g1224(n1072 ,n357 ,n106);
    or g1225(n1377 ,n1353 ,n1367);
    dff g1226(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1304), .Q(n10[17]));
    not g1227(n329 ,n20[5]);
    nor g1228(n1781 ,n380 ,n1447);
    nor g1229(n660 ,n97 ,n609);
    nor g1230(n1502 ,n203 ,n1370);
    dff g1231(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1130), .Q(n13[0]));
    not g1232(n349 ,n25[1]);
    dff g1233(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1955), .Q(n28[6]));
    nor g1234(n678 ,n97 ,n653);
    nor g1235(n1434 ,n445 ,n1371);
    or g1236(n1968 ,n568 ,n1526);
    nor g1237(n1399 ,n257 ,n1371);
    nor g1238(n1739 ,n392 ,n1444);
    not g1239(n2087 ,n24[27]);
    nor g1240(n1450 ,n408 ,n1371);
    not g1241(n45 ,n27[6]);
    nor g1242(n1408 ,n358 ,n1369);
    nor g1243(n997 ,n165 ,n96);
    or g1244(n2011 ,n1805 ,n1851);
    nor g1245(n1463 ,n368 ,n1368);
    or g1246(n528 ,n8[5] ,n8[4]);
    nor g1247(n1626 ,n1104 ,n1443);
    not g1248(n515 ,n30[3]);
    not g1249(n315 ,n24[16]);
    or g1250(n1277 ,n837 ,n993);
    dff g1251(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1132), .Q(n11[3]));
    nor g1252(n657 ,n97 ,n607);
    nor g1253(n1435 ,n237 ,n1370);
    or g1254(n41 ,n27[1] ,n39);
    buf g1255(n14[16], n10[12]);
    dff g1256(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1922), .Q(n30[7]));
    nor g1257(n1505 ,n377 ,n1369);
    nor g1258(n894 ,n507 ,n98);
    buf g1259(n14[25], n10[21]);
    not g1260(n474 ,n9[26]);
    nor g1261(n738 ,n113 ,n104);
    or g1262(n1214 ,n917 ,n830);
    nor g1263(n1607 ,n875 ,n1443);
    or g1264(n1308 ,n972 ,n1089);
    or g1265(n1170 ,n793 ,n1048);
    dff g1266(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2024), .Q(n25[1]));
    nor g1267(n981 ,n329 ,n101);
    nor g1268(n536 ,n443 ,n3);
    not g1269(n195 ,n11[15]);
    nor g1270(n942 ,n496 ,n99);
    nor g1271(n1625 ,n1103 ,n1443);
    nor g1272(n698 ,n638 ,n609);
    nor g1273(n1431 ,n439 ,n1371);
    not g1274(n344 ,n25[25]);
    dff g1275(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1210), .Q(n20[8]));
    nor g1276(n936 ,n123 ,n104);
    not g1277(n330 ,n21[0]);
    not g1278(n500 ,n30[0]);
    dff g1279(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1200), .Q(n19[0]));
    dff g1280(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1921), .Q(n30[8]));
    not g1281(n69 ,n29[6]);
    nor g1282(n1001 ,n336 ,n96);
    dff g1283(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1936), .Q(n28[25]));
    or g1284(n2024 ,n1831 ,n1872);
    nor g1285(n1429 ,n159 ,n1369);
    dff g1286(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1952), .Q(n28[9]));
    nor g1287(n1509 ,n344 ,n1368);
    dff g1288(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1169), .Q(n24[8]));
    not g1289(n385 ,n22[2]);
    or g1290(n1575 ,n1506 ,n1507);
    not g1291(n553 ,n554);
    dff g1292(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1180), .Q(n24[5]));
    dff g1293(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1209), .Q(n13[30]));
    not g1294(n264 ,n10[9]);
    buf g1295(n17[13], n10[5]);
    dff g1296(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1900), .Q(n30[29]));
    not g1297(n520 ,n12[24]);
    nor g1298(n579 ,n268 ,n3);
    dff g1299(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1232), .Q(n13[13]));
    not g1300(n213 ,n5[14]);
    nor g1301(n1802 ,n386 ,n1447);
    or g1302(n1518 ,n1387 ,n1386);
    xnor g1303(n602 ,n20[31] ,n24[31]);
    or g1304(n2110 ,n2100 ,n2104);
    or g1305(n1913 ,n1723 ,n1631);
    not g1306(n208 ,n10[17]);
    nor g1307(n1042 ,n160 ,n106);
    dff g1308(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1211), .Q(n13[29]));
    dff g1309(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2052), .Q(n9[30]));
    buf g1310(n17[6], 1'b0);
    or g1311(n2034 ,n1531 ,n1970);
    nor g1312(n777 ,n305 ,n101);
    or g1313(n1863 ,n704 ,n1820);
    nor g1314(n1086 ,n389 ,n105);
    not g1315(n421 ,n9[30]);
    dff g1316(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1226), .Q(n13[17]));
    or g1317(n2050 ,n1563 ,n1986);
    or g1318(n1862 ,n1677 ,n1597);
    or g1319(n1916 ,n1724 ,n1654);
    or g1320(n1871 ,n1681 ,n1601);
    or g1321(n1904 ,n1712 ,n1590);
    not g1322(n440 ,n13[3]);
    not g1323(n378 ,n22[10]);
    dff g1324(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1183), .Q(n20[18]));
    nor g1325(n1013 ,n126 ,n101);
    not g1326(n497 ,n28[28]);
    or g1327(n1193 ,n833 ,n755);
    nor g1328(n1016 ,n333 ,n96);
    nor g1329(n911 ,n190 ,n99);
    or g1330(n1188 ,n838 ,n1064);
    nor g1331(n812 ,n317 ,n103);
    nor g1332(n959 ,n492 ,n102);
    nor g1333(n944 ,n458 ,n99);
    or g1334(n1285 ,n834 ,n1018);
    dff g1335(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1889), .Q(n22[8]));
    nor g1336(n1150 ,n641 ,n790);
    nor g1337(n1610 ,n1102 ,n1443);
    buf g1338(n17[8], n10[0]);
    dff g1339(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1121), .Q(n12[24]));
    dff g1340(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2049), .Q(n9[1]));
    dff g1341(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1937), .Q(n28[24]));
    nor g1342(n1715 ,n502 ,n1440);
    or g1343(n1220 ,n889 ,n657);
    nor g1344(n1394 ,n173 ,n1370);
    nor g1345(n1052 ,n384 ,n105);
    or g1346(n1212 ,n802 ,n839);
    not g1347(n238 ,n14[4]);
    nor g1348(n1833 ,n240 ,n1444);
    nor g1349(n1089 ,n216 ,n105);
    not g1350(n457 ,n10[23]);
    nor g1351(n740 ,n116 ,n103);
    not g1352(n243 ,n13[21]);
    dff g1353(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1957), .Q(n28[4]));
    not g1354(n321 ,n20[3]);
    buf g1355(n14[26], n10[22]);
    nor g1356(n1439 ,n157 ,n1368);
    nor g1357(n1097 ,n2059 ,n638);
    nor g1358(n1436 ,n342 ,n1369);
    or g1359(n1293 ,n941 ,n1011);
    dff g1360(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1288), .Q(n10[27]));
    nor g1361(n692 ,n638 ,n596);
    nor g1362(n893 ,n201 ,n99);
    or g1363(n632 ,n532 ,n538);
    nor g1364(n814 ,n325 ,n104);
    nor g1365(n1832 ,n367 ,n1447);
    or g1366(n1139 ,n747 ,n1021);
    not g1367(n221 ,n13[7]);
    nor g1368(n1629 ,n878 ,n1441);
    xnor g1369(n614 ,n20[8] ,n24[8]);
    nor g1370(n1655 ,n1105 ,n1445);
    nor g1371(n1479 ,n367 ,n1368);
    or g1372(n1517 ,n1383 ,n1382);
    or g1373(n1861 ,n703 ,n1818);
    dff g1374(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1177), .Q(n26[1]));
    or g1375(n2053 ,n1569 ,n1989);
    nor g1376(n1027 ,n151 ,n106);
    not g1377(n495 ,n30[31]);
    not g1378(n180 ,n10[8]);
    or g1379(n1906 ,n1714 ,n1588);
    dff g1380(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2020), .Q(n25[5]));
    dff g1381(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1170), .Q(n20[21]));
    nor g1382(n1741 ,n497 ,n1444);
    not g1383(n242 ,n5[19]);
    nor g1384(n673 ,n97 ,n596);
    not g1385(n222 ,n28[17]);
    or g1386(n1947 ,n1755 ,n1656);
    nor g1387(n714 ,n21[3] ,n593);
    nor g1388(n733 ,n112 ,n104);
    or g1389(n1880 ,n1687 ,n1609);
    not g1390(n517 ,n12[31]);
    nor g1391(n897 ,n278 ,n98);
    nor g1392(n1504 ,n380 ,n1368);
    nor g1393(n641 ,n293 ,n545);
    buf g1394(n14[19], n10[15]);
    nor g1395(n1077 ,n356 ,n105);
    or g1396(n2041 ,n1544 ,n1977);
    not g1397(n182 ,n13[17]);
    xnor g1398(n611 ,n20[15] ,n24[15]);
    not g1399(n466 ,n13[8]);
    nor g1400(n914 ,n466 ,n99);
    dff g1401(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1914), .Q(n30[16]));
    or g1402(n1221 ,n905 ,n1072);
    or g1403(n1926 ,n1733 ,n1635);
    dff g1404(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1997), .Q(n25[27]));
    xnor g1405(n593 ,n24[3] ,n321);
    or g1406(n20[1] ,n19[1] ,n2119);
    or g1407(n1098 ,n135 ,n645);
    dff g1408(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1888), .Q(n22[9]));
    or g1409(n1253 ,n932 ,n779);
    not g1410(n417 ,n30[25]);
    nor g1411(n1792 ,n346 ,n1447);
    not g1412(n300 ,n26[1]);
    nor g1413(n668 ,n96 ,n615);
    not g1414(n506 ,n12[29]);
    or g1415(n1295 ,n822 ,n763);
    nor g1416(n1705 ,n372 ,n1442);
    nor g1417(n2075 ,n77 ,n76);
    nor g1418(n1587 ,n877 ,n1445);
    or g1419(n2048 ,n1559 ,n1984);
    or g1420(n1124 ,n825 ,n784);
    nor g1421(n707 ,n638 ,n655);
    or g1422(n1932 ,n1740 ,n1643);
    or g1423(n2116 ,n2115 ,n2113);
    dff g1424(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1870), .Q(n22[25]));
    not g1425(n290 ,n2062);
    not g1426(n492 ,n10[11]);
    nor g1427(n908 ,n279 ,n98);
    dff g1428(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1929), .Q(n30[1]));
    or g1429(n1569 ,n1495 ,n1494);
    dff g1430(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1250), .Q(n10[0]));
    nor g1431(n1830 ,n187 ,n1446);
    or g1432(n1148 ,n749 ,n1028);
    or g1433(n1894 ,n1702 ,n1623);
    not g1434(n138 ,n22[12]);
    not g1435(n178 ,n5[30]);
    nor g1436(n1787 ,n153 ,n1447);
    dff g1437(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1135), .Q(n11[1]));
    buf g1438(n17[12], n10[4]);
    dff g1439(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2071), .Q(n29[5]));
    or g1440(n1866 ,n706 ,n1824);
    dff g1441(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1953), .Q(n28[8]));
    nor g1442(n697 ,n638 ,n611);
    not g1443(n452 ,n30[4]);
    dff g1444(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1240), .Q(n13[5]));
    or g1445(n1127 ,n820 ,n1063);
    or g1446(n1185 ,n819 ,n1056);
    nor g1447(n970 ,n224 ,n639);
    dff g1448(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2035), .Q(n9[15]));
    not g1449(n335 ,n21[2]);
    xnor g1450(n600 ,n26[0] ,n330);
    not g1451(n158 ,n15[4]);
    not g1452(n116 ,n24[21]);
    not g1453(n1341 ,n1150);
    nor g1454(n1697 ,n147 ,n1442);
    or g1455(n1536 ,n1420 ,n1421);
    buf g1456(n17[1], n14[5]);
    nor g1457(n1710 ,n487 ,n1440);
    nor g1458(n1382 ,n244 ,n1370);
    not g1459(n205 ,n18[0]);
    or g1460(n1884 ,n1692 ,n1613);
    nor g1461(n1771 ,n150 ,n1447);
    dff g1462(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1187), .Q(n11[6]));
    nor g1463(n702 ,n638 ,n614);
    xnor g1464(n598 ,n26[1] ,n331);
    not g1465(n489 ,n27[1]);
    nor g1466(n2071 ,n88 ,n89);
    nor g1467(n1395 ,n420 ,n1371);
    or g1468(n1899 ,n1703 ,n1625);
    nor g1469(n809 ,n338 ,n103);
    not g1470(n160 ,n25[13]);
    not g1471(n445 ,n30[10]);
    or g1472(n1864 ,n1678 ,n1598);
    or g1473(n1197 ,n844 ,n1065);
    not g1474(n499 ,n12[16]);
    nor g1475(n1811 ,n177 ,n1446);
    not g1476(n110 ,n8[0]);
    nor g1477(n727 ,n115 ,n103);
    or g1478(n1233 ,n904 ,n661);
    nor g1479(n1637 ,n1106 ,n1441);
    xnor g1480(n608 ,n20[20] ,n24[20]);
    or g1481(n2060 ,n27[6] ,n44);
    not g1482(n461 ,n10[27]);
    or g1483(n1208 ,n866 ,n851);
    not g1484(n501 ,n10[21]);
    nor g1485(n104 ,n295 ,n558);
    nor g1486(n758 ,n306 ,n96);
    nor g1487(n932 ,n275 ,n99);
    not g1488(n1442 ,n1443);
    nor g1489(n736 ,n307 ,n103);
    nor g1490(n1764 ,n231 ,n1444);
    or g1491(n526 ,n4[13] ,n4[12]);
    or g1492(n1562 ,n1513 ,n1479);
    dff g1493(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2037), .Q(n9[13]));
    or g1494(n33 ,n29[3] ,n29[2]);
    nor g1495(n843 ,n97 ,n603);
    nor g1496(n1472 ,n385 ,n1369);
    nor g1497(n1048 ,n343 ,n105);
    not g1498(n413 ,n13[6]);
    nor g1499(n926 ,n503 ,n99);
    not g1500(n283 ,n10[16]);
    nor g1501(n1401 ,n384 ,n1369);
    nor g1502(n1812 ,n166 ,n1447);
    buf g1503(n14[31], n10[27]);
    not g1504(n2082 ,n24[16]);
    nor g1505(n1427 ,n235 ,n1371);
    not g1506(n259 ,n9[15]);
    buf g1507(n12[15], n10[15]);
    or g1508(n1225 ,n841 ,n853);
    or g1509(n1335 ,n987 ,n1262);
    or g1510(n1120 ,n791 ,n770);
    nor g1511(n629 ,n546 ,n524);
    nor g1512(n1600 ,n881 ,n1443);
    not g1513(n504 ,n9[22]);
    or g1514(n1355 ,n627 ,n93);
    or g1515(n1942 ,n1750 ,n1652);
    nor g1516(n1699 ,n351 ,n1442);
    or g1517(n1982 ,n562 ,n1556);
    nor g1518(n1404 ,n365 ,n1369);
    not g1519(n262 ,n30[24]);
    or g1520(n1103 ,n247 ,n640);
    nor g1521(n1410 ,n430 ,n1370);
    or g1522(n1967 ,n584 ,n1524);
    nor g1523(n1590 ,n881 ,n1441);
    nor g1524(n1498 ,n497 ,n1370);
    nor g1525(n1494 ,n181 ,n1370);
    not g1526(n488 ,n9[14]);
    or g1527(n1351 ,n1327 ,n1341);
    not g1528(n84 ,n83);
    dff g1529(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1206), .Q(n14[0]));
    or g1530(n1878 ,n1686 ,n1607);
    not g1531(n439 ,n30[11]);
    nor g1532(n1608 ,n874 ,n1443);
    dff g1533(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1932), .Q(n28[29]));
    dff g1534(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1191), .Q(n11[14]));
    not g1535(n131 ,n20[8]);
    or g1536(n2023 ,n1829 ,n1869);
    not g1537(n496 ,n12[20]);
    nor g1538(n866 ,n428 ,n98);
    dff g1539(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1155), .Q(n20[24]));
    dff g1540(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1238), .Q(n13[7]));
    not g1541(n429 ,n13[11]);
    dff g1542(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1181), .Q(n24[4]));
    not g1543(n250 ,n11[1]);
    nor g1544(n991 ,n319 ,n96);
    nor g1545(n763 ,n310 ,n101);
    nor g1546(n1653 ,n874 ,n1445);
    not g1547(n187 ,n5[1]);
    xnor g1548(n591 ,n24[2] ,n323);
    nor g1549(n1579 ,n1102 ,n1445);
    nor g1550(n1716 ,n399 ,n1440);
    nor g1551(n941 ,n457 ,n102);
    or g1552(n2098 ,n2078 ,n24[2]);
    nor g1553(n1760 ,n404 ,n1444);
    or g1554(n1201 ,n845 ,n1067);
    xnor g1555(n607 ,n20[21] ,n24[21]);
    buf g1556(n11[19], n10[19]);
    or g1557(n1559 ,n1473 ,n1474);
    dff g1558(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2048), .Q(n9[2]));
    not g1559(n189 ,n5[12]);
    nor g1560(n980 ,n131 ,n101);
    or g1561(n1230 ,n894 ,n675);
    nor g1562(n1352 ,n645 ,n1345);
    nor g1563(n1437 ,n390 ,n1368);
    nor g1564(n773 ,n297 ,n96);
    or g1565(n1981 ,n588 ,n1552);
    dff g1566(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1995), .Q(n25[30]));
    nor g1567(n1513 ,n374 ,n1369);
    or g1568(n1574 ,n1505 ,n1504);
    dff g1569(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1174), .Q(n27[2]));
    or g1570(n1992 ,n548 ,n1574);
    nor g1571(n1055 ,n192 ,n106);
    dff g1572(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2029), .Q(n9[20]));
    dff g1573(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1126), .Q(n12[28]));
    nor g1574(n1748 ,n282 ,n1444);
    buf g1575(n14[9], 1'b0);
    or g1576(n1144 ,n742 ,n1025);
    nor g1577(n859 ,n125 ,n103);
    or g1578(n882 ,n255 ,n640);
    buf g1579(n11[20], n10[20]);
    or g1580(n1911 ,n1719 ,n1630);
    not g1581(n468 ,n28[0]);
    not g1582(n249 ,n28[25]);
    or g1583(n1919 ,n1727 ,n1632);
    dff g1584(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1951), .Q(n28[10]));
    or g1585(n1100 ,n198 ,n640);
    not g1586(n246 ,n11[10]);
    dff g1587(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2034), .Q(n9[16]));
    xor g1588(n2062 ,n27[7] ,n68);
    dff g1589(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2017), .Q(n25[8]));
    nor g1590(n1740 ,n181 ,n1444);
    not g1591(n463 ,n30[13]);
    dff g1592(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1268), .Q(n10[15]));
    not g1593(n317 ,n20[19]);
    nor g1594(n1075 ,n145 ,n106);
    or g1595(n1363 ,n94 ,n1355);
    xnor g1596(n654 ,n20[18] ,n24[18]);
    nor g1597(n2063 ,n67 ,n68);
    dff g1598(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1935), .Q(n28[27]));
    or g1599(n1953 ,n1761 ,n1651);
    or g1600(n1181 ,n730 ,n1051);
    not g1601(n177 ,n5[10]);
    or g1602(n1925 ,n1737 ,n1640);
    nor g1603(n1396 ,n350 ,n1368);
    nor g1604(n1668 ,n1106 ,n1445);
    or g1605(n2003 ,n1789 ,n1843);
    nor g1606(n1797 ,n141 ,n1447);
    or g1607(n1112 ,n211 ,n640);
    nor g1608(n852 ,n410 ,n99);
    dff g1609(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1156), .Q(n24[17]));
    nor g1610(n1484 ,n155 ,n1369);
    dff g1611(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1896), .Q(n22[1]));
    not g1612(n102 ,n101);
    nor g1613(n1682 ,n362 ,n1442);
    not g1614(n592 ,n591);
    nor g1615(n903 ,n411 ,n99);
    not g1616(n275 ,n12[21]);
    not g1617(n411 ,n12[30]);
    not g1618(n179 ,n13[28]);
    nor g1619(n713 ,n21[2] ,n591);
    buf g1620(n17[4], 1'b0);
    not g1621(n194 ,n5[31]);
    or g1622(n1848 ,n687 ,n1798);
    nor g1623(n1801 ,n277 ,n1446);
    nor g1624(n1499 ,n447 ,n1371);
    or g1625(n1990 ,n573 ,n1570);
    xnor g1626(n613 ,n20[9] ,n24[9]);
    or g1627(n880 ,n272 ,n640);
    or g1628(n1278 ,n821 ,n982);
    xnor g1629(n609 ,n20[14] ,n24[14]);
    or g1630(n1555 ,n1467 ,n1466);
    dff g1631(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1215), .Q(n13[25]));
    nor g1632(n644 ,n23[2] ,n556);
    not g1633(n455 ,n13[13]);
    not g1634(n154 ,n25[22]);
    dff g1635(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2018), .Q(n25[7]));
    dff g1636(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1197), .Q(n20[12]));
    dff g1637(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1172), .Q(n24[7]));
    nor g1638(n42 ,n40 ,n41);
    nor g1639(n567 ,n423 ,n3);
    or g1640(n1290 ,n953 ,n1010);
    or g1641(n1843 ,n692 ,n1788);
    nor g1642(n1627 ,n884 ,n1441);
    nor g1643(n1005 ,n337 ,n96);
    not g1644(n210 ,n8[3]);
    nor g1645(n1500 ,n364 ,n1368);
    dff g1646(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1883), .Q(n22[14]));
    nor g1647(n800 ,n132 ,n103);
    nor g1648(n1074 ,n351 ,n106);
    nor g1649(n696 ,n638 ,n654);
    dff g1650(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1280), .Q(n10[8]));
    nor g1651(n551 ,n453 ,n3);
    dff g1652(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1144), .Q(n24[26]));
    not g1653(n453 ,n9[0]);
    nor g1654(n757 ,n298 ,n101);
    or g1655(n1865 ,n705 ,n1822);
    not g1656(n282 ,n28[21]);
    not g1657(n419 ,n9[20]);
    buf g1658(n11[31], n10[31]);
    or g1659(n715 ,n630 ,n633);
    nor g1660(n786 ,n112 ,n96);
    or g1661(n2035 ,n1533 ,n1971);
    nor g1662(n570 ,n398 ,n3);
    nor g1663(n1388 ,n343 ,n1369);
    nor g1664(n1071 ,n142 ,n106);
    dff g1665(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2055), .Q(n9[27]));
    nor g1666(n1732 ,n414 ,n1440);
    buf g1667(n11[22], n10[22]);
    nor g1668(n575 ,n469 ,n3);
    nor g1669(n1615 ,n1109 ,n1443);
    xnor g1670(n655 ,n20[16] ,n24[16]);
    nor g1671(n1611 ,n1105 ,n1443);
    or g1672(n1200 ,n913 ,n1079);
    not g1673(n185 ,n5[18]);
    nor g1674(n969 ,n195 ,n102);
    or g1675(n1563 ,n1482 ,n1481);
    or g1676(n1516 ,n1380 ,n1381);
    or g1677(n1846 ,n695 ,n1794);
    dff g1678(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2016), .Q(n25[9]));
    nor g1679(n1743 ,n462 ,n1444);
    nor g1680(n1073 ,n364 ,n106);
    nor g1681(n1701 ,n145 ,n1442);
    buf g1682(n12[12], n10[12]);
    or g1683(n1128 ,n815 ,n756);
    nor g1684(n930 ,n481 ,n102);
    dff g1685(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1999), .Q(n25[26]));
    not g1686(n199 ,n30[23]);
    not g1687(n367 ,n25[0]);
    nor g1688(n689 ,n638 ,n595);
    nor g1689(n1490 ,n392 ,n1370);
    dff g1690(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1277), .Q(n10[10]));
    dff g1691(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1274), .Q(n10[12]));
    or g1692(n1177 ,n732 ,n1050);
    dff g1693(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1229), .Q(n20[3]));
    dff g1694(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1928), .Q(n30[2]));
    nor g1695(n1704 ,n385 ,n1442);
    nor g1696(n1512 ,n417 ,n1371);
    nor g1697(n1328 ,n370 ,n1324);
    nor g1698(n1349 ,n645 ,n1344);
    nor g1699(n1088 ,n360 ,n106);
    dff g1700(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1154), .Q(n24[18]));
    not g1701(n233 ,n5[21]);
    dff g1702(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2025), .Q(n9[25]));
    dff g1703(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1287), .Q(n10[3]));
    nor g1704(n987 ,n375 ,n101);
    nor g1705(n1036 ,n347 ,n106);
    or g1706(n571 ,n127 ,n4[3]);
    not g1707(n2088 ,n24[25]);
    dff g1708(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1218), .Q(n13[23]));
    nor g1709(n899 ,n371 ,n643);
    nor g1710(n1041 ,n352 ,n105);
    xnor g1711(n610 ,n20[17] ,n24[17]);
    not g1712(n114 ,n24[5]);
    dff g1713(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1886), .Q(n22[11]));
    nor g1714(n1029 ,n154 ,n106);
    not g1715(n302 ,n24[26]);
    nor g1716(n982 ,n125 ,n101);
    or g1717(n1997 ,n1780 ,n1838);
    or g1718(n1291 ,n751 ,n1026);
    or g1719(n2047 ,n1557 ,n1982);
    dff g1720(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1272), .Q(n20[5]));
    buf g1721(n11[30], n10[30]);
    or g1722(n545 ,n295 ,n23[1]);
    nor g1723(n1656 ,n1108 ,n1445);
    nor g1724(n965 ,n441 ,n102);
    or g1725(n1169 ,n754 ,n1088);
    dff g1726(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1880), .Q(n22[17]));
    nor g1727(n1698 ,n142 ,n1442);
    nor g1728(n935 ,n449 ,n99);
    or g1729(n1568 ,n1492 ,n1493);
    nor g1730(n1662 ,n1109 ,n1445);
    not g1731(n235 ,n30[12]);
    dff g1732(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1282), .Q(n10[5]));
    nor g1733(n1466 ,n416 ,n1370);
    not g1734(n376 ,n22[24]);
    not g1735(n145 ,n22[4]);
    nor g1736(n924 ,n435 ,n98);
    or g1737(n1940 ,n1748 ,n1587);
    not g1738(n240 ,n28[15]);
    or g1739(n1179 ,n729 ,n1046);
    dff g1740(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1163), .Q(n24[12]));
    nor g1741(n820 ,n331 ,n103);
    buf g1742(n14[11], 1'b0);
    nor g1743(n1460 ,n352 ,n1368);
    not g1744(n123 ,n20[30]);
    or g1745(n1573 ,n1503 ,n1502);
    or g1746(n1106 ,n214 ,n640);
    nor g1747(n1772 ,n369 ,n1447);
    nor g1748(n1336 ,n857 ,n1316);
    nor g1749(n573 ,n412 ,n3);
    or g1750(n1323 ,n810 ,n776);
    dff g1751(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1296), .Q(n10[22]));
    dff g1752(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1924), .Q(n30[5]));
    not g1753(n175 ,n28[7]);
    not g1754(n207 ,n5[4]);
    not g1755(n57 ,n56);
    nor g1756(n557 ,n23[1] ,n23[2]);
    nor g1757(n1353 ,n97 ,n1333);
    dff g1758(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1241), .Q(n20[2]));
    nor g1759(n554 ,n109 ,n23[0]);
    nor g1760(n745 ,n299 ,n103);
    nor g1761(n802 ,n179 ,n99);
    or g1762(n537 ,n4[19] ,n4[18]);
    nor g1763(n886 ,n424 ,n98);
    dff g1764(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1245), .Q(n10[20]));
    dff g1765(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1255), .Q(n19[1]));
    or g1766(n1571 ,n1499 ,n1498);
    or g1767(n2103 ,n2086 ,n2085);
    dff g1768(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1310), .Q(n11[13]));
    dff g1769(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1917), .Q(n30[12]));
    or g1770(n37 ,n29[7] ,n36);
    not g1771(n422 ,n9[25]);
    not g1772(n143 ,n25[2]);
    dff g1773(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1188), .Q(n20[14]));
    nor g1774(n1023 ,n139 ,n106);
    nor g1775(n1726 ,n439 ,n1440);
    not g1776(n441 ,n10[0]);
    dff g1777(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1185), .Q(n20[17]));
    nor g1778(n891 ,n373 ,n643);
    or g1779(n1111 ,n225 ,n640);
    nor g1780(n2074 ,n79 ,n80);
    buf g1781(n14[24], n10[20]);
    or g1782(n1549 ,n1454 ,n1453);
    nor g1783(n1622 ,n1110 ,n1443);
    buf g1784(n14[15], n10[11]);
    dff g1785(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1301), .Q(n10[18]));
    or g1786(n1989 ,n575 ,n1568);
    dff g1787(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1249), .Q(n12[22]));
    or g1788(n1168 ,n738 ,n1049);
    dff g1789(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1941), .Q(n28[20]));
    not g1790(n350 ,n25[19]);
    or g1791(n1326 ,n715 ,n718);
    or g1792(n1860 ,n1676 ,n1595);
    nor g1793(n928 ,n337 ,n103);
    dff g1794(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2072), .Q(n29[4]));
    not g1795(n375 ,n16[3]);
    dff g1796(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1949), .Q(n28[11]));
    nor g1797(n1820 ,n152 ,n1447);
    or g1798(n1187 ,n795 ,n764);
    not g1799(n147 ,n22[8]);
    not g1800(n112 ,n24[14]);
    nor g1801(n1385 ,n363 ,n1369);
    nor g1802(n955 ,n124 ,n104);
    dff g1803(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1958), .Q(n28[3]));
    nor g1804(n1750 ,n446 ,n1444);
    buf g1805(n12[7], n10[7]);
    nor g1806(n958 ,n256 ,n102);
    nor g1807(n1333 ,n530 ,n1322);
    not g1808(n402 ,n11[6]);
    dff g1809(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1927), .Q(n30[3]));
    nor g1810(n1432 ,n354 ,n1368);
    nor g1811(n811 ,n442 ,n99);
    not g1812(n556 ,n555);
    or g1813(n2108 ,n2094 ,n2102);
    nor g1814(n962 ,n461 ,n102);
    nor g1815(n1807 ,n160 ,n1447);
    or g1816(n2044 ,n1550 ,n1980);
    or g1817(n2097 ,n2083 ,n24[20]);
    dff g1818(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1278), .Q(n10[9]));
    or g1819(n1115 ,n193 ,n640);
    nor g1820(n960 ,n520 ,n102);
    buf g1821(n18[10], 1'b0);
    buf g1822(n14[2], 1'b0);
    or g1823(n1210 ,n863 ,n1070);
    not g1824(n491 ,n13[4]);
    not g1825(n432 ,n28[14]);
    dff g1826(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1236), .Q(n13[9]));
    dff g1827(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1264), .Q(n12[16]));
    nor g1828(n1672 ,n881 ,n1445);
    dff g1829(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1878), .Q(n22[19]));
    or g1830(n1359 ,n867 ,n1349);
    or g1831(n1538 ,n1425 ,n1424);
    nor g1832(n580 ,n493 ,n3);
    nor g1833(n1677 ,n387 ,n1442);
    or g1834(n1272 ,n895 ,n1074);
    dff g1835(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1899), .Q(n22[0]));
    nor g1836(n951 ,n518 ,n99);
    nor g1837(n887 ,n248 ,n99);
    or g1838(n1855 ,n1514 ,n1593);
    not g1839(n164 ,n20[0]);
    nor g1840(n1514 ,n155 ,n1442);
    dff g1841(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1925), .Q(n30[0]));
    dff g1842(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1998), .Q(n25[28]));
    not g1843(n510 ,n13[0]);
    nor g1844(n1737 ,n500 ,n1440);
    nor g1845(n853 ,n97 ,n635);
    not g1846(n446 ,n28[19]);
    nor g1847(n1024 ,n387 ,n105);
    nor g1848(n1722 ,n273 ,n1440);
    not g1849(n71 ,n29[4]);
    or g1850(n870 ,n641 ,n639);
    not g1851(n365 ,n22[17]);
    nor g1852(n1768 ,n498 ,n1444);
    nor g1853(n1423 ,n463 ,n1371);
    nor g1854(n842 ,n345 ,n643);
    or g1855(n1166 ,n796 ,n1032);
    not g1856(n458 ,n10[20]);
    dff g1857(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2051), .Q(n9[31]));
    dff g1858(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1351), .Q(n16[0]));
    or g1859(n1266 ,n641 ,n974);
    or g1860(n883 ,n169 ,n640);
    nor g1861(n862 ,n486 ,n99);
    dff g1862(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1894), .Q(n22[3]));
    nor g1863(n1669 ,n1104 ,n1445);
    not g1864(n244 ,n28[23]);
    nor g1865(n1720 ,n263 ,n1440);
    not g1866(n339 ,n19[0]);
    nor g1867(n988 ,n324 ,n101);
    nor g1868(n562 ,n438 ,n3);
    nor g1869(n1623 ,n1107 ,n1443);
    not g1870(n347 ,n22[19]);
    not g1871(n159 ,n22[11]);
    not g1872(n2076 ,n24[5]);
    nor g1873(n1591 ,n880 ,n1445);
    nor g1874(n1628 ,n1101 ,n1441);
    nor g1875(n1657 ,n1118 ,n1445);
    nor g1876(n35 ,n33 ,n32);
    not g1877(n153 ,n25[23]);
    or g1878(n1237 ,n914 ,n664);
    dff g1879(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1233), .Q(n13[12]));
    nor g1880(n737 ,n111 ,n104);
    dff g1881(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1943), .Q(n28[18]));
    or g1882(n1570 ,n1497 ,n1496);
    nor g1883(n979 ,n124 ,n101);
    or g1884(n627 ,n535 ,n95);
    nor g1885(n1485 ,n150 ,n1368);
    or g1886(n1890 ,n1698 ,n1619);
    not g1887(n286 ,n7[0]);
    not g1888(n130 ,n20[21]);
    buf g1889(n12[9], n10[9]);
    or g1890(n1222 ,n886 ,n658);
    dff g1891(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1160), .Q(n24[15]));
    or g1892(n1524 ,n1397 ,n1396);
    nor g1893(n705 ,n638 ,n615);
    nor g1894(n1636 ,n1107 ,n1441);
    or g1895(n1206 ,n865 ,n773);
    dff g1896(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1913), .Q(n30[14]));
    or g1897(n1219 ,n898 ,n673);
    dff g1898(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1923), .Q(n30[6]));
    nor g1899(n788 ,n297 ,n638);
    nor g1900(n921 ,n471 ,n99);
    nor g1901(n973 ,n479 ,n639);
    nor g1902(n858 ,n499 ,n98);
    nor g1903(n720 ,n108 ,n103);
    dff g1904(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1332), .Q(n15[1]));
    nor g1905(n1047 ,n354 ,n106);
    buf g1906(n14[13], n10[9]);
    nor g1907(n798 ,n451 ,n102);
    not g1908(n366 ,n15[1]);
    nor g1909(n76 ,n29[1] ,n29[0]);
    nor g1910(n1381 ,n153 ,n1368);
    nor g1911(n1066 ,n167 ,n105);
    or g1912(n1838 ,n683 ,n1778);
    not g1913(n358 ,n22[16]);
    nor g1914(n1469 ,n218 ,n1370);
    or g1915(n1525 ,n1399 ,n1398);
    not g1916(n173 ,n28[20]);
    nor g1917(n706 ,n638 ,n616);
    not g1918(n414 ,n30[5]);
    or g1919(n2027 ,n1517 ,n1963);
    or g1920(n1547 ,n1450 ,n1449);
    not g1921(n51 ,n27[2]);
    nor g1922(n1007 ,n340 ,n100);
    buf g1923(n11[25], n10[25]);
    or g1924(n1521 ,n1391 ,n1390);
    nor g1925(n1327 ,n383 ,n1324);
    dff g1926(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1898), .Q(n30[31]));
    dff g1927(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1947), .Q(n28[14]));
    nor g1928(n744 ,n311 ,n103);
    or g1929(n1566 ,n1489 ,n1488);
    not g1930(n448 ,n29[0]);
    nor g1931(n742 ,n302 ,n103);
    dff g1932(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1890), .Q(n22[7]));
    not g1933(n115 ,n24[3]);
    not g1934(n373 ,n15[6]);
    not g1935(n170 ,n28[13]);
    nor g1936(n1804 ,n213 ,n1446);
    nor g1937(n699 ,n638 ,n612);
    not g1938(n99 ,n101);
    nor g1939(n1621 ,n1111 ,n1443);
    nor g1940(n895 ,n329 ,n103);
    dff g1941(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1959), .Q(n28[2]));
    not g1942(n508 ,n14[7]);
    buf g1943(n12[3], n10[3]);
    or g1944(n1250 ,n965 ,n1002);
    nor g1945(n1631 ,n1108 ,n1441);
    nor g1946(n1507 ,n462 ,n1370);
    not g1947(n303 ,n24[24]);
    nor g1948(n1689 ,n358 ,n1442);
    nor g1949(n1666 ,n1110 ,n1445);
    nor g1950(n1706 ,n495 ,n1440);
    dff g1951(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1307), .Q(n10[16]));
    not g1952(n227 ,n28[18]);
    or g1953(n1264 ,n858 ,n767);
    not g1954(n357 ,n22[6]);
    dff g1955(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1145), .Q(n20[28]));
    nor g1956(n1486 ,n485 ,n1370);
    or g1957(n1354 ,n626 ,n93);
    nor g1958(n1059 ,n358 ,n105);
    not g1959(n599 ,n598);
    or g1960(n1174 ,n966 ,n1095);
    or g1961(n1958 ,n1766 ,n1667);
    not g1962(n46 ,n27[0]);
    or g1963(n710 ,n8[0] ,n634);
    buf g1964(n14[29], n10[25]);
    dff g1965(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2022), .Q(n25[3]));
    dff g1966(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1323), .Q(n18[0]));
    nor g1967(n1818 ,n140 ,n1447);
    dff g1968(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1161), .Q(n24[14]));
    or g1969(n1881 ,n1689 ,n1610);
    or g1970(n1334 ,n842 ,n1263);
    or g1971(n1368 ,n107 ,n1363);
    or g1972(n1141 ,n725 ,n1080);
    nor g1973(n1796 ,n185 ,n1446);
    buf g1974(n17[9], n10[1]);
    or g1975(n1889 ,n1697 ,n1618);
    nor g1976(n1428 ,n166 ,n1368);
    nor g1977(n1004 ,n128 ,n96);
    not g1978(n197 ,n5[9]);
    nor g1979(n1593 ,n885 ,n1443);
    not g1980(n165 ,n8[2]);
    nor g1981(n1815 ,n197 ,n1446);
    or g1982(n2017 ,n1817 ,n1859);
    not g1983(n74 ,n29[5]);
    buf g1984(n14[10], 1'b0);
    or g1985(n2020 ,n1823 ,n1865);
    nor g1986(n747 ,n120 ,n103);
    nor g1987(n1664 ,n1112 ,n1445);
    or g1988(n1540 ,n1429 ,n1428);
    dff g1989(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1357), .Q(n16[2]));
    nor g1990(n850 ,n335 ,n592);
    not g1991(n323 ,n20[2]);
    dff g1992(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1151), .Q(n24[21]));
    nor g1993(n898 ,n280 ,n98);
    nor g1994(n923 ,n133 ,n103);
    or g1995(n2029 ,n1523 ,n1966);
    or g1996(n547 ,n4[15] ,n4[14]);
    nor g1997(n1809 ,n146 ,n1447);
    dff g1998(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1259), .Q(n12[18]));
    nor g1999(n1619 ,n1114 ,n1443);
    nor g2000(n1598 ,n882 ,n1443);
    or g2001(n2106 ,n2103 ,n2092);
    nor g2002(n1793 ,n171 ,n1446);
    or g2003(n40 ,n27[2] ,n27[0]);
    or g2004(n1196 ,n903 ,n765);
    buf g2005(n14[28], n10[24]);
    dff g2006(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1217), .Q(n13[24]));
    not g2007(n400 ,n13[23]);
    or g2008(n1371 ,n107 ,n1364);
    dff g2009(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1148), .Q(n24[23]));
    nor g2010(n817 ,n229 ,n99);
    or g2011(n32 ,n29[1] ,n29[0]);
    not g2012(n49 ,n27[1]);
    not g2013(n359 ,n25[28]);
    or g2014(n2043 ,n1549 ,n1979);
    nor g2015(n1078 ,n372 ,n106);
    nor g2016(n779 ,n116 ,n101);
    nor g2017(n1828 ,n214 ,n1446);
    nor g2018(n1746 ,n244 ,n1444);
    nor g2019(n1758 ,n258 ,n1444);
    dff g2020(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1279), .Q(n10[2]));
    not g2021(n311 ,n24[27]);
    or g2022(n1995 ,n1773 ,n1835);
    dff g2023(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2031), .Q(n9[19]));
    or g2024(n2038 ,n1539 ,n1974);
    not g2025(n202 ,n28[12]);
    nor g2026(n694 ,n638 ,n608);
    or g2027(n1262 ,n641 ,n869);
    nor g2028(n1046 ,n286 ,n106);
    or g2029(n1532 ,n1412 ,n1413);
    nor g2030(n967 ,n444 ,n639);
    dff g2031(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1897), .Q(n30[30]));
    nor g2032(n586 ,n431 ,n3);
    nor g2033(n1776 ,n198 ,n1446);
    nor g2034(n1468 ,n348 ,n1368);
    nor g2035(n1049 ,n390 ,n105);
    nor g2036(n952 ,n407 ,n102);
    nor g2037(n746 ,n305 ,n103);
    nor g2038(n759 ,n301 ,n96);
    buf g2039(n14[30], n10[26]);
    nor g2040(n2067 ,n55 ,n56);
    nor g2041(n676 ,n97 ,n621);
    not g2042(n406 ,n9[19]);
    nor g2043(n1329 ,n375 ,n1324);
    nor g2044(n766 ,n117 ,n101);
    xnor g2045(n621 ,n20[23] ,n24[23]);
    or g2046(n873 ,n183 ,n640);
    nor g2047(n1648 ,n879 ,n1445);
    or g2048(n1105 ,n277 ,n640);
    not g2049(n310 ,n24[25]);
    or g2050(n1870 ,n1680 ,n1600);
    nor g2051(n1099 ,n226 ,n102);
    nor g2052(n825 ,n241 ,n98);
    nor g2053(n1670 ,n1103 ,n1445);
    not g2054(n260 ,n30[29]);
    buf g2055(n14[21], n10[17]);
    nor g2056(n735 ,n301 ,n104);
    dff g2057(.RN(n2058), .SN(1'b1), .CK(n0), .D(n448), .Q(n29[0]));
    or g2058(n1537 ,n1423 ,n1422);
    or g2059(n1156 ,n743 ,n1038);
    not g2060(n217 ,n28[6]);
    dff g2061(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1860), .Q(n22[29]));
    or g2062(n1991 ,n570 ,n1572);
    nor g2063(n722 ,n294 ,n96);
    nor g2064(n1015 ,n335 ,n101);
    or g2065(n1243 ,n925 ,n670);
    or g2066(n1109 ,n254 ,n640);
    dff g2067(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1139), .Q(n24[30]));
    nor g2068(n581 ,n176 ,n3);
    or g2069(n1931 ,n1739 ,n1642);
    dff g2070(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1291), .Q(n24[25]));
    nor g2071(n1580 ,n885 ,n1445);
    nor g2072(n1761 ,n514 ,n1444);
    dff g2073(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2002), .Q(n25[23]));
    nor g2074(n901 ,n321 ,n104);
    nor g2075(n860 ,n652 ,n599);
    or g2076(n1242 ,n922 ,n669);
    buf g2077(n18[8], 1'b0);
    buf g2078(n18[12], n10[0]);
    or g2079(n1245 ,n944 ,n1014);
    nor g2080(n1595 ,n883 ,n1443);
    or g2081(n1839 ,n690 ,n1779);
    or g2082(n1161 ,n733 ,n1040);
    not g2083(n273 ,n30[15]);
    buf g2084(n11[27], n10[27]);
    nor g2085(n561 ,n267 ,n3);
    not g2086(n81 ,n80);
    dff g2087(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1230), .Q(n13[15]));
    nor g2088(n1816 ,n360 ,n1447);
    not g2089(n223 ,n13[1]);
    dff g2090(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1876), .Q(n22[21]));
    nor g2091(n828 ,n238 ,n102);
    nor g2092(n1343 ,n641 ,n1320);
    xnor g2093(n612 ,n20[13] ,n24[13]);
    nor g2094(n1618 ,n1115 ,n1443);
    not g2095(n140 ,n25[7]);
    not g2096(n209 ,n30[14]);
    dff g2097(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1231), .Q(n13[14]));
    or g2098(n1286 ,n804 ,n781);
    or g2099(n1138 ,n955 ,n1019);
    or g2100(n2036 ,n1535 ,n1972);
    dff g2101(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2073), .Q(n29[3]));
    dff g2102(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1204), .Q(n24[19]));
    dff g2103(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1335), .Q(n15[3]));
    or g2104(n1313 ,n638 ,n714);
    dff g2105(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2030), .Q(n9[21]));
    nor g2106(n977 ,n122 ,n100);
    not g2107(n473 ,n12[25]);
    not g2108(n287 ,n2063);
    nor g2109(n1679 ,n377 ,n1442);
    nor g2110(n85 ,n29[4] ,n83);
    dff g2111(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1251), .Q(n24[31]));
    nor g2112(n1094 ,n288 ,n638);
    or g2113(n1364 ,n94 ,n1356);
    nor g2114(n1043 ,n362 ,n106);
    or g2115(n1988 ,n583 ,n1566);
    dff g2116(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1140), .Q(n24[29]));
    not g2117(n119 ,n24[15]);
    not g2118(n229 ,n10[5]);
    buf g2119(n14[3], 1'b0);
    dff g2120(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1221), .Q(n20[6]));
    nor g2121(n588 ,n467 ,n3);
    not g2122(n1324 ,n1325);
    not g2123(n484 ,n13[25]);
    nor g2124(n708 ,n638 ,n613);
    or g2125(n1544 ,n1405 ,n1438);
    nor g2126(n1694 ,n159 ,n1442);
    nor g2127(n1729 ,n408 ,n1440);
    nor g2128(n934 ,n427 ,n102);
    nor g2129(n577 ,n259 ,n3);
    nor g2130(n964 ,n182 ,n102);
    or g2131(n1305 ,n970 ,n1091);
    or g2132(n1939 ,n1747 ,n1649);
    nor g2133(n848 ,n126 ,n594);
    or g2134(n1983 ,n536 ,n1554);
    nor g2135(n1346 ,n1342 ,n1325);
    or g2136(n1300 ,n943 ,n996);
    nor g2137(n1467 ,n452 ,n1371);
    nor g2138(n847 ,n101 ,n597);
    nor g2139(n569 ,n215 ,n3);
    not g2140(n493 ,n9[16]);
    not g2141(n511 ,n13[30]);
    nor g2142(n996 ,n317 ,n101);
    dff g2143(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1956), .Q(n28[5]));
    not g2144(n560 ,n559);
    or g2145(n1296 ,n938 ,n1001);
    or g2146(n540 ,n4[31] ,n4[30]);
    not g2147(n87 ,n86);
    or g2148(n2055 ,n1573 ,n1991);
    not g2149(n146 ,n25[12]);
    nor g2150(n1738 ,n485 ,n1444);
    dff g2151(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2045), .Q(n9[5]));
    nor g2152(n1643 ,n883 ,n1445);
    dff g2153(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1862), .Q(n22[28]));
    dff g2154(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1254), .Q(n18[3]));
    not g2155(n502 ,n30[22]);
    or g2156(n1966 ,n550 ,n1522);
    buf g2157(n14[27], n10[23]);
    dff g2158(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1309), .Q(n14[5]));
    not g2159(n412 ,n9[28]);
    nor g2160(n791 ,n246 ,n102);
    not g2161(n507 ,n13[15]);
    nor g2162(n643 ,n555 ,n557);
    nor g2163(n729 ,n297 ,n103);
    nor g2164(n1383 ,n199 ,n1371);
    nor g2165(n574 ,n478 ,n3);
    xnor g2166(n617 ,n20[26] ,n24[26]);
    nor g2167(n1489 ,n382 ,n1369);
    or g2168(n1261 ,n945 ,n997);
    or g2169(n2026 ,n1515 ,n1962);
    nor g2170(n1438 ,n404 ,n1370);
    nor g2171(n675 ,n97 ,n611);
    or g2172(n1577 ,n1512 ,n1511);
    nor g2173(n1584 ,n873 ,n1445);
    nor g2174(n813 ,n394 ,n99);
    nor g2175(n53 ,n49 ,n46);
    nor g2176(n1378 ,n251 ,n1370);
    nor g2177(n922 ,n491 ,n98);
    dff g2178(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1293), .Q(n10[23]));
    or g2179(n1934 ,n1741 ,n1644);
    nor g2180(n1034 ,n348 ,n106);
    not g2181(n106 ,n104);
    dff g2182(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1874), .Q(n22[22]));
    or g2183(n1362 ,n94 ,n1347);
    not g2184(n137 ,n2);
    or g2185(n1921 ,n1729 ,n1673);
    or g2186(n1209 ,n868 ,n847);
    not g2187(n2086 ,n24[13]);
    or g2188(n1885 ,n1693 ,n1614);
    nor g2189(n1644 ,n1100 ,n1445);
    dff g2190(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1306), .Q(n14[4]));
    nor g2191(n1785 ,n151 ,n1447);
    or g2192(n1936 ,n1744 ,n1672);
    buf g2193(n11[18], n10[18]);
    not g2194(n462 ,n28[26]);
    dff g2195(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2014), .Q(n25[11]));
    or g2196(n1977 ,n581 ,n1545);
    or g2197(n1370 ,n107 ,n1362);
    nor g2198(n818 ,n456 ,n99);
    dff g2199(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1885), .Q(n22[12]));
    nor g2200(n1025 ,n380 ,n106);
    nor g2201(n782 ,n113 ,n101);
    not g2202(n103 ,n106);
    dff g2203(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1167), .Q(n27[7]));
    nor g2204(n1096 ,n284 ,n638);
    nor g2205(n59 ,n48 ,n57);
    or g2206(n93 ,n646 ,n1326);
    or g2207(n538 ,n4[21] ,n4[20]);
    not g2208(n269 ,n9[31]);
    buf g2209(n11[26], n10[26]);
    or g2210(n1965 ,n565 ,n1520);
    or g2211(n1853 ,n700 ,n1808);
    not g2212(n296 ,n24[18]);
    not g2213(n274 ,n30[9]);
    or g2214(n1548 ,n1451 ,n1452);
    dff g2215(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1227), .Q(n15[7]));
    nor g2216(n927 ,n477 ,n98);
    or g2217(n1519 ,n1385 ,n1384);
    nor g2218(n1330 ,n355 ,n1324);
    nor g2219(n1496 ,n359 ,n1368);
    nor g2220(n1586 ,n876 ,n1445);
    nor g2221(n1775 ,n169 ,n1446);
    not g2222(n245 ,n14[6]);
    nor g2223(n966 ,n494 ,n639);
    dff g2224(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1178), .Q(n20[20]));
    nor g2225(n572 ,n450 ,n3);
    not g2226(n193 ,n5[8]);
    dff g2227(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1946), .Q(n28[15]));
    nor g2228(n1483 ,n361 ,n1369);
    nor g2229(n1387 ,n502 ,n1371);
    not g2230(n220 ,n10[10]);
    or g2231(n1901 ,n1709 ,n1602);
    or g2232(n1117 ,n177 ,n640);
    not g2233(n415 ,n9[21]);
    or g2234(n1143 ,n800 ,n1023);
    or g2235(n1902 ,n1710 ,n1592);
    dff g2236(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2043), .Q(n9[7]));
    nor g2237(n1767 ,n191 ,n1444);
    or g2238(n1303 ,n968 ,n1092);
    or g2239(n1849 ,n707 ,n1800);
    dff g2240(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1294), .Q(n10[1]));
    or g2241(n1229 ,n901 ,n1077);
    nor g2242(n1725 ,n235 ,n1440);
    or g2243(n2092 ,n2081 ,n24[15]);
    not g2244(n305 ,n24[20]);
    not g2245(n301 ,n24[12]);
    dff g2246(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2026), .Q(n9[24]));
    or g2247(n539 ,n4[7] ,n4[6]);
    or g2248(n1146 ,n752 ,n1027);
    or g2249(n1236 ,n911 ,n667);
    nor g2250(n1810 ,n254 ,n1446);
    nor g2251(n945 ,n405 ,n102);
    dff g2252(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2069), .Q(n29[7]));
    nor g2253(n1508 ,n376 ,n1369);
    not g2254(n203 ,n28[27]);
    or g2255(n1104 ,n187 ,n640);
    nor g2256(n985 ,n330 ,n101);
    nor g2257(n704 ,n638 ,n606);
    dff g2258(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2042), .Q(n9[8]));
    buf g2259(n1340 ,n641);
    not g2260(n139 ,n22[29]);
    or g2261(n1994 ,n1771 ,n1834);
    not g2262(n271 ,n10[25]);
    dff g2263(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1136), .Q(n20[30]));
    nor g2264(n1022 ,n144 ,n105);
    buf g2265(n11[24], n10[24]);
    or g2266(n564 ,n129 ,n4[2]);
    dff g2267(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1377), .Q(n23[0]));
    xor g2268(n2069 ,n29[7] ,n92);
    nor g2269(n821 ,n264 ,n102);
    dff g2270(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1212), .Q(n13[28]));
    not g2271(n487 ,n30[27]);
    or g2272(n523 ,n8[7] ,n8[6]);
    dff g2273(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1933), .Q(n28[26]));
    nor g2274(n1011 ,n332 ,n101);
    not g2275(n348 ,n25[3]);
    nor g2276(n1379 ,n262 ,n1371);
    nor g2277(n1782 ,n196 ,n1446);
    dff g2278(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1950), .Q(n28[12]));
    nor g2279(n1511 ,n249 ,n1370);
    nor g2280(n559 ,n293 ,n23[0]);
    not g2281(n505 ,n10[13]);
    nor g2282(n1800 ,n200 ,n1446);
    or g2283(n2012 ,n1807 ,n1852);
    dff g2284(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1871), .Q(n22[24]));
    nor g2285(n1707 ,n472 ,n1440);
    or g2286(n1284 ,n927 ,n990);
    nor g2287(n1777 ,n359 ,n1447);
    nor g2288(n1454 ,n490 ,n1371);
    or g2289(n1113 ,n189 ,n640);
    or g2290(n1134 ,n737 ,n1045);
    nor g2291(n989 ,n370 ,n101);
    dff g2292(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1247), .Q(n12[29]));
    not g2293(n128 ,n20[14]);
    nor g2294(n1031 ,n346 ,n106);
    nor g2295(n1476 ,n349 ,n1368);
    or g2296(n533 ,n15[6] ,n15[7]);
    nor g2297(n1703 ,n374 ,n1442);
    or g2298(n1287 ,n803 ,n978);
    or g2299(n1556 ,n1465 ,n1468);
    or g2300(n1356 ,n637 ,n93);
    not g2301(n125 ,n20[9]);
    nor g2302(n929 ,n508 ,n102);
    dff g2303(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1907), .Q(n30[22]));
    or g2304(n1552 ,n1459 ,n1460);
    not g2305(n201 ,n13[16]);
    or g2306(n1951 ,n1759 ,n1659);
    not g2307(n328 ,n20[25]);
    not g2308(n204 ,n9[10]);
    nor g2309(n1079 ,n374 ,n105);
    nor g2310(n1453 ,n175 ,n1370);
    nor g2311(n983 ,n123 ,n96);
    nor g2312(n1814 ,n390 ,n1447);
    not g2313(n387 ,n22[28]);
    dff g2314(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1228), .Q(n13[16]));
    not g2315(n149 ,n22[14]);
    or g2316(n1332 ,n1266 ,n1265);
    nor g2317(n1492 ,n139 ,n1369);
    dff g2318(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1149), .Q(n24[22]));
    or g2319(n1576 ,n1483 ,n1509);
    dff g2320(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1248), .Q(n12[27]));
    or g2321(n1276 ,n959 ,n991);
    or g2322(n1528 ,n1404 ,n1439);
    or g2323(n1674 ,n1508 ,n1510);
    nor g2324(n1003 ,n383 ,n96);
    nor g2325(n1696 ,n342 ,n1442);
    nor g2326(n1827 ,n186 ,n1446);
    nor g2327(n1790 ,n233 ,n1446);
    dff g2328(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1879), .Q(n22[18]));
    buf g2329(n11[23], n10[23]);
    not g2330(n503 ,n13[2]);
    nor g2331(n1421 ,n160 ,n1368);
    not g2332(n443 ,n9[4]);
    dff g2333(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2044), .Q(n9[6]));
    not g2334(n47 ,n27[4]);
    nor g2335(n978 ,n321 ,n101);
    buf g2336(n18[4], n14[4]);
    dff g2337(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1143), .Q(n20[29]));
    nor g2338(n768 ,n119 ,n101);
    nor g2339(n1457 ,n217 ,n1370);
    not g2340(n172 ,n2061);
    dff g2341(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1162), .Q(n24[13]));
    dff g2342(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1175), .Q(n27[1]));
    nor g2343(n1663 ,n1114 ,n1445);
    nor g2344(n890 ,n232 ,n98);
    nor g2345(n1391 ,n399 ,n1371);
    nor g2346(n1639 ,n1104 ,n1441);
    nor g2347(n1687 ,n365 ,n1442);
    not g2348(n284 ,n2068);
    nor g2349(n992 ,n135 ,n101);
    or g2350(n2056 ,n1575 ,n1992);
    dff g2351(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1312), .Q(n11[11]));
    nor g2352(n1409 ,n386 ,n1368);
    or g2353(n1955 ,n1763 ,n1664);
    or g2354(n1874 ,n1683 ,n1604);
    not g2355(n336 ,n20[22]);
    not g2356(n464 ,n13[29]);
    or g2357(n1900 ,n1708 ,n1596);
    or g2358(n884 ,n178 ,n640);
    dff g2359(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1252), .Q(n12[23]));
    not g2360(n404 ,n28[9]);
    or g2361(n1315 ,n638 ,n716);
    not g2362(n371 ,n15[5]);
    not g2363(n126 ,n21[3]);
    not g2364(n1373 ,n1372);
    nor g2365(n761 ,n308 ,n101);
    nor g2366(n1742 ,n203 ,n1444);
    nor g2367(n1638 ,n1111 ,n1441);
    nor g2368(n1053 ,n143 ,n106);
    not g2369(n200 ,n5[16]);
    nor g2370(n968 ,n482 ,n639);
    or g2371(n1108 ,n213 ,n640);
    or g2372(n1191 ,n831 ,n786);
    not g2373(n181 ,n28[29]);
    not g2374(n72 ,n29[3]);
    buf g2375(n18[14], n10[2]);
    dff g2376(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2036), .Q(n9[14]));
    nor g2377(n1717 ,n420 ,n1440);
    dff g2378(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1275), .Q(n11[0]));
    or g2379(n1949 ,n1758 ,n1662);
    or g2380(n1288 ,n962 ,n1008);
    or g2381(n1249 ,n937 ,n780);
    dff g2382(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1270), .Q(n18[1]));
    nor g2383(n869 ,n341 ,n643);
    dff g2384(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1916), .Q(n30[13]));
    nor g2385(n64 ,n27[5] ,n62);
    nor g2386(n1085 ,n152 ,n106);
    nor g2387(n1317 ,n8[0] ,n1098);
    nor g2388(n1714 ,n199 ,n1440);
    not g2389(n345 ,n15[2]);
    not g2390(n364 ,n25[27]);
    dff g2391(.RN(n2058), .SN(1'b1), .CK(n0), .D(n2074), .Q(n29[2]));
    not g2392(n485 ,n28[31]);
    nor g2393(n804 ,n234 ,n99);
    or g2394(n1216 ,n928 ,n1071);
    nor g2395(n831 ,n454 ,n102);
    not g2396(n157 ,n25[17]);
    xnor g2397(n604 ,n20[25] ,n24[25]);
    nor g2398(n1684 ,n343 ,n1442);
    dff g2399(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1931), .Q(n28[30]));
    or g2400(n1265 ,n789 ,n989);
    or g2401(n1259 ,n946 ,n774);
    dff g2402(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1887), .Q(n22[10]));
    nor g2403(n1035 ,n350 ,n106);
    not g2404(n486 ,n14[1]);
    dff g2405(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1237), .Q(n13[8]));
    or g2406(n1151 ,n740 ,n1081);
    nor g2407(n664 ,n97 ,n614);
    nor g2408(n1646 ,n1101 ,n1445);
    or g2409(n2030 ,n1521 ,n1965);
    xnor g2410(n636 ,n108 ,n164);
    nor g2411(n1415 ,n273 ,n1371);
    dff g2412(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1242), .Q(n13[4]));
    dff g2413(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1271), .Q(n10[14]));
    nor g2414(n1058 ,n386 ,n105);
    or g2415(n1876 ,n1684 ,n1605);
    not g2416(n337 ,n20[7]);
    dff g2417(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1153), .Q(n20[26]));
    nor g2418(n1050 ,n289 ,n105);
    nor g2419(n1478 ,n397 ,n1371);
    not g2420(n54 ,n53);
    nor g2421(n931 ,n228 ,n99);
    nor g2422(n1700 ,n357 ,n1442);
    or g2423(n1985 ,n590 ,n1560);
    not g2424(n405 ,n18[2]);
    not g2425(n186 ,n5[3]);
    nor g2426(n857 ,n650 ,n601);
    nor g2427(n1829 ,n143 ,n1447);
    or g2428(n1136 ,n936 ,n1020);
    or g2429(n1895 ,n1704 ,n1624);
    nor g2430(n52 ,n27[1] ,n27[0]);
    nor g2431(n690 ,n638 ,n617);
    nor g2432(n725 ,n306 ,n103);
    not g2433(n247 ,n5[0]);
    nor g2434(n999 ,n130 ,n101);
    or g2435(n2093 ,n24[29] ,n24[28]);
    nor g2436(n686 ,n638 ,n620);
    nor g2437(n724 ,n313 ,n103);
    or g2438(n648 ,n542 ,n541);
    or g2439(n1903 ,n1711 ,n1628);
    not g2440(n449 ,n10[31]);
    or g2441(n2040 ,n1543 ,n1976);
    nor g2442(n1620 ,n1112 ,n1443);
    not g2443(n334 ,n20[15]);
    nor g2444(n868 ,n511 ,n99);
    dff g2445(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1159), .Q(n24[3]));
    or g2446(n1858 ,n708 ,n1814);
    not g2447(n361 ,n22[25]);
    nor g2448(n1808 ,n189 ,n1446);
    not g2449(n163 ,n22[15]);
    xnor g2450(n615 ,n20[5] ,n24[5]);
    nor g2451(n1412 ,n163 ,n1369);
    or g2452(n626 ,n571 ,n95);
    or g2453(n1365 ,n94 ,n1354);
    or g2454(n1877 ,n1685 ,n1606);
    or g2455(n1126 ,n826 ,n758);
    nor g2456(n829 ,n122 ,n103);
    nor g2457(n1473 ,n418 ,n1371);
    not g2458(n425 ,n30[26]);
    nor g2459(n1038 ,n157 ,n105);
    not g2460(n379 ,n15[7]);
    or g2461(n1950 ,n1757 ,n1658);
    nor g2462(n1033 ,n361 ,n105);
    nor g2463(n841 ,n223 ,n102);
    not g2464(n2058 ,n1);
    nor g2465(n1320 ,n534 ,n948);
    nor g2466(n1585 ,n1102 ,n1441);
    dff g2467(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1961), .Q(n28[0]));
    nor g2468(n753 ,n119 ,n103);
    or g2469(n1515 ,n1379 ,n1378);
    buf g2470(n18[9], 1'b0);
    nor g2471(n1718 ,n257 ,n1440);
    or g2472(n1888 ,n1696 ,n1617);
    not g2473(n494 ,n27[2]);
    nor g2474(n1783 ,n344 ,n1447);
    or g2475(n1891 ,n1700 ,n1620);
    nor g2476(n1749 ,n173 ,n1444);
    nor g2477(n89 ,n74 ,n87);
    or g2478(n948 ,n165 ,n645);
    or g2479(n1567 ,n1491 ,n1490);
    nor g2480(n1686 ,n347 ,n1442);
    not g2481(n50 ,n27[5]);
    dff g2482(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1954), .Q(n28[7]));
    not g2483(n642 ,n643);
    nor g2484(n888 ,n459 ,n98);
    buf g2485(n14[20], n10[16]);
    nor g2486(n669 ,n96 ,n616);
    nor g2487(n1068 ,n378 ,n106);
    nor g2488(n909 ,n379 ,n643);
    not g2489(n124 ,n20[31]);
    nor g2490(n1652 ,n875 ,n1445);
    or g2491(n1918 ,n1726 ,n1647);
    not g2492(n150 ,n25[31]);
    not g2493(n265 ,n30[16]);
    nor g2494(n1713 ,n262 ,n1440);
    nor g2495(n1076 ,n385 ,n105);
    nor g2496(n1778 ,n255 ,n1446);
    dff g2497(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1996), .Q(n25[29]));
    nor g2498(n1398 ,n446 ,n1370);
    or g2499(n101 ,n23[1] ,n560);
    nor g2500(n716 ,n651 ,n598);
    nor g2501(n855 ,n158 ,n643);
    or g2502(n1173 ,n812 ,n1036);
    or g2503(n1297 ,n967 ,n1094);
    or g2504(n1302 ,n912 ,n1015);
    not g2505(n234 ,n12[26]);
    nor g2506(n1798 ,n157 ,n1447);
    nor g2507(n1510 ,n151 ,n1368);
    or g2508(n1227 ,n641 ,n909);
    nor g2509(n1012 ,n323 ,n100);
    or g2510(n1223 ,n890 ,n679);
    or g2511(n1162 ,n728 ,n1042);
    nor g2512(n778 ,n309 ,n96);
    not g2513(n460 ,n11[8]);
    nor g2514(n1045 ,n166 ,n105);
    nor g2515(n1390 ,n282 ,n1370);
    or g2516(n1137 ,n806 ,n1006);
    not g2517(n38 ,n27[5]);
    or g2518(n1534 ,n1417 ,n1416);
    or g2519(n874 ,n185 ,n640);
    nor g2520(n1040 ,n388 ,n106);
    xnor g2521(n1119 ,n638 ,n27[0]);
    not g2522(n498 ,n28[1]);
    not g2523(n291 ,n2064);
    nor g2524(n1728 ,n274 ,n1440);
    or g2525(n1248 ,n939 ,n783);
    or g2526(n1218 ,n902 ,n676);
    nor g2527(n1823 ,n225 ,n1446);
    or g2528(n1975 ,n561 ,n1540);
    nor g2529(n693 ,n638 ,n607);
    dff g2530(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1902), .Q(n30[27]));
    or g2531(n94 ,n648 ,n647);
    nor g2532(n1624 ,n1106 ,n1443);
    not g2533(n444 ,n27[3]);
    not g2534(n652 ,n651);
    or g2535(n1986 ,n551 ,n1562);
    dff g2536(.RN(n2058), .SN(1'b1), .CK(n0), .D(n1196), .Q(n12[30]));
    nor g2537(n993 ,n134 ,n96);
    or g2538(n1929 ,n1736 ,n1639);
    nor g2539(n830 ,n97 ,n617);
    not g2540(n354 ,n25[10]);
    not g2541(n451 ,n11[0]);
    or g2542(n1993 ,n585 ,n1576);
    not g2543(n212 ,n5[22]);
endmodule
