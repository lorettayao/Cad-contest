module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11);
    input [127:0] n0;
    input [255:0] n1;
    input [63:0] n2;
    input [3:0] n3;
    input [31:0] n4;
    input [4:0] n5;
    input n6, n7, n8;
    output [127:0] n9;
    output [31:0] n10;
    output n11;
    wire [127:0] n0;
    wire [255:0] n1;
    wire [63:0] n2;
    wire [3:0] n3;
    wire [31:0] n4;
    wire [4:0] n5;
    wire n6, n7, n8;
    wire [127:0] n9;
    wire [31:0] n10;
    wire n11;
    wire n12, n13, n14, n15, n16, n17, n18, n19;
    wire n20, n21, n22, n23, n24, n25, n26, n27;
    wire n28, n29, n30, n31, n32, n33, n34, n35;
    wire n36, n37, n38, n39, n40, n41, n42, n43;
    wire n44, n45, n46, n47, n48, n49, n50, n51;
    wire n52, n53, n54, n55, n56, n57, n58, n59;
    wire n60, n61, n62, n63, n64, n65, n66, n67;
    wire n68, n69, n70, n71, n72, n73, n74, n75;
    wire n76, n77, n78, n79, n80, n81, n82, n83;
    wire n84, n85, n86, n87, n88, n89, n90, n91;
    wire n92, n93, n94, n95, n96, n97, n98, n99;
    wire n100, n101, n102, n103, n104, n105, n106, n107;
    wire n108, n109, n110, n111, n112, n113, n114, n115;
    wire n116, n117, n118, n119, n120, n121, n122, n123;
    wire n124, n125, n126, n127, n128, n129, n130, n131;
    wire n132, n133, n134, n135, n136, n137, n138, n139;
    wire n140, n141, n142, n143, n144, n145, n146, n147;
    wire n148, n149, n150, n151, n152, n153, n154, n155;
    wire n156, n157, n158, n159, n160, n161, n162, n163;
    wire n164, n165, n166, n167, n168, n169, n170, n171;
    wire n172, n173, n174, n175, n176, n177, n178, n179;
    wire n180, n181, n182, n183, n184, n185, n186, n187;
    wire n188, n189, n190, n191, n192, n193, n194, n195;
    wire n196, n197, n198, n199, n200, n201, n202, n203;
    wire n204, n205, n206, n207, n208, n209, n210, n211;
    wire n212, n213, n214, n215, n216, n217, n218, n219;
    wire n220, n221, n222, n223, n224, n225, n226, n227;
    wire n228, n229, n230, n231, n232, n233, n234, n235;
    wire n236, n237, n238, n239, n240, n241, n242, n243;
    wire n244, n245, n246, n247, n248, n249, n250, n251;
    wire n252, n253, n254, n255, n256, n257, n258, n259;
    wire n260, n261, n262, n263, n264, n265, n266, n267;
    wire n268, n269, n270, n271, n272, n273, n274, n275;
    wire n276, n277, n278, n279, n280, n281, n282, n283;
    wire n284, n285, n286, n287, n288, n289, n290, n291;
    wire n292, n293, n294, n295, n296, n297, n298, n299;
    wire n300, n301, n302, n303, n304, n305, n306, n307;
    wire n308, n309, n310, n311, n312, n313, n314, n315;
    wire n316, n317, n318, n319, n320, n321, n322, n323;
    wire n324, n325, n326, n327, n328, n329, n330, n331;
    wire n332, n333, n334, n335, n336, n337, n338, n339;
    wire n340, n341, n342, n343, n344, n345, n346, n347;
    wire n348, n349, n350, n351, n352, n353, n354, n355;
    wire n356, n357, n358, n359, n360, n361, n362, n363;
    wire n364, n365, n366, n367, n368, n369, n370, n371;
    wire n372, n373, n374, n375, n376, n377, n378, n379;
    wire n380, n381, n382, n383, n384, n385, n386, n387;
    wire n388, n389, n390, n391, n392, n393, n394, n395;
    wire n396, n397, n398, n399, n400, n401, n402, n403;
    wire n404, n405, n406, n407, n408, n409, n410, n411;
    wire n412, n413, n414, n415, n416, n417, n418, n419;
    wire n420, n421, n422, n423, n424, n425, n426, n427;
    wire n428, n429, n430, n431, n432, n433, n434, n435;
    wire n436, n437, n438, n439, n440, n441, n442, n443;
    wire n444, n445, n446, n447, n448, n449, n450, n451;
    wire n452, n453, n454, n455, n456, n457, n458, n459;
    wire n460, n461, n462, n463, n464, n465, n466, n467;
    wire n468, n469, n470, n471, n472, n473, n474, n475;
    wire n476, n477, n478, n479, n480, n481, n482, n483;
    wire n484, n485, n486, n487, n488, n489, n490, n491;
    wire n492, n493, n494, n495, n496, n497, n498, n499;
    wire n500, n501, n502, n503, n504, n505, n506, n507;
    wire n508, n509, n510, n511, n512, n513, n514, n515;
    wire n516, n517, n518, n519, n520, n521, n522, n523;
    wire n524, n525, n526, n527, n528, n529, n530, n531;
    wire n532, n533, n534, n535, n536, n537, n538, n539;
    wire n540, n541, n542, n543, n544, n545, n546, n547;
    wire n548, n549, n550, n551, n552, n553, n554, n555;
    wire n556, n557, n558, n559, n560, n561, n562, n563;
    wire n564, n565, n566, n567, n568, n569, n570, n571;
    wire n572, n573, n574, n575, n576, n577, n578, n579;
    wire n580, n581, n582, n583, n584, n585, n586, n587;
    wire n588, n589, n590, n591, n592, n593, n594, n595;
    wire n596, n597, n598, n599, n600, n601, n602, n603;
    wire n604, n605, n606, n607, n608, n609, n610, n611;
    wire n612, n613, n614, n615, n616, n617, n618, n619;
    wire n620, n621, n622, n623, n624, n625, n626, n627;
    wire n628, n629, n630, n631, n632, n633, n634, n635;
    wire n636, n637, n638, n639, n640, n641, n642, n643;
    wire n644, n645, n646, n647, n648, n649, n650, n651;
    wire n652, n653, n654, n655, n656, n657, n658, n659;
    wire n660, n661, n662, n663, n664, n665, n666, n667;
    wire n668, n669, n670, n671, n672, n673, n674, n675;
    wire n676, n677, n678, n679, n680, n681, n682, n683;
    wire n684, n685, n686, n687, n688, n689, n690, n691;
    wire n692, n693, n694, n695, n696, n697, n698, n699;
    wire n700, n701, n702, n703, n704, n705, n706, n707;
    wire n708, n709, n710, n711, n712, n713, n714, n715;
    wire n716, n717, n718, n719, n720, n721, n722, n723;
    wire n724, n725, n726, n727, n728, n729, n730, n731;
    wire n732, n733, n734, n735, n736, n737, n738, n739;
    wire n740, n741, n742, n743, n744, n745, n746, n747;
    wire n748, n749, n750, n751, n752, n753, n754, n755;
    wire n756, n757, n758, n759, n760, n761, n762, n763;
    wire n764, n765, n766, n767, n768, n769, n770, n771;
    wire n772, n773, n774, n775, n776, n777, n778, n779;
    wire n780, n781, n782, n783, n784, n785, n786, n787;
    wire n788, n789, n790, n791, n792, n793, n794, n795;
    wire n796, n797, n798, n799, n800, n801, n802, n803;
    wire n804, n805, n806, n807, n808, n809, n810, n811;
    wire n812, n813, n814, n815, n816, n817, n818, n819;
    wire n820, n821, n822, n823, n824, n825, n826, n827;
    wire n828, n829, n830, n831, n832, n833, n834, n835;
    wire n836, n837, n838, n839, n840, n841, n842, n843;
    wire n844, n845, n846, n847, n848, n849, n850, n851;
    wire n852, n853, n854, n855, n856, n857, n858, n859;
    wire n860, n861, n862, n863, n864, n865, n866, n867;
    wire n868, n869, n870, n871, n872, n873, n874, n875;
    wire n876, n877, n878, n879, n880, n881, n882, n883;
    wire n884, n885, n886, n887, n888, n889, n890, n891;
    wire n892, n893, n894, n895, n896, n897, n898, n899;
    wire n900, n901, n902, n903, n904, n905, n906, n907;
    wire n908, n909, n910, n911, n912, n913, n914, n915;
    wire n916, n917, n918, n919, n920, n921, n922, n923;
    wire n924, n925, n926, n927, n928, n929, n930, n931;
    wire n932, n933, n934, n935, n936, n937, n938, n939;
    wire n940, n941, n942, n943, n944, n945, n946, n947;
    wire n948, n949, n950, n951, n952, n953, n954, n955;
    wire n956, n957, n958, n959, n960, n961, n962, n963;
    wire n964, n965, n966, n967, n968, n969, n970, n971;
    wire n972, n973, n974, n975, n976, n977, n978, n979;
    wire n980, n981, n982, n983, n984, n985, n986, n987;
    wire n988, n989, n990, n991, n992, n993, n994, n995;
    wire n996, n997, n998, n999, n1000, n1001, n1002, n1003;
    wire n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011;
    wire n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
    wire n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
    wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
    wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
    wire n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051;
    wire n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
    wire n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067;
    wire n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075;
    wire n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083;
    wire n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;
    wire n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099;
    wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107;
    wire n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115;
    wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
    wire n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131;
    wire n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139;
    wire n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147;
    wire n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155;
    wire n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163;
    wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171;
    wire n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179;
    wire n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187;
    wire n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195;
    wire n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203;
    wire n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211;
    wire n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219;
    wire n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227;
    wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235;
    wire n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243;
    wire n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251;
    wire n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259;
    wire n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267;
    wire n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
    wire n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283;
    wire n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291;
    wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299;
    wire n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307;
    wire n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315;
    wire n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323;
    wire n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331;
    wire n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339;
    wire n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347;
    wire n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355;
    wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363;
    wire n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371;
    wire n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379;
    wire n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387;
    wire n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395;
    wire n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403;
    wire n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411;
    wire n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419;
    wire n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427;
    wire n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435;
    wire n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443;
    wire n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451;
    wire n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459;
    wire n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467;
    wire n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475;
    wire n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
    wire n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491;
    wire n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499;
    wire n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507;
    wire n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515;
    wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
    wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;
    wire n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539;
    wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
    wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
    wire n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563;
    wire n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571;
    wire n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579;
    wire n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587;
    wire n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595;
    wire n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603;
    wire n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611;
    wire n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619;
    wire n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627;
    wire n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635;
    wire n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643;
    wire n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651;
    wire n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659;
    wire n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667;
    wire n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675;
    wire n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683;
    wire n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691;
    wire n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699;
    wire n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707;
    wire n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715;
    wire n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723;
    wire n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731;
    wire n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739;
    wire n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747;
    wire n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755;
    wire n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763;
    wire n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771;
    wire n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779;
    wire n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787;
    wire n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795;
    wire n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803;
    wire n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811;
    wire n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819;
    wire n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827;
    wire n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835;
    wire n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843;
    wire n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851;
    wire n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859;
    wire n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867;
    wire n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
    wire n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883;
    wire n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891;
    wire n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899;
    wire n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907;
    wire n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915;
    wire n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923;
    wire n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931;
    wire n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939;
    wire n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947;
    wire n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955;
    wire n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963;
    wire n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971;
    wire n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979;
    wire n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987;
    wire n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995;
    wire n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;
    wire n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011;
    wire n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019;
    wire n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027;
    wire n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035;
    wire n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043;
    wire n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051;
    wire n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059;
    wire n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067;
    wire n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075;
    wire n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083;
    wire n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091;
    wire n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099;
    wire n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107;
    wire n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115;
    wire n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123;
    wire n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131;
    wire n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139;
    wire n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147;
    wire n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155;
    wire n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163;
    wire n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
    wire n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179;
    wire n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187;
    wire n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195;
    wire n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203;
    wire n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211;
    wire n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219;
    wire n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227;
    wire n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235;
    wire n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243;
    wire n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251;
    wire n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259;
    wire n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267;
    wire n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275;
    wire n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283;
    wire n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291;
    wire n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299;
    wire n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307;
    wire n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315;
    wire n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323;
    wire n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331;
    wire n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339;
    wire n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347;
    wire n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355;
    wire n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363;
    wire n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371;
    wire n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379;
    wire n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387;
    wire n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395;
    wire n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403;
    wire n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411;
    wire n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419;
    wire n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427;
    wire n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435;
    wire n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443;
    wire n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451;
    wire n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459;
    wire n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467;
    wire n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475;
    wire n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483;
    wire n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491;
    wire n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499;
    wire n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507;
    wire n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515;
    wire n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523;
    wire n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531;
    wire n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539;
    wire n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547;
    wire n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555;
    wire n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563;
    wire n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571;
    wire n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579;
    wire n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587;
    wire n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595;
    wire n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603;
    wire n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611;
    wire n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619;
    wire n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627;
    wire n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635;
    wire n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643;
    wire n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651;
    wire n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659;
    wire n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667;
    wire n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675;
    wire n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683;
    wire n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691;
    wire n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699;
    wire n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707;
    wire n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715;
    wire n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723;
    wire n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731;
    wire n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739;
    wire n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747;
    wire n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755;
    wire n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763;
    wire n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771;
    wire n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779;
    wire n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787;
    wire n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795;
    wire n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803;
    wire n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811;
    wire n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819;
    wire n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827;
    wire n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835;
    wire n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843;
    wire n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851;
    wire n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859;
    wire n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867;
    wire n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875;
    wire n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883;
    wire n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891;
    wire n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899;
    wire n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907;
    wire n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915;
    wire n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923;
    wire n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931;
    wire n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939;
    wire n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947;
    wire n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955;
    wire n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963;
    wire n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971;
    wire n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979;
    wire n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987;
    wire n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995;
    wire n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003;
    wire n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011;
    wire n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019;
    wire n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027;
    wire n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035;
    wire n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043;
    wire n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051;
    wire n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059;
    wire n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067;
    wire n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075;
    wire n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083;
    wire n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091;
    wire n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099;
    wire n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107;
    wire n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115;
    wire n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123;
    wire n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131;
    wire n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139;
    wire n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147;
    wire n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155;
    wire n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163;
    wire n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171;
    wire n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179;
    wire n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187;
    wire n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195;
    wire n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203;
    wire n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211;
    wire n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219;
    wire n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227;
    wire n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235;
    wire n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243;
    wire n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251;
    wire n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259;
    wire n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267;
    wire n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275;
    wire n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283;
    wire n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291;
    wire n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299;
    wire n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307;
    wire n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315;
    wire n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323;
    wire n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331;
    wire n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339;
    wire n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347;
    wire n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355;
    wire n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363;
    wire n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371;
    wire n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379;
    wire n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387;
    wire n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395;
    wire n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403;
    wire n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411;
    wire n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419;
    wire n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427;
    wire n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435;
    wire n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443;
    wire n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451;
    wire n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459;
    wire n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467;
    wire n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475;
    wire n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483;
    wire n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491;
    wire n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499;
    wire n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507;
    wire n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515;
    wire n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523;
    wire n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531;
    wire n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539;
    wire n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547;
    wire n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555;
    wire n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563;
    wire n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571;
    wire n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579;
    wire n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587;
    wire n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595;
    wire n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603;
    wire n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611;
    wire n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619;
    wire n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627;
    wire n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635;
    wire n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643;
    wire n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651;
    wire n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659;
    wire n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667;
    wire n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675;
    wire n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683;
    wire n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691;
    wire n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699;
    wire n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707;
    wire n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715;
    wire n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723;
    wire n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731;
    wire n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739;
    wire n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747;
    wire n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755;
    wire n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763;
    wire n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771;
    wire n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779;
    wire n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787;
    wire n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795;
    wire n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803;
    wire n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811;
    wire n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819;
    wire n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827;
    wire n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835;
    wire n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843;
    wire n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851;
    wire n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859;
    wire n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867;
    wire n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875;
    wire n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883;
    wire n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891;
    wire n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899;
    wire n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907;
    wire n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915;
    wire n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923;
    wire n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931;
    wire n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939;
    wire n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947;
    wire n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955;
    wire n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963;
    wire n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971;
    wire n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979;
    wire n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987;
    wire n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995;
    wire n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003;
    wire n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011;
    wire n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019;
    wire n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027;
    wire n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035;
    wire n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043;
    wire n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051;
    wire n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059;
    wire n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067;
    wire n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075;
    wire n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083;
    wire n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091;
    wire n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099;
    wire n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107;
    wire n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115;
    wire n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123;
    wire n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131;
    wire n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139;
    wire n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147;
    wire n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155;
    wire n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163;
    wire n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171;
    wire n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179;
    wire n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187;
    wire n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195;
    wire n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203;
    wire n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211;
    wire n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219;
    wire n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227;
    wire n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235;
    wire n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243;
    wire n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251;
    wire n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259;
    wire n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267;
    wire n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275;
    wire n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283;
    wire n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291;
    wire n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299;
    wire n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307;
    wire n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315;
    wire n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323;
    wire n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331;
    wire n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339;
    wire n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347;
    wire n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355;
    wire n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363;
    wire n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371;
    wire n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379;
    wire n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387;
    wire n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395;
    wire n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403;
    wire n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411;
    wire n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419;
    wire n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427;
    wire n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435;
    wire n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443;
    wire n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451;
    wire n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459;
    wire n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467;
    wire n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475;
    wire n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483;
    wire n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491;
    wire n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499;
    wire n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507;
    wire n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515;
    wire n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523;
    wire n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531;
    wire n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539;
    wire n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547;
    wire n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555;
    wire n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563;
    wire n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571;
    wire n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579;
    wire n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587;
    wire n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595;
    wire n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603;
    wire n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611;
    wire n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619;
    wire n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627;
    wire n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635;
    wire n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643;
    wire n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651;
    wire n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659;
    wire n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667;
    wire n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675;
    wire n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683;
    wire n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691;
    wire n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699;
    wire n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707;
    wire n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715;
    wire n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723;
    wire n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731;
    wire n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739;
    wire n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747;
    wire n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755;
    wire n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763;
    wire n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771;
    wire n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779;
    wire n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787;
    wire n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795;
    wire n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803;
    wire n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811;
    wire n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819;
    wire n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827;
    wire n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835;
    wire n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843;
    wire n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851;
    wire n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859;
    wire n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867;
    wire n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875;
    wire n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883;
    wire n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891;
    wire n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899;
    wire n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907;
    wire n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915;
    wire n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923;
    wire n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931;
    wire n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939;
    wire n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947;
    wire n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955;
    wire n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963;
    wire n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971;
    wire n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979;
    wire n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987;
    wire n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995;
    wire n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003;
    wire n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011;
    wire n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019;
    wire n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027;
    wire n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035;
    wire n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043;
    wire n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051;
    wire n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059;
    wire n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067;
    wire n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075;
    wire n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083;
    wire n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091;
    wire n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099;
    wire n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107;
    wire n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115;
    wire n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123;
    wire n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131;
    wire n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139;
    wire n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147;
    wire n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155;
    wire n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163;
    wire n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171;
    wire n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179;
    wire n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187;
    wire n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195;
    wire n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203;
    wire n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211;
    wire n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219;
    wire n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227;
    wire n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235;
    wire n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243;
    wire n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251;
    wire n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259;
    wire n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267;
    wire n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275;
    wire n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283;
    wire n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291;
    wire n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299;
    wire n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307;
    wire n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315;
    wire n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323;
    wire n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331;
    wire n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339;
    wire n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347;
    wire n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355;
    wire n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363;
    wire n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371;
    wire n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379;
    wire n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387;
    wire n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395;
    wire n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403;
    wire n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411;
    wire n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419;
    wire n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427;
    wire n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435;
    wire n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443;
    wire n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451;
    wire n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459;
    wire n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467;
    wire n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475;
    wire n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483;
    wire n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491;
    wire n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499;
    wire n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507;
    wire n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515;
    wire n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523;
    wire n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531;
    wire n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539;
    wire n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547;
    wire n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555;
    wire n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563;
    wire n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571;
    wire n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579;
    wire n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587;
    wire n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595;
    wire n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603;
    wire n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611;
    wire n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619;
    wire n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627;
    wire n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635;
    wire n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643;
    wire n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651;
    wire n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659;
    wire n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667;
    wire n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675;
    wire n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683;
    wire n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691;
    wire n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699;
    wire n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707;
    wire n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715;
    wire n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723;
    wire n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731;
    wire n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739;
    wire n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747;
    wire n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755;
    wire n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763;
    wire n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771;
    wire n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779;
    wire n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787;
    wire n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795;
    wire n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803;
    wire n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811;
    wire n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819;
    wire n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827;
    wire n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835;
    wire n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843;
    wire n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851;
    wire n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859;
    wire n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867;
    wire n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875;
    wire n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883;
    wire n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891;
    wire n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899;
    wire n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907;
    wire n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915;
    wire n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923;
    wire n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931;
    wire n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939;
    wire n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947;
    wire n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955;
    wire n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963;
    wire n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971;
    wire n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979;
    wire n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987;
    wire n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995;
    wire n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003;
    wire n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011;
    wire n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019;
    wire n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027;
    wire n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035;
    wire n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043;
    wire n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051;
    wire n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059;
    wire n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067;
    wire n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075;
    wire n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083;
    wire n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091;
    wire n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099;
    wire n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107;
    wire n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115;
    wire n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123;
    wire n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131;
    wire n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139;
    wire n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147;
    wire n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155;
    wire n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163;
    wire n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171;
    wire n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179;
    wire n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187;
    wire n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195;
    wire n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203;
    wire n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211;
    wire n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219;
    wire n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227;
    wire n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235;
    wire n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243;
    wire n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251;
    wire n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259;
    wire n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267;
    wire n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275;
    wire n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283;
    wire n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291;
    wire n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299;
    wire n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307;
    wire n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315;
    wire n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323;
    wire n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331;
    wire n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339;
    wire n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347;
    wire n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355;
    wire n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363;
    wire n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371;
    wire n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379;
    wire n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387;
    wire n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395;
    wire n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403;
    wire n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411;
    wire n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419;
    wire n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427;
    wire n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435;
    wire n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443;
    wire n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451;
    wire n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459;
    wire n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467;
    wire n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475;
    wire n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483;
    wire n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491;
    wire n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499;
    wire n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507;
    wire n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515;
    wire n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523;
    wire n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531;
    wire n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539;
    wire n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547;
    wire n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555;
    wire n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563;
    wire n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571;
    wire n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579;
    wire n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587;
    wire n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595;
    wire n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603;
    wire n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611;
    wire n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619;
    wire n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627;
    wire n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635;
    wire n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643;
    wire n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651;
    wire n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659;
    wire n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667;
    wire n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675;
    wire n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683;
    wire n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691;
    wire n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699;
    wire n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707;
    wire n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715;
    wire n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723;
    wire n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731;
    wire n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739;
    wire n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747;
    wire n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755;
    wire n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763;
    wire n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771;
    wire n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779;
    wire n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787;
    wire n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795;
    wire n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803;
    wire n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811;
    wire n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819;
    wire n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827;
    wire n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835;
    wire n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843;
    wire n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851;
    wire n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859;
    wire n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867;
    wire n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875;
    wire n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883;
    wire n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891;
    wire n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899;
    wire n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907;
    wire n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915;
    wire n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923;
    wire n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931;
    wire n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939;
    wire n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947;
    wire n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955;
    wire n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963;
    wire n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971;
    wire n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979;
    wire n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987;
    wire n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995;
    wire n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003;
    wire n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011;
    wire n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019;
    wire n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027;
    wire n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035;
    wire n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043;
    wire n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051;
    wire n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059;
    wire n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067;
    wire n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075;
    wire n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083;
    wire n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091;
    wire n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099;
    wire n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107;
    wire n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115;
    wire n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123;
    wire n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131;
    wire n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139;
    wire n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147;
    wire n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155;
    wire n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163;
    wire n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171;
    wire n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179;
    wire n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187;
    wire n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195;
    wire n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203;
    wire n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211;
    wire n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219;
    wire n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227;
    wire n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235;
    wire n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243;
    wire n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251;
    wire n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259;
    wire n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267;
    wire n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275;
    wire n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283;
    wire n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291;
    wire n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299;
    wire n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307;
    wire n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315;
    wire n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323;
    wire n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331;
    wire n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339;
    wire n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347;
    wire n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355;
    wire n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363;
    wire n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371;
    wire n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379;
    wire n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387;
    wire n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395;
    wire n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403;
    wire n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411;
    wire n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419;
    wire n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427;
    wire n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435;
    wire n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443;
    wire n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451;
    wire n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459;
    wire n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467;
    wire n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475;
    wire n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483;
    wire n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491;
    wire n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499;
    wire n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507;
    wire n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515;
    wire n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523;
    wire n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531;
    wire n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539;
    wire n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547;
    wire n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555;
    wire n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563;
    wire n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571;
    wire n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579;
    wire n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587;
    wire n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595;
    wire n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603;
    wire n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611;
    wire n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619;
    wire n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627;
    wire n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635;
    wire n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643;
    wire n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651;
    wire n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659;
    wire n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667;
    wire n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675;
    wire n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683;
    wire n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691;
    wire n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699;
    wire n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707;
    wire n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715;
    wire n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723;
    wire n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731;
    wire n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739;
    wire n7740, n7741, n7742;
    not g0(n7377 ,n7379);
    not g1(n7376 ,n7382);
    not g2(n7375 ,n7698);
    not g3(n7374 ,n7731);
    not g4(n7373 ,n7730);
    not g5(n7372 ,n7396);
    not g6(n7371 ,n7381);
    not g7(n7370 ,n7729);
    not g8(n7369 ,n7394);
    not g9(n7368 ,n7390);
    not g10(n7367 ,n7728);
    not g11(n7366 ,n7707);
    not g12(n7365 ,n7380);
    not g13(n7364 ,n7727);
    not g14(n7363 ,n7389);
    not g15(n7362 ,n7726);
    not g16(n7361 ,n7699);
    not g17(n7360 ,n7725);
    not g18(n7359 ,n7724);
    not g19(n7358 ,n7378);
    not g20(n7357 ,n7723);
    not g21(n7356 ,n7393);
    not g22(n7355 ,n7388);
    not g23(n7354 ,n7708);
    not g24(n7353 ,n7722);
    not g25(n7352 ,n7742);
    not g26(n7351 ,n7721);
    not g27(n7350 ,n7720);
    not g28(n7349 ,n7741);
    not g29(n7348 ,n7719);
    not g30(n7347 ,n7387);
    not g31(n7346 ,n7718);
    not g32(n7345 ,n7709);
    not g33(n7344 ,n7740);
    not g34(n7343 ,n7716);
    not g35(n7342 ,n7395);
    not g36(n7341 ,n7739);
    not g37(n7340 ,n7715);
    not g38(n7339 ,n7392);
    not g39(n7338 ,n7386);
    not g40(n7337 ,n7714);
    not g41(n7336 ,n7738);
    not g42(n7335 ,n7713);
    not g43(n7334 ,n7737);
    not g44(n7333 ,n7711);
    not g45(n7332 ,n7385);
    not g46(n7331 ,n7710);
    not g47(n7330 ,n7736);
    not g48(n7329 ,n7717);
    not g49(n7328 ,n7712);
    not g50(n7327 ,n7735);
    not g51(n7326 ,n7391);
    not g52(n7325 ,n7384);
    not g53(n7324 ,n7706);
    not g54(n7323 ,n7734);
    not g55(n7322 ,n7705);
    not g56(n7321 ,n7704);
    not g57(n7320 ,n7733);
    not g58(n7319 ,n7703);
    not g59(n7318 ,n7383);
    not g60(n7317 ,n7702);
    not g61(n7316 ,n7732);
    not g62(n7315 ,n7701);
    not g63(n7314 ,n7700);
    not g64(n7313 ,n7401);
    not g65(n7312 ,n6);
    not g66(n7311 ,n7);
    or g67(n7528 ,n7262 ,n7310);
    or g68(n7557 ,n7260 ,n7289);
    or g69(n7554 ,n7268 ,n7302);
    or g70(n7548 ,n7274 ,n7306);
    or g71(n7535 ,n7276 ,n7308);
    or g72(n7547 ,n7270 ,n7305);
    or g73(n7534 ,n7273 ,n7307);
    or g74(n7533 ,n7271 ,n7304);
    or g75(n7546 ,n7266 ,n7299);
    or g76(n7532 ,n7269 ,n7303);
    or g77(n7531 ,n7267 ,n7301);
    or g78(n7530 ,n7256 ,n7298);
    or g79(n7553 ,n7277 ,n7291);
    or g80(n7545 ,n7263 ,n7279);
    or g81(n7529 ,n7264 ,n7296);
    or g82(n7558 ,n7265 ,n7297);
    or g83(n7536 ,n7246 ,n7309);
    or g84(n7527 ,n7261 ,n7293);
    or g85(n7552 ,n7258 ,n7287);
    or g86(n7543 ,n7259 ,n7290);
    or g87(n7556 ,n7252 ,n7280);
    or g88(n7551 ,n7254 ,n7286);
    or g89(n7542 ,n7257 ,n7288);
    or g90(n7541 ,n7255 ,n7285);
    or g91(n7540 ,n7253 ,n7284);
    or g92(n7539 ,n7251 ,n7283);
    or g93(n7555 ,n7275 ,n7300);
    or g94(n7550 ,n7250 ,n7282);
    or g95(n7538 ,n7249 ,n7281);
    or g96(n7549 ,n7247 ,n7295);
    or g97(n7537 ,n7248 ,n7294);
    or g98(n7544 ,n7272 ,n7292);
    nor g99(n7310 ,n7229 ,n7278);
    nor g100(n7309 ,n7183 ,n7278);
    nor g101(n7308 ,n7237 ,n7278);
    nor g102(n7307 ,n7177 ,n7278);
    nor g103(n7306 ,n7175 ,n7278);
    nor g104(n7305 ,n7226 ,n7278);
    nor g105(n7304 ,n7239 ,n7278);
    nor g106(n7303 ,n7230 ,n7278);
    nor g107(n7302 ,n7184 ,n7278);
    nor g108(n7301 ,n7225 ,n7278);
    nor g109(n7300 ,n7176 ,n7278);
    nor g110(n7299 ,n7215 ,n7278);
    nor g111(n7298 ,n7214 ,n7278);
    nor g112(n7297 ,n7191 ,n7278);
    nor g113(n7296 ,n7186 ,n7278);
    nor g114(n7295 ,n7212 ,n7278);
    nor g115(n7294 ,n7203 ,n7278);
    nor g116(n7293 ,n7178 ,n7278);
    nor g117(n7292 ,n7197 ,n7278);
    nor g118(n7291 ,n7223 ,n7278);
    nor g119(n7290 ,n7192 ,n7278);
    nor g120(n7289 ,n7202 ,n7278);
    nor g121(n7288 ,n7213 ,n7278);
    nor g122(n7287 ,n7210 ,n7278);
    nor g123(n7286 ,n7173 ,n7278);
    nor g124(n7285 ,n7228 ,n7278);
    nor g125(n7284 ,n7205 ,n7278);
    nor g126(n7283 ,n7227 ,n7278);
    nor g127(n7282 ,n7224 ,n7278);
    nor g128(n7281 ,n7233 ,n7278);
    nor g129(n7280 ,n7238 ,n7278);
    nor g130(n7279 ,n7174 ,n7278);
    not g131(n7662 ,n7278);
    nor g132(n7278 ,n7240 ,n7401);
    nor g133(n7277 ,n7181 ,n7171);
    nor g134(n7276 ,n7199 ,n7171);
    nor g135(n7275 ,n7198 ,n7171);
    nor g136(n7274 ,n7182 ,n7171);
    nor g137(n7273 ,n7180 ,n7171);
    nor g138(n7272 ,n7194 ,n7171);
    nor g139(n7271 ,n7236 ,n7171);
    nor g140(n7270 ,n7220 ,n7171);
    nor g141(n7269 ,n7231 ,n7171);
    nor g142(n7268 ,n7232 ,n7171);
    nor g143(n7267 ,n7217 ,n7171);
    nor g144(n7266 ,n7219 ,n7171);
    nor g145(n7265 ,n7189 ,n7171);
    nor g146(n7264 ,n7201 ,n7171);
    nor g147(n7263 ,n7185 ,n7171);
    nor g148(n7262 ,n7196 ,n7171);
    nor g149(n7261 ,n7209 ,n7171);
    nor g150(n7260 ,n7218 ,n7171);
    nor g151(n7259 ,n7187 ,n7171);
    nor g152(n7258 ,n7193 ,n7171);
    nor g153(n7257 ,n7190 ,n7171);
    nor g154(n7256 ,n7235 ,n7171);
    nor g155(n7255 ,n7179 ,n7171);
    nor g156(n7254 ,n7188 ,n7171);
    nor g157(n7253 ,n7204 ,n7171);
    nor g158(n7252 ,n7234 ,n7171);
    nor g159(n7251 ,n7195 ,n7171);
    nor g160(n7250 ,n7200 ,n7171);
    nor g161(n7249 ,n7221 ,n7171);
    nor g162(n7248 ,n7222 ,n7171);
    nor g163(n7247 ,n7211 ,n7171);
    nor g164(n7246 ,n7216 ,n7171);
    or g165(n7401 ,n7241 ,n7244);
    not g166(n7171 ,n7245);
    not g167(n7400 ,n7245);
    nor g168(n7245 ,n3[0] ,n7243);
    not g169(n7397 ,n7244);
    nor g170(n7244 ,n3[1] ,n7242);
    or g171(n7243 ,n7206 ,n7664);
    or g172(n7242 ,n7208 ,n7663);
    not g173(n7398 ,n7241);
    not g174(n7399 ,n7240);
    nor g175(n7241 ,n7663 ,n7664);
    nor g176(n7240 ,n7664 ,n7665);
    or g177(n7664 ,n7207 ,n3[2]);
    or g178(n7665 ,n3[3] ,n3[0]);
    or g179(n7663 ,n7172 ,n3[3]);
    not g180(n7239 ,n1[102]);
    not g181(n7238 ,n1[125]);
    not g182(n7237 ,n1[104]);
    not g183(n7236 ,n0[38]);
    not g184(n7235 ,n0[35]);
    not g185(n7234 ,n0[61]);
    not g186(n7233 ,n1[107]);
    not g187(n7232 ,n0[59]);
    not g188(n7231 ,n0[37]);
    not g189(n7230 ,n1[101]);
    not g190(n7229 ,n1[97]);
    not g191(n7228 ,n1[110]);
    not g192(n7227 ,n1[108]);
    not g193(n7226 ,n1[116]);
    not g194(n7225 ,n1[100]);
    not g195(n7224 ,n1[119]);
    not g196(n7223 ,n1[122]);
    not g197(n7222 ,n0[42]);
    not g198(n7221 ,n0[43]);
    not g199(n7220 ,n0[52]);
    not g200(n7219 ,n0[51]);
    not g201(n7218 ,n0[62]);
    not g202(n7217 ,n0[36]);
    not g203(n7216 ,n0[41]);
    not g204(n7215 ,n1[115]);
    not g205(n7214 ,n1[99]);
    not g206(n7213 ,n1[111]);
    not g207(n7212 ,n1[118]);
    not g208(n7211 ,n0[54]);
    not g209(n7210 ,n1[121]);
    not g210(n7209 ,n0[32]);
    not g211(n7208 ,n3[2]);
    not g212(n7207 ,n3[1]);
    not g213(n7206 ,n3[3]);
    not g214(n7205 ,n1[109]);
    not g215(n7204 ,n0[45]);
    not g216(n7203 ,n1[106]);
    not g217(n7202 ,n1[126]);
    not g218(n7201 ,n0[34]);
    not g219(n7200 ,n0[55]);
    not g220(n7199 ,n0[40]);
    not g221(n7198 ,n0[60]);
    not g222(n7197 ,n1[113]);
    not g223(n7196 ,n0[33]);
    not g224(n7195 ,n0[44]);
    not g225(n7194 ,n0[49]);
    not g226(n7193 ,n0[57]);
    not g227(n7192 ,n1[112]);
    not g228(n7191 ,n1[127]);
    not g229(n7190 ,n0[47]);
    not g230(n7189 ,n0[63]);
    not g231(n7188 ,n0[56]);
    not g232(n7187 ,n0[48]);
    not g233(n7186 ,n1[98]);
    not g234(n7185 ,n0[50]);
    not g235(n7184 ,n1[123]);
    not g236(n7183 ,n1[105]);
    not g237(n7182 ,n0[53]);
    not g238(n7181 ,n0[58]);
    not g239(n7180 ,n0[39]);
    not g240(n7179 ,n0[46]);
    not g241(n7178 ,n1[96]);
    not g242(n7177 ,n1[103]);
    not g243(n7176 ,n1[124]);
    not g244(n7175 ,n1[117]);
    not g245(n7174 ,n1[114]);
    not g246(n7173 ,n1[120]);
    not g247(n7172 ,n3[0]);
    or g248(n7622 ,n7004 ,n7169);
    or g249(n7589 ,n6985 ,n7119);
    or g250(n7587 ,n6995 ,n7125);
    or g251(n7584 ,n7002 ,n7135);
    or g252(n7577 ,n7013 ,n7139);
    or g253(n7595 ,n7014 ,n7141);
    or g254(n7594 ,n7042 ,n7140);
    or g255(n7562 ,n7011 ,n7122);
    or g256(n7593 ,n7010 ,n7137);
    or g257(n7592 ,n7009 ,n7136);
    or g258(n7576 ,n7007 ,n7133);
    or g259(n7561 ,n7008 ,n7134);
    or g260(n7560 ,n7006 ,n7132);
    or g261(n7583 ,n6997 ,n7129);
    or g262(n7575 ,n7003 ,n7130);
    or g263(n7623 ,n7005 ,n7154);
    or g264(n7591 ,n6989 ,n7127);
    or g265(n7574 ,n6999 ,n7128);
    or g266(n7621 ,n7001 ,n7168);
    or g267(n7620 ,n6998 ,n7167);
    or g268(n7582 ,n6990 ,n7124);
    or g269(n7573 ,n6992 ,n7126);
    or g270(n7619 ,n6994 ,n7166);
    or g271(n7618 ,n6993 ,n7165);
    or g272(n7572 ,n6987 ,n7123);
    or g273(n7617 ,n6991 ,n7164);
    or g274(n7616 ,n6988 ,n7163);
    or g275(n7581 ,n6980 ,n7121);
    or g276(n7571 ,n6981 ,n7138);
    or g277(n7615 ,n6986 ,n7162);
    or g278(n7614 ,n6983 ,n7161);
    or g279(n7613 ,n6952 ,n7160);
    or g280(n7604 ,n6966 ,n7151);
    or g281(n7590 ,n6954 ,n7109);
    or g282(n7586 ,n6976 ,n7118);
    or g283(n7580 ,n6996 ,n7115);
    or g284(n7570 ,n6978 ,n7120);
    or g285(n7611 ,n6977 ,n7158);
    or g286(n7610 ,n6975 ,n7157);
    or g287(n7569 ,n6973 ,n7117);
    or g288(n7609 ,n6974 ,n7156);
    or g289(n7608 ,n6972 ,n7155);
    or g290(n7579 ,n6962 ,n7113);
    or g291(n7568 ,n6969 ,n7116);
    or g292(n7607 ,n6970 ,n7170);
    or g293(n7606 ,n6968 ,n7153);
    or g294(n7567 ,n7000 ,n7114);
    or g295(n7605 ,n6967 ,n7152);
    or g296(n7612 ,n6979 ,n7159);
    or g297(n7588 ,n6982 ,n7131);
    or g298(n7585 ,n6961 ,n7111);
    or g299(n7566 ,n6957 ,n7112);
    or g300(n7603 ,n6965 ,n7150);
    or g301(n7602 ,n6963 ,n7149);
    or g302(n7565 ,n6958 ,n7110);
    or g303(n7601 ,n6960 ,n7148);
    or g304(n7600 ,n6959 ,n7147);
    or g305(n7578 ,n6955 ,n7108);
    or g306(n7564 ,n6964 ,n7107);
    or g307(n7599 ,n6956 ,n7146);
    or g308(n7598 ,n6953 ,n7145);
    or g309(n7563 ,n6984 ,n7142);
    or g310(n7597 ,n6951 ,n7144);
    or g311(n7596 ,n6971 ,n7143);
    not g312(n7714 ,n7170);
    not g313(n7699 ,n7169);
    not g314(n7700 ,n7168);
    not g315(n7701 ,n7167);
    not g316(n7702 ,n7166);
    not g317(n7703 ,n7165);
    not g318(n7704 ,n7164);
    not g319(n7705 ,n7163);
    not g320(n7706 ,n7162);
    not g321(n7707 ,n7161);
    not g322(n7708 ,n7160);
    not g323(n7709 ,n7159);
    not g324(n7710 ,n7158);
    not g325(n7711 ,n7157);
    not g326(n7712 ,n7156);
    not g327(n7713 ,n7155);
    not g328(n7698 ,n7154);
    not g329(n7715 ,n7153);
    not g330(n7716 ,n7152);
    not g331(n7717 ,n7151);
    not g332(n7718 ,n7150);
    not g333(n7719 ,n7149);
    not g334(n7720 ,n7148);
    not g335(n7721 ,n7147);
    not g336(n7722 ,n7146);
    not g337(n7723 ,n7145);
    not g338(n7724 ,n7144);
    not g339(n7725 ,n7143);
    not g340(n7393 ,n7142);
    not g341(n7726 ,n7141);
    not g342(n7727 ,n7140);
    not g343(n7379 ,n7139);
    nor g344(n7170 ,n7026 ,n7085);
    nor g345(n7169 ,n7041 ,n7100);
    nor g346(n7168 ,n7040 ,n7099);
    nor g347(n7167 ,n7039 ,n7098);
    nor g348(n7166 ,n7038 ,n7097);
    nor g349(n7165 ,n7037 ,n7096);
    nor g350(n7164 ,n7036 ,n7095);
    nor g351(n7163 ,n7035 ,n7094);
    nor g352(n7162 ,n7034 ,n7093);
    nor g353(n7161 ,n7033 ,n7092);
    nor g354(n7160 ,n7032 ,n7091);
    nor g355(n7159 ,n7031 ,n7090);
    nor g356(n7158 ,n7030 ,n7089);
    nor g357(n7157 ,n7029 ,n7088);
    nor g358(n7156 ,n7028 ,n7087);
    nor g359(n7155 ,n7027 ,n7102);
    nor g360(n7154 ,n7012 ,n7101);
    nor g361(n7153 ,n7025 ,n7084);
    nor g362(n7152 ,n7023 ,n7083);
    nor g363(n7151 ,n7022 ,n7082);
    nor g364(n7150 ,n7021 ,n7081);
    nor g365(n7149 ,n7020 ,n7080);
    nor g366(n7148 ,n7018 ,n7079);
    nor g367(n7147 ,n7017 ,n7078);
    nor g368(n7146 ,n7016 ,n7077);
    nor g369(n7145 ,n7019 ,n7076);
    nor g370(n7144 ,n7024 ,n7075);
    nor g371(n7143 ,n7015 ,n7086);
    nor g372(n7142 ,n6821 ,n7104);
    nor g373(n7141 ,n6821 ,n7105);
    nor g374(n7140 ,n6821 ,n7106);
    nor g375(n7139 ,n6821 ,n7058);
    not g376(n7385 ,n7138);
    not g377(n7728 ,n7137);
    not g378(n7729 ,n7136);
    not g379(n7737 ,n7135);
    not g380(n7395 ,n7134);
    not g381(n7380 ,n7133);
    not g382(n7396 ,n7132);
    not g383(n7733 ,n7131);
    not g384(n7381 ,n7130);
    not g385(n7738 ,n7129);
    not g386(n7382 ,n7128);
    not g387(n7730 ,n7127);
    not g388(n7383 ,n7126);
    not g389(n7734 ,n7125);
    not g390(n7739 ,n7124);
    not g391(n7384 ,n7123);
    not g392(n7394 ,n7122);
    not g393(n7740 ,n7121);
    not g394(n7386 ,n7120);
    not g395(n7732 ,n7119);
    not g396(n7735 ,n7118);
    not g397(n7387 ,n7117);
    not g398(n7388 ,n7116);
    not g399(n7741 ,n7115);
    not g400(n7389 ,n7114);
    not g401(n7742 ,n7113);
    not g402(n7390 ,n7112);
    not g403(n7736 ,n7111);
    not g404(n7391 ,n7110);
    not g405(n7731 ,n7109);
    not g406(n7378 ,n7108);
    not g407(n7392 ,n7107);
    nor g408(n7138 ,n6821 ,n7074);
    nor g409(n7137 ,n6821 ,n7073);
    nor g410(n7136 ,n6821 ,n7071);
    nor g411(n7135 ,n6821 ,n7068);
    nor g412(n7134 ,n6821 ,n7069);
    nor g413(n7133 ,n6821 ,n7067);
    nor g414(n7132 ,n6821 ,n7066);
    nor g415(n7131 ,n6821 ,n7070);
    nor g416(n7130 ,n6821 ,n7065);
    nor g417(n7129 ,n6821 ,n7064);
    nor g418(n7128 ,n6821 ,n7063);
    nor g419(n7127 ,n6821 ,n7057);
    nor g420(n7126 ,n6821 ,n7061);
    nor g421(n7125 ,n6821 ,n7062);
    nor g422(n7124 ,n6821 ,n7059);
    nor g423(n7123 ,n6820 ,n7060);
    nor g424(n7122 ,n6821 ,n7072);
    nor g425(n7121 ,n6821 ,n7056);
    nor g426(n7120 ,n6821 ,n7055);
    nor g427(n7119 ,n6821 ,n7054);
    nor g428(n7118 ,n6821 ,n7052);
    nor g429(n7117 ,n6820 ,n7053);
    nor g430(n7116 ,n6820 ,n7050);
    nor g431(n7115 ,n6821 ,n7051);
    nor g432(n7114 ,n6821 ,n7049);
    nor g433(n7113 ,n6821 ,n7048);
    nor g434(n7112 ,n6821 ,n7047);
    nor g435(n7111 ,n6821 ,n7045);
    nor g436(n7110 ,n6821 ,n7046);
    nor g437(n7109 ,n6821 ,n7103);
    nor g438(n7108 ,n6821 ,n7044);
    nor g439(n7107 ,n6820 ,n7043);
    not g440(n7626 ,n7106);
    not g441(n7627 ,n7105);
    not g442(n7669 ,n7104);
    not g443(n7696 ,n7103);
    or g444(n7102 ,n6820 ,n6931);
    or g445(n7101 ,n6820 ,n6945);
    or g446(n7100 ,n6820 ,n6944);
    or g447(n7099 ,n6820 ,n6943);
    or g448(n7098 ,n6820 ,n6942);
    or g449(n7097 ,n6820 ,n6926);
    or g450(n7096 ,n6820 ,n6941);
    or g451(n7095 ,n6820 ,n6940);
    or g452(n7094 ,n6820 ,n6950);
    or g453(n7093 ,n6820 ,n6938);
    or g454(n7092 ,n6820 ,n6937);
    or g455(n7091 ,n6820 ,n6936);
    or g456(n7090 ,n6820 ,n6934);
    or g457(n7089 ,n6820 ,n6925);
    or g458(n7088 ,n6820 ,n6933);
    or g459(n7087 ,n6820 ,n6932);
    or g460(n7086 ,n6820 ,n6948);
    or g461(n7085 ,n6820 ,n6924);
    or g462(n7084 ,n6820 ,n6929);
    or g463(n7083 ,n6820 ,n6928);
    or g464(n7082 ,n6820 ,n6947);
    or g465(n7081 ,n6820 ,n6923);
    or g466(n7080 ,n6820 ,n6935);
    or g467(n7079 ,n6820 ,n6939);
    or g468(n7078 ,n6820 ,n6949);
    or g469(n7077 ,n6820 ,n6946);
    or g470(n7076 ,n6820 ,n6927);
    or g471(n7075 ,n6820 ,n6930);
    xnor g472(n7106 ,n0[98] ,n0[66]);
    xnor g473(n7105 ,n0[99] ,n0[67]);
    xnor g474(n7104 ,n0[35] ,n0[3]);
    xnor g475(n7103 ,n0[62] ,n0[30]);
    not g476(n7677 ,n7074);
    not g477(n7625 ,n7073);
    not g478(n7668 ,n7072);
    not g479(n7624 ,n7071);
    not g480(n7694 ,n7070);
    not g481(n7667 ,n7069);
    not g482(n7690 ,n7068);
    not g483(n7682 ,n7067);
    not g484(n7666 ,n7066);
    not g485(n7681 ,n7065);
    not g486(n7689 ,n7064);
    not g487(n7680 ,n7063);
    not g488(n7693 ,n7062);
    not g489(n7679 ,n7061);
    not g490(n7678 ,n7060);
    not g491(n7688 ,n7059);
    not g492(n7683 ,n7058);
    not g493(n7697 ,n7057);
    not g494(n7687 ,n7056);
    not g495(n7676 ,n7055);
    not g496(n7695 ,n7054);
    not g497(n7675 ,n7053);
    not g498(n7692 ,n7052);
    not g499(n7686 ,n7051);
    not g500(n7674 ,n7050);
    not g501(n7673 ,n7049);
    not g502(n7685 ,n7048);
    not g503(n7672 ,n7047);
    not g504(n7671 ,n7046);
    not g505(n7691 ,n7045);
    not g506(n7684 ,n7044);
    not g507(n7670 ,n7043);
    xnor g508(n7074 ,n0[43] ,n0[11]);
    xnor g509(n7073 ,n0[97] ,n0[65]);
    xnor g510(n7072 ,n0[34] ,n0[2]);
    xnor g511(n7071 ,n0[96] ,n0[64]);
    xnor g512(n7070 ,n0[60] ,n0[28]);
    xnor g513(n7069 ,n0[33] ,n0[1]);
    xnor g514(n7068 ,n0[56] ,n0[24]);
    xnor g515(n7067 ,n0[48] ,n0[16]);
    xnor g516(n7066 ,n0[32] ,n0[0]);
    xnor g517(n7065 ,n0[47] ,n0[15]);
    xnor g518(n7064 ,n0[55] ,n0[23]);
    xnor g519(n7063 ,n0[46] ,n0[14]);
    xnor g520(n7062 ,n0[59] ,n0[27]);
    xnor g521(n7061 ,n0[45] ,n0[13]);
    xnor g522(n7060 ,n0[44] ,n0[12]);
    xnor g523(n7059 ,n0[54] ,n0[22]);
    xnor g524(n7058 ,n0[49] ,n0[17]);
    xnor g525(n7057 ,n0[63] ,n0[31]);
    xnor g526(n7056 ,n0[53] ,n0[21]);
    xnor g527(n7055 ,n0[42] ,n0[10]);
    xnor g528(n7054 ,n0[61] ,n0[29]);
    xnor g529(n7053 ,n0[41] ,n0[9]);
    xnor g530(n7052 ,n0[58] ,n0[26]);
    xnor g531(n7051 ,n0[52] ,n0[20]);
    xnor g532(n7050 ,n0[40] ,n0[8]);
    xnor g533(n7049 ,n0[39] ,n0[7]);
    xnor g534(n7048 ,n0[51] ,n0[19]);
    xnor g535(n7047 ,n0[38] ,n0[6]);
    xnor g536(n7046 ,n0[37] ,n0[5]);
    xnor g537(n7045 ,n0[57] ,n0[25]);
    xnor g538(n7044 ,n0[50] ,n0[18]);
    xnor g539(n7043 ,n0[36] ,n0[4]);
    nor g540(n7042 ,n6910 ,n6826);
    nor g541(n7041 ,n6896 ,n6838);
    nor g542(n7040 ,n6902 ,n6844);
    nor g543(n7039 ,n6908 ,n6887);
    nor g544(n7038 ,n6859 ,n6883);
    nor g545(n7037 ,n6852 ,n6890);
    nor g546(n7036 ,n6895 ,n6833);
    nor g547(n7035 ,n6847 ,n6886);
    nor g548(n7034 ,n6901 ,n6832);
    nor g549(n7033 ,n6855 ,n6880);
    nor g550(n7032 ,n6897 ,n6837);
    nor g551(n7031 ,n6906 ,n6881);
    nor g552(n7030 ,n6905 ,n6892);
    nor g553(n7029 ,n6851 ,n6839);
    nor g554(n7028 ,n6898 ,n6836);
    nor g555(n7027 ,n6848 ,n6894);
    nor g556(n7026 ,n6850 ,n6843);
    nor g557(n7025 ,n6853 ,n6893);
    nor g558(n7024 ,n6854 ,n6884);
    nor g559(n7023 ,n6900 ,n6835);
    nor g560(n7022 ,n6904 ,n6830);
    nor g561(n7021 ,n6899 ,n6891);
    nor g562(n7020 ,n6903 ,n6834);
    nor g563(n7019 ,n6907 ,n6882);
    nor g564(n7018 ,n6858 ,n6831);
    nor g565(n7017 ,n6857 ,n6840);
    nor g566(n7016 ,n6856 ,n6842);
    nor g567(n7015 ,n6846 ,n6845);
    nor g568(n7014 ,n6916 ,n6829);
    nor g569(n7013 ,n6836 ,n6822);
    nor g570(n7012 ,n6849 ,n6841);
    nor g571(n7011 ,n6879 ,n6828);
    nor g572(n7010 ,n6861 ,n6829);
    nor g573(n7009 ,n6917 ,n6827);
    nor g574(n7008 ,n6888 ,n6824);
    nor g575(n7007 ,n6894 ,n6822);
    nor g576(n7006 ,n6889 ,n6826);
    nor g577(n7005 ,n6860 ,n6823);
    nor g578(n7004 ,n6872 ,n6824);
    nor g579(n7003 ,n6843 ,n6823);
    nor g580(n7002 ,n6886 ,n6825);
    nor g581(n7001 ,n6909 ,n6824);
    nor g582(n7000 ,n6842 ,n6822);
    nor g583(n6999 ,n6893 ,n6828);
    nor g584(n6998 ,n6920 ,n6828);
    nor g585(n6997 ,n6832 ,n6827);
    nor g586(n6996 ,n6881 ,n6825);
    nor g587(n6995 ,n6883 ,n6827);
    nor g588(n6994 ,n6912 ,n6825);
    nor g589(n6993 ,n6873 ,n6826);
    nor g590(n6992 ,n6835 ,n6826);
    nor g591(n6991 ,n6877 ,n6826);
    nor g592(n6990 ,n6880 ,n6825);
    nor g593(n6989 ,n6841 ,n6828);
    nor g594(n6988 ,n6874 ,n6828);
    nor g595(n6987 ,n6830 ,n6824);
    nor g596(n6986 ,n6870 ,n6825);
    nor g597(n6985 ,n6844 ,n6823);
    nor g598(n6984 ,n6885 ,n6826);
    nor g599(n6983 ,n6922 ,n6824);
    nor g600(n6982 ,n6887 ,n6827);
    nor g601(n6981 ,n6891 ,n6829);
    nor g602(n6980 ,n6837 ,n6829);
    nor g603(n6979 ,n6919 ,n6828);
    nor g604(n6978 ,n6834 ,n6829);
    nor g605(n6977 ,n6915 ,n6822);
    nor g606(n6976 ,n6890 ,n6824);
    nor g607(n6975 ,n6864 ,n6823);
    nor g608(n6974 ,n6913 ,n6823);
    nor g609(n6973 ,n6831 ,n6823);
    nor g610(n6972 ,n6875 ,n6825);
    nor g611(n6971 ,n6869 ,n6826);
    nor g612(n6970 ,n6911 ,n6827);
    nor g613(n6969 ,n6840 ,n6822);
    nor g614(n6968 ,n6867 ,n6823);
    nor g615(n6967 ,n6876 ,n6822);
    nor g616(n6966 ,n6865 ,n6829);
    nor g617(n6965 ,n6862 ,n6828);
    nor g618(n6964 ,n6845 ,n6829);
    nor g619(n6963 ,n6918 ,n6824);
    nor g620(n6962 ,n6892 ,n6827);
    nor g621(n6961 ,n6833 ,n6825);
    nor g622(n6960 ,n6914 ,n6825);
    nor g623(n6959 ,n6866 ,n6824);
    nor g624(n6958 ,n6884 ,n6828);
    nor g625(n6957 ,n6882 ,n6822);
    nor g626(n6956 ,n6863 ,n6827);
    nor g627(n6955 ,n6839 ,n6827);
    nor g628(n6954 ,n6838 ,n6822);
    nor g629(n6953 ,n6868 ,n6823);
    nor g630(n6952 ,n6921 ,n6826);
    nor g631(n6951 ,n6871 ,n6829);
    nor g632(n6950 ,n0[120] ,n0[88]);
    nor g633(n6949 ,n0[104] ,n0[72]);
    nor g634(n6948 ,n0[100] ,n0[68]);
    nor g635(n6947 ,n0[108] ,n0[76]);
    nor g636(n6946 ,n0[103] ,n0[71]);
    nor g637(n6945 ,n0[127] ,n0[95]);
    nor g638(n6944 ,n0[126] ,n0[94]);
    nor g639(n6943 ,n0[125] ,n0[93]);
    nor g640(n6942 ,n0[124] ,n0[92]);
    nor g641(n6941 ,n0[122] ,n0[90]);
    nor g642(n6940 ,n0[121] ,n0[89]);
    nor g643(n6939 ,n0[105] ,n0[73]);
    nor g644(n6938 ,n0[119] ,n0[87]);
    nor g645(n6937 ,n0[118] ,n0[86]);
    nor g646(n6936 ,n0[117] ,n0[85]);
    nor g647(n6935 ,n0[106] ,n0[74]);
    nor g648(n6934 ,n0[116] ,n0[84]);
    nor g649(n6933 ,n0[114] ,n0[82]);
    nor g650(n6932 ,n0[113] ,n0[81]);
    nor g651(n6931 ,n0[112] ,n0[80]);
    nor g652(n6930 ,n0[101] ,n0[69]);
    nor g653(n6929 ,n0[110] ,n0[78]);
    nor g654(n6928 ,n0[109] ,n0[77]);
    nor g655(n6927 ,n0[102] ,n0[70]);
    nor g656(n6926 ,n0[123] ,n0[91]);
    nor g657(n6925 ,n0[115] ,n0[83]);
    nor g658(n6924 ,n0[111] ,n0[79]);
    nor g659(n6923 ,n0[107] ,n0[75]);
    not g660(n6922 ,n1[86]);
    not g661(n6921 ,n1[85]);
    not g662(n6920 ,n1[92]);
    not g663(n6919 ,n1[84]);
    not g664(n6918 ,n1[74]);
    not g665(n6917 ,n1[64]);
    not g666(n6916 ,n1[67]);
    not g667(n6915 ,n1[83]);
    not g668(n6914 ,n1[73]);
    not g669(n6913 ,n1[81]);
    not g670(n6912 ,n1[91]);
    not g671(n6911 ,n1[79]);
    not g672(n6910 ,n1[66]);
    not g673(n6909 ,n1[93]);
    not g674(n6908 ,n0[124]);
    not g675(n6907 ,n0[102]);
    not g676(n6906 ,n0[116]);
    not g677(n6905 ,n0[115]);
    not g678(n6904 ,n0[108]);
    not g679(n6903 ,n0[106]);
    not g680(n6902 ,n0[125]);
    not g681(n6901 ,n0[119]);
    not g682(n6900 ,n0[109]);
    not g683(n6899 ,n0[107]);
    not g684(n6898 ,n0[113]);
    not g685(n6897 ,n0[117]);
    not g686(n6896 ,n0[126]);
    not g687(n6895 ,n0[121]);
    not g688(n6894 ,n0[80]);
    not g689(n6893 ,n0[78]);
    not g690(n6892 ,n0[83]);
    not g691(n6891 ,n0[75]);
    not g692(n6890 ,n0[90]);
    not g693(n6889 ,n0[64]);
    not g694(n6888 ,n0[65]);
    not g695(n6887 ,n0[92]);
    not g696(n6886 ,n0[88]);
    not g697(n6885 ,n0[67]);
    not g698(n6884 ,n0[69]);
    not g699(n6883 ,n0[91]);
    not g700(n6882 ,n0[70]);
    not g701(n6881 ,n0[84]);
    not g702(n6880 ,n0[86]);
    not g703(n6879 ,n0[66]);
    not g704(n6821 ,n6878);
    not g705(n6820 ,n6878);
    not g706(n6878 ,n7400);
    not g707(n6877 ,n1[89]);
    not g708(n6876 ,n1[77]);
    not g709(n6875 ,n1[80]);
    not g710(n6874 ,n1[88]);
    not g711(n6873 ,n1[90]);
    not g712(n6872 ,n1[94]);
    not g713(n6871 ,n1[69]);
    not g714(n6870 ,n1[87]);
    not g715(n6869 ,n1[68]);
    not g716(n6868 ,n1[70]);
    not g717(n6867 ,n1[78]);
    not g718(n6866 ,n1[72]);
    not g719(n6865 ,n1[76]);
    not g720(n6864 ,n1[82]);
    not g721(n6863 ,n1[71]);
    not g722(n6862 ,n1[75]);
    not g723(n6861 ,n1[65]);
    not g724(n6860 ,n1[95]);
    not g725(n6859 ,n0[123]);
    not g726(n6858 ,n0[105]);
    not g727(n6857 ,n0[104]);
    not g728(n6856 ,n0[103]);
    not g729(n6855 ,n0[118]);
    not g730(n6854 ,n0[101]);
    not g731(n6853 ,n0[110]);
    not g732(n6852 ,n0[122]);
    not g733(n6851 ,n0[114]);
    not g734(n6850 ,n0[111]);
    not g735(n6849 ,n0[127]);
    not g736(n6848 ,n0[112]);
    not g737(n6847 ,n0[120]);
    not g738(n6846 ,n0[100]);
    not g739(n6845 ,n0[68]);
    not g740(n6844 ,n0[93]);
    not g741(n6843 ,n0[79]);
    not g742(n6842 ,n0[71]);
    not g743(n6841 ,n0[95]);
    not g744(n6840 ,n0[72]);
    not g745(n6839 ,n0[82]);
    not g746(n6838 ,n0[94]);
    not g747(n6837 ,n0[85]);
    not g748(n6836 ,n0[81]);
    not g749(n6835 ,n0[77]);
    not g750(n6834 ,n0[74]);
    not g751(n6833 ,n0[89]);
    not g752(n6832 ,n0[87]);
    not g753(n6831 ,n0[73]);
    not g754(n6830 ,n0[76]);
    not g755(n6829 ,n7662);
    not g756(n6828 ,n7662);
    not g757(n6827 ,n7662);
    not g758(n6826 ,n7662);
    not g759(n6825 ,n7662);
    not g760(n6824 ,n7662);
    not g761(n6823 ,n7662);
    not g762(n6822 ,n7662);
    or g763(n9[107] ,n5861 ,n6819);
    or g764(n9[96] ,n5492 ,n6818);
    or g765(n9[72] ,n6783 ,n6817);
    or g766(n9[67] ,n6782 ,n6815);
    or g767(n9[19] ,n6806 ,n6816);
    or g768(n9[0] ,n6803 ,n6814);
    or g769(n6819 ,n4941 ,n6813);
    or g770(n6818 ,n5348 ,n6812);
    or g771(n9[32] ,n5680 ,n6795);
    or g772(n9[73] ,n6047 ,n6796);
    or g773(n9[105] ,n5854 ,n6808);
    or g774(n9[104] ,n5851 ,n6807);
    or g775(n9[81] ,n6756 ,n6810);
    or g776(n9[112] ,n6786 ,n6802);
    or g777(n9[80] ,n6811 ,n6745);
    or g778(n6817 ,n5704 ,n6799);
    or g779(n6816 ,n5718 ,n6794);
    or g780(n6815 ,n5397 ,n6798);
    or g781(n9[65] ,n6596 ,n6809);
    or g782(n9[123] ,n6805 ,n6730);
    or g783(n9[115] ,n6787 ,n6800);
    or g784(n6814 ,n5400 ,n6804);
    or g785(n6813 ,n6731 ,n6797);
    or g786(n6812 ,n6741 ,n6801);
    or g787(n9[16] ,n6792 ,n6626);
    or g788(n6811 ,n5506 ,n6785);
    or g789(n9[120] ,n5850 ,n6771);
    or g790(n9[97] ,n5675 ,n6770);
    or g791(n9[9] ,n6748 ,n6778);
    or g792(n6810 ,n5714 ,n6777);
    or g793(n9[83] ,n6729 ,n6789);
    or g794(n9[75] ,n6521 ,n6784);
    or g795(n6809 ,n6719 ,n6775);
    or g796(n6808 ,n5158 ,n6773);
    or g797(n6807 ,n5042 ,n6772);
    or g798(n9[27] ,n6780 ,n6627);
    or g799(n6806 ,n5491 ,n6793);
    or g800(n6805 ,n5681 ,n6781);
    nor g801(n6804 ,n6768 ,n6693);
    or g802(n9[8] ,n6791 ,n6623);
    or g803(n9[91] ,n6725 ,n6790);
    or g804(n6803 ,n5672 ,n6788);
    nor g805(n6802 ,n1034 ,n6766);
    nor g806(n6801 ,n1038 ,n6762);
    nor g807(n6800 ,n1034 ,n6767);
    nor g808(n6799 ,n1036 ,n6765);
    nor g809(n6798 ,n1034 ,n6764);
    nor g810(n6797 ,n1034 ,n6763);
    or g811(n6796 ,n6707 ,n6776);
    or g812(n6795 ,n6703 ,n6774);
    nor g813(n6794 ,n6769 ,n6689);
    or g814(n9[11] ,n6779 ,n6625);
    nor g815(n6793 ,n1036 ,n6735);
    or g816(n9[56] ,n4423 ,n6754);
    or g817(n9[41] ,n4409 ,n6753);
    or g818(n9[33] ,n4911 ,n6752);
    or g819(n9[99] ,n5496 ,n6750);
    or g820(n9[24] ,n5846 ,n6751);
    or g821(n6792 ,n5674 ,n6749);
    or g822(n6791 ,n5488 ,n6747);
    or g823(n6790 ,n5375 ,n6746);
    or g824(n6789 ,n5508 ,n6757);
    nor g825(n6788 ,n1036 ,n6733);
    or g826(n6787 ,n6014 ,n6758);
    or g827(n9[88] ,n5864 ,n6724);
    or g828(n9[113] ,n6710 ,n6740);
    or g829(n6786 ,n6051 ,n6755);
    or g830(n6785 ,n5713 ,n6728);
    or g831(n6784 ,n6662 ,n6727);
    or g832(n6783 ,n5190 ,n6743);
    or g833(n6782 ,n5335 ,n6732);
    or g834(n6781 ,n5622 ,n6726);
    or g835(n6780 ,n6647 ,n6760);
    or g836(n6779 ,n6655 ,n6759);
    or g837(n6778 ,n5880 ,n6734);
    nor g838(n6777 ,n1038 ,n6723);
    nor g839(n6776 ,n1038 ,n6722);
    nor g840(n6775 ,n1036 ,n6721);
    nor g841(n6774 ,n1034 ,n6720);
    or g842(n6773 ,n6638 ,n6739);
    or g843(n6772 ,n6738 ,n6742);
    or g844(n6771 ,n6637 ,n6737);
    or g845(n6770 ,n6636 ,n6736);
    nor g846(n6769 ,n1047 ,n6744);
    nor g847(n6768 ,n1047 ,n6761);
    xnor g848(n6767 ,n6663 ,n2479);
    xnor g849(n6766 ,n6664 ,n1756);
    xnor g850(n6765 ,n6667 ,n2469);
    xnor g851(n6764 ,n6666 ,n2084);
    xnor g852(n6763 ,n6665 ,n1750);
    xnor g853(n6762 ,n6668 ,n2116);
    nor g854(n6761 ,n1038 ,n6692);
    or g855(n6760 ,n5847 ,n6699);
    or g856(n6759 ,n6034 ,n6688);
    nor g857(n6758 ,n6643 ,n6705);
    or g858(n6757 ,n5718 ,n6702);
    or g859(n6756 ,n5507 ,n6706);
    nor g860(n6755 ,n6634 ,n6704);
    or g861(n9[64] ,n5633 ,n6701);
    or g862(n9[57] ,n6589 ,n6718);
    or g863(n6754 ,n5159 ,n6717);
    or g864(n6753 ,n5156 ,n6716);
    or g865(n6752 ,n5155 ,n6714);
    or g866(n6751 ,n5154 ,n6698);
    or g867(n6750 ,n4936 ,n6700);
    or g868(n9[17] ,n6526 ,n6709);
    or g869(n6749 ,n5713 ,n6697);
    or g870(n6748 ,n5489 ,n6713);
    or g871(n6747 ,n5704 ,n6686);
    or g872(n9[3] ,n6525 ,n6708);
    or g873(n6746 ,n5615 ,n6685);
    nor g874(n6745 ,n1046 ,n1011);
    nor g875(n6744 ,n1038 ,n6696);
    or g876(n9[40] ,n5360 ,n6715);
    nor g877(n6743 ,n2365 ,n6677);
    nor g878(n6742 ,n1045 ,n6683);
    nor g879(n6741 ,n1045 ,n6680);
    nor g880(n6740 ,n1034 ,n6671);
    nor g881(n6739 ,n1038 ,n6675);
    nor g882(n6738 ,n1036 ,n6672);
    nor g883(n6737 ,n1034 ,n6676);
    nor g884(n6736 ,n1038 ,n6679);
    or g885(n6735 ,n6695 ,n6690);
    nor g886(n6734 ,n6687 ,n6575);
    or g887(n6733 ,n6691 ,n6694);
    nor g888(n6732 ,n1046 ,n6678);
    nor g889(n6731 ,n1046 ,n6684);
    nor g890(n6730 ,n2365 ,n6681);
    nor g891(n6729 ,n1038 ,n6670);
    nor g892(n6728 ,n1038 ,n6669);
    nor g893(n6727 ,n1034 ,n6674);
    nor g894(n6726 ,n1038 ,n6673);
    nor g895(n6725 ,n1038 ,n6682);
    nor g896(n6724 ,n6712 ,n6711);
    xnor g897(n6723 ,n2181 ,n1015);
    xnor g898(n6722 ,n1014 ,n2091);
    xnor g899(n6721 ,n6608 ,n2083);
    xnor g900(n6720 ,n2179 ,n1013);
    or g901(n9[122] ,n5865 ,n6654);
    or g902(n9[121] ,n5827 ,n6661);
    or g903(n6719 ,n5504 ,n6652);
    or g904(n6718 ,n5857 ,n6619);
    or g905(n6717 ,n5722 ,n6618);
    or g906(n9[43] ,n4913 ,n6649);
    or g907(n6716 ,n5712 ,n6617);
    or g908(n6715 ,n5720 ,n6616);
    or g909(n9[35] ,n4912 ,n6648);
    or g910(n6714 ,n5303 ,n6615);
    or g911(n9[98] ,n5495 ,n6646);
    or g912(n9[89] ,n5631 ,n6644);
    nor g913(n6713 ,n1038 ,n6641);
    nor g914(n6712 ,n4090 ,n6622);
    nor g915(n6711 ,n3940 ,n6639);
    or g916(n6710 ,n6053 ,n6653);
    or g917(n9[25] ,n6487 ,n6660);
    or g918(n6709 ,n6520 ,n6659);
    or g919(n6708 ,n6658 ,n6583);
    or g920(n9[1] ,n6657 ,n6635);
    nor g921(n6707 ,n2365 ,n6611);
    nor g922(n6706 ,n2365 ,n6610);
    or g923(n6705 ,n2365 ,n6621);
    or g924(n6704 ,n2365 ,n6633);
    nor g925(n6703 ,n2365 ,n6609);
    nor g926(n6702 ,n6642 ,n6620);
    nor g927(n6701 ,n6651 ,n6650);
    or g928(n6700 ,n6628 ,n6630);
    or g929(n6699 ,n5372 ,n6656);
    or g930(n6698 ,n6486 ,n6629);
    nor g931(n6697 ,n6632 ,n6614);
    not g932(n6696 ,n6695);
    not g933(n6694 ,n6693);
    not g934(n6692 ,n6691);
    not g935(n6690 ,n6689);
    or g936(n6688 ,n4935 ,n6645);
    nor g937(n6687 ,n1047 ,n6624);
    nor g938(n6686 ,n6631 ,n6613);
    nor g939(n6685 ,n6640 ,n6612);
    xnor g940(n6684 ,n6154 ,n6553);
    xnor g941(n6683 ,n6367 ,n6558);
    xnor g942(n6682 ,n3216 ,n6564);
    xnor g943(n6681 ,n6153 ,n6559);
    xnor g944(n6680 ,n6360 ,n6562);
    xnor g945(n6679 ,n6533 ,n2144);
    xnor g946(n6678 ,n6059 ,n6566);
    xnor g947(n6677 ,n6057 ,n6563);
    xnor g948(n6676 ,n3167 ,n6532);
    xnor g949(n6675 ,n6531 ,n2195);
    xnor g950(n6674 ,n6534 ,n2476);
    xnor g951(n6673 ,n6559 ,n3206);
    xnor g952(n6672 ,n6558 ,n3208);
    xnor g953(n6671 ,n6529 ,n2184);
    xnor g954(n6670 ,n3243 ,n6569);
    xnor g955(n6669 ,n3239 ,n6567);
    xnor g956(n6668 ,n6562 ,n2422);
    xnor g957(n6667 ,n2086 ,n6563);
    xnor g958(n6666 ,n2121 ,n6566);
    xnor g959(n6665 ,n6553 ,n2467);
    xnor g960(n6664 ,n6551 ,n2474);
    xnor g961(n6663 ,n6556 ,n1755);
    xnor g962(n6695 ,n6530 ,n2374);
    xnor g963(n6693 ,n6081 ,n6561);
    xnor g964(n6691 ,n6528 ,n2413);
    xnor g965(n6689 ,n6059 ,n6556);
    or g966(n6662 ,n4951 ,n6599);
    or g967(n9[74] ,n6300 ,n6598);
    or g968(n6661 ,n5705 ,n6580);
    or g969(n9[106] ,n5858 ,n6579);
    or g970(n9[51] ,n5126 ,n6606);
    or g971(n9[49] ,n4916 ,n6605);
    or g972(n9[48] ,n5122 ,n6604);
    or g973(n6660 ,n5824 ,n6549);
    or g974(n6659 ,n5490 ,n6595);
    or g975(n6658 ,n5376 ,n6593);
    or g976(n6657 ,n5486 ,n6591);
    or g977(n9[90] ,n6031 ,n6548);
    nor g978(n6656 ,n6159 ,n6560);
    nor g979(n6655 ,n6156 ,n6554);
    or g980(n6654 ,n4673 ,n6582);
    or g981(n9[82] ,n6191 ,n6600);
    nor g982(n6653 ,n6490 ,n6584);
    or g983(n9[66] ,n6189 ,n6597);
    or g984(n6652 ,n5453 ,n6601);
    nor g985(n6651 ,n4084 ,n6581);
    nor g986(n6650 ,n3936 ,n6590);
    or g987(n6649 ,n4938 ,n6603);
    or g988(n6648 ,n4937 ,n6602);
    nor g989(n6647 ,n6231 ,n6559);
    or g990(n6646 ,n4662 ,n6535);
    nor g991(n6645 ,n6233 ,n6553);
    or g992(n9[10] ,n6468 ,n6594);
    or g993(n9[2] ,n6186 ,n6592);
    or g994(n6644 ,n5431 ,n6547);
    nor g995(n6643 ,n6151 ,n6555);
    nor g996(n6642 ,n6157 ,n6568);
    or g997(n6641 ,n6573 ,n6574);
    nor g998(n6640 ,n6155 ,n6565);
    or g999(n6639 ,n6228 ,n6571);
    nor g1000(n6638 ,n1045 ,n6541);
    nor g1001(n6637 ,n2365 ,n6542);
    nor g1002(n6636 ,n2365 ,n6539);
    nor g1003(n6635 ,n2365 ,n6545);
    nor g1004(n6634 ,n6365 ,n6552);
    nor g1005(n6633 ,n6366 ,n6551);
    nor g1006(n6632 ,n6161 ,n6551);
    nor g1007(n6631 ,n6162 ,n6558);
    nor g1008(n6630 ,n1045 ,n6540);
    nor g1009(n6629 ,n1045 ,n6546);
    nor g1010(n6628 ,n1038 ,n6550);
    nor g1011(n6627 ,n1038 ,n6536);
    nor g1012(n6626 ,n1038 ,n6537);
    nor g1013(n6625 ,n1034 ,n6538);
    nor g1014(n6624 ,n1038 ,n6572);
    nor g1015(n6623 ,n1034 ,n6543);
    or g1016(n6622 ,n6162 ,n6570);
    nor g1017(n6621 ,n6152 ,n6556);
    nor g1018(n6620 ,n6229 ,n6569);
    or g1019(n6619 ,n5160 ,n6578);
    or g1020(n6618 ,n6588 ,n6577);
    or g1021(n6617 ,n6587 ,n6576);
    or g1022(n6616 ,n6585 ,n6607);
    or g1023(n6615 ,n6586 ,n6544);
    nor g1024(n6614 ,n6227 ,n6552);
    nor g1025(n6613 ,n6228 ,n6557);
    nor g1026(n6612 ,n6232 ,n6564);
    xnor g1027(n6611 ,n6080 ,n6496);
    xnor g1028(n6610 ,n6058 ,n6499);
    xnor g1029(n6609 ,n6495 ,n5978);
    xnor g1030(n6608 ,n2132 ,n6498);
    nor g1031(n6607 ,n6278 ,n6500);
    or g1032(n9[77] ,n6050 ,n6523);
    or g1033(n9[76] ,n6049 ,n6522);
    or g1034(n9[59] ,n5859 ,n6481);
    or g1035(n6606 ,n5721 ,n6480);
    or g1036(n6605 ,n5715 ,n6478);
    or g1037(n6604 ,n5707 ,n6477);
    or g1038(n6603 ,n5710 ,n6476);
    or g1039(n6602 ,n5394 ,n6475);
    nor g1040(n6601 ,n6234 ,n6498);
    or g1041(n9[114] ,n6467 ,n6494);
    or g1042(n6600 ,n6398 ,n6517);
    or g1043(n6599 ,n5879 ,n6527);
    or g1044(n6598 ,n6048 ,n6516);
    or g1045(n6597 ,n6396 ,n6515);
    nor g1046(n6596 ,n6160 ,n6497);
    or g1047(n6595 ,n5714 ,n6485);
    or g1048(n6594 ,n6033 ,n6489);
    or g1049(n6593 ,n5397 ,n6519);
    or g1050(n6592 ,n6386 ,n6484);
    or g1051(n6591 ,n5453 ,n6483);
    or g1052(n6590 ,n6227 ,n6503);
    nor g1053(n6589 ,n6298 ,n6511);
    nor g1054(n6588 ,n6308 ,n6509);
    nor g1055(n6587 ,n6281 ,n6506);
    nor g1056(n6586 ,n6276 ,n6505);
    nor g1057(n6585 ,n6279 ,n6501);
    or g1058(n6584 ,n2365 ,n6488);
    nor g1059(n6583 ,n1034 ,n6474);
    or g1060(n6582 ,n6382 ,n6493);
    or g1061(n6581 ,n6161 ,n6502);
    or g1062(n6580 ,n6513 ,n6479);
    or g1063(n6579 ,n6341 ,n6492);
    nor g1064(n6578 ,n6301 ,n6510);
    nor g1065(n6577 ,n6334 ,n6508);
    nor g1066(n6576 ,n6280 ,n6507);
    or g1067(n9[79] ,n6052 ,n6524);
    not g1068(n6575 ,n6574);
    not g1069(n6573 ,n6572);
    not g1070(n6571 ,n6570);
    not g1071(n6569 ,n6568);
    not g1072(n6565 ,n6564);
    not g1073(n6562 ,n6561);
    not g1074(n6560 ,n6559);
    not g1075(n6558 ,n6557);
    not g1076(n6555 ,n6556);
    not g1077(n6554 ,n6553);
    not g1078(n6551 ,n6552);
    xnor g1079(n6550 ,n6435 ,n3200);
    or g1080(n6549 ,n5431 ,n6518);
    or g1081(n6548 ,n6384 ,n6514);
    or g1082(n6547 ,n6512 ,n6482);
    xnor g1083(n6546 ,n6436 ,n6057);
    xnor g1084(n6545 ,n6427 ,n6058);
    nor g1085(n6544 ,n6275 ,n6504);
    xnor g1086(n6543 ,n6405 ,n2178);
    xnor g1087(n6542 ,n6436 ,n6149);
    xnor g1088(n6541 ,n6364 ,n6430);
    xnor g1089(n6540 ,n6150 ,n6435);
    xnor g1090(n6539 ,n6363 ,n6428);
    xnor g1091(n6538 ,n6403 ,n2197);
    xnor g1092(n6537 ,n6406 ,n2196);
    xnor g1093(n6536 ,n6404 ,n2194);
    or g1094(n6535 ,n6358 ,n6491);
    xnor g1095(n6574 ,n5969 ,n6429);
    xnor g1096(n6572 ,n6402 ,n2376);
    xnor g1097(n6534 ,n2087 ,n6438);
    xnor g1098(n6533 ,n6428 ,n1754);
    xnor g1099(n6532 ,n0[120] ,n6436);
    xnor g1100(n6531 ,n6430 ,n2475);
    xnor g1101(n6530 ,n6471 ,n1812);
    xnor g1102(n6529 ,n6431 ,n2437);
    xnor g1103(n6528 ,n6433 ,n2154);
    xnor g1104(n6570 ,n6149 ,n6472);
    xnor g1105(n6568 ,n6151 ,n6473);
    xnor g1106(n6567 ,n6366 ,n6437);
    xnor g1107(n6566 ,n6150 ,n6440);
    xnor g1108(n6564 ,n6153 ,n6471);
    xnor g1109(n6563 ,n6367 ,n6433);
    xnor g1110(n6561 ,n6433 ,n5978);
    xnor g1111(n6559 ,n5800 ,n6440);
    xnor g1112(n6557 ,n6071 ,n6437);
    xnor g1113(n6556 ,n6471 ,n5802);
    xnor g1114(n6553 ,n5797 ,n6473);
    xnor g1115(n6552 ,n6075 ,n6472);
    or g1116(n9[71] ,n6046 ,n6449);
    or g1117(n9[109] ,n5863 ,n6446);
    or g1118(n9[68] ,n6045 ,n6447);
    or g1119(n9[125] ,n5499 ,n6418);
    or g1120(n9[42] ,n4411 ,n6464);
    or g1121(n9[34] ,n4405 ,n6463);
    or g1122(n9[93] ,n5673 ,n6419);
    or g1123(n9[124] ,n5509 ,n6448);
    or g1124(n9[116] ,n5844 ,n6417);
    nor g1125(n6527 ,n6159 ,n6439);
    nor g1126(n6526 ,n6234 ,n6431);
    nor g1127(n6525 ,n6158 ,n6434);
    or g1128(n6524 ,n4127 ,n6453);
    or g1129(n6523 ,n4125 ,n6451);
    or g1130(n6522 ,n4124 ,n6450);
    nor g1131(n6521 ,n6231 ,n6438);
    or g1132(n9[69] ,n5823 ,n6466);
    or g1133(n9[58] ,n6345 ,n6465);
    or g1134(n9[102] ,n6122 ,n6469);
    or g1135(n9[26] ,n6188 ,n6462);
    or g1136(n9[18] ,n6187 ,n6461);
    nor g1137(n6520 ,n6160 ,n6432);
    or g1138(n9[95] ,n5825 ,n6460);
    nor g1139(n6519 ,n6230 ,n6435);
    nor g1140(n6518 ,n1045 ,n6413);
    nor g1141(n6517 ,n1036 ,n6408);
    nor g1142(n6516 ,n1038 ,n6410);
    nor g1143(n6515 ,n1036 ,n6414);
    nor g1144(n6514 ,n2364 ,n6426);
    nor g1145(n6513 ,n6356 ,n6442);
    nor g1146(n6512 ,n6271 ,n6444);
    not g1147(n6511 ,n6510);
    not g1148(n6509 ,n6508);
    not g1149(n6507 ,n6506);
    not g1150(n6505 ,n6504);
    not g1151(n6503 ,n6502);
    not g1152(n6501 ,n6500);
    not g1153(n6498 ,n6497);
    nor g1154(n6494 ,n1038 ,n6407);
    nor g1155(n6493 ,n1034 ,n6409);
    nor g1156(n6492 ,n1034 ,n6415);
    nor g1157(n6491 ,n1035 ,n6416);
    nor g1158(n6490 ,n6361 ,n6432);
    nor g1159(n6489 ,n6420 ,n6297);
    nor g1160(n6488 ,n6362 ,n6431);
    nor g1161(n6487 ,n1036 ,n1012);
    nor g1162(n6486 ,n1038 ,n6412);
    nor g1163(n6485 ,n1035 ,n6411);
    nor g1164(n6484 ,n2364 ,n6421);
    nor g1165(n6483 ,n1035 ,n6423);
    nor g1166(n6482 ,n6303 ,n6443);
    or g1167(n6481 ,n6459 ,n6445);
    or g1168(n6480 ,n6458 ,n6452);
    nor g1169(n6479 ,n6357 ,n6441);
    or g1170(n6478 ,n6454 ,n6470);
    or g1171(n6477 ,n6455 ,n6425);
    or g1172(n6476 ,n6457 ,n6424);
    or g1173(n6475 ,n6456 ,n6422);
    xnor g1174(n6474 ,n6338 ,n2157);
    xnor g1175(n6510 ,n5969 ,n6363);
    xnor g1176(n6508 ,n6060 ,n6360);
    xnor g1177(n6506 ,n6362 ,n6080);
    xnor g1178(n6504 ,n6078 ,n6364);
    xnor g1179(n6502 ,n6360 ,n6290);
    xnor g1180(n6500 ,n6057 ,n6365);
    xnor g1181(n6499 ,n6362 ,n6289);
    xnor g1182(n6497 ,n6363 ,n6288);
    xnor g1183(n6496 ,n6364 ,n6292);
    xnor g1184(n6495 ,n6072 ,n6367);
    nor g1185(n6470 ,n6285 ,n6381);
    or g1186(n6469 ,n4410 ,n6392);
    nor g1187(n6468 ,n2364 ,n6383);
    or g1188(n9[87] ,n6144 ,n6389);
    or g1189(n6467 ,n6055 ,n6385);
    or g1190(n9[85] ,n6107 ,n6400);
    or g1191(n9[84] ,n6142 ,n6399);
    or g1192(n9[70] ,n6133 ,n6397);
    or g1193(n6466 ,n6221 ,n6349);
    or g1194(n6465 ,n6044 ,n6355);
    or g1195(n9[103] ,n6123 ,n6394);
    or g1196(n6464 ,n4666 ,n6393);
    or g1197(n6463 ,n4664 ,n6391);
    or g1198(n6462 ,n6390 ,n6344);
    or g1199(n6461 ,n6401 ,n6343);
    or g1200(n6460 ,n6199 ,n6342);
    or g1201(n9[94] ,n6115 ,n6388);
    or g1202(n9[92] ,n6112 ,n6387);
    nor g1203(n6459 ,n6089 ,n6371);
    nor g1204(n6458 ,n6087 ,n6373);
    nor g1205(n6457 ,n6091 ,n6375);
    nor g1206(n6456 ,n6130 ,n6377);
    nor g1207(n6455 ,n6284 ,n6379);
    nor g1208(n6454 ,n6286 ,n6380);
    or g1209(n9[50] ,n4917 ,n6395);
    or g1210(n6453 ,n6139 ,n6353);
    nor g1211(n6452 ,n6086 ,n6372);
    or g1212(n6451 ,n6137 ,n6352);
    or g1213(n6450 ,n6136 ,n6351);
    or g1214(n6449 ,n6134 ,n6350);
    or g1215(n6448 ,n6141 ,n6346);
    or g1216(n6447 ,n6132 ,n6348);
    or g1217(n6446 ,n6131 ,n6347);
    nor g1218(n6445 ,n6088 ,n6370);
    nor g1219(n6473 ,n4920 ,n6369);
    nor g1220(n6472 ,n5023 ,n6368);
    nor g1221(n6471 ,n5143 ,n6369);
    not g1222(n6444 ,n6443);
    not g1223(n6442 ,n6441);
    not g1224(n6439 ,n6438);
    not g1225(n6434 ,n6435);
    not g1226(n6431 ,n6432);
    not g1227(n6430 ,n6429);
    not g1228(n6428 ,n6427);
    xnor g1229(n6426 ,n2149 ,n1010);
    nor g1230(n6425 ,n6283 ,n6378);
    nor g1231(n6424 ,n6111 ,n6374);
    xnor g1232(n6423 ,n6247 ,n3177);
    nor g1233(n6422 ,n6135 ,n6376);
    xnor g1234(n6421 ,n6237 ,n2090);
    nor g1235(n6420 ,n1047 ,n6359);
    or g1236(n6419 ,n6114 ,n6340);
    or g1237(n6418 ,n6116 ,n6339);
    or g1238(n6417 ,n6110 ,n6354);
    xnor g1239(n6416 ,n6248 ,n2402);
    xnor g1240(n6415 ,n6249 ,n2161);
    xnor g1241(n6414 ,n6239 ,n2066);
    xnor g1242(n6413 ,n6288 ,n6293);
    xnor g1243(n6412 ,n6245 ,n6235);
    xnor g1244(n6411 ,n6242 ,n6236);
    xnor g1245(n6410 ,n2182 ,n6243);
    xnor g1246(n6409 ,n6250 ,n2150);
    xnor g1247(n6408 ,n2172 ,n6246);
    xnor g1248(n6407 ,n6251 ,n1758);
    xnor g1249(n6406 ,n6241 ,n2385);
    xnor g1250(n6443 ,n6148 ,n6335);
    xnor g1251(n6441 ,n6067 ,n6288);
    xnor g1252(n6405 ,n6238 ,n2415);
    xnor g1253(n6404 ,n6244 ,n2375);
    xnor g1254(n6403 ,n6240 ,n2416);
    xnor g1255(n6402 ,n6289 ,n2193);
    nor g1256(n6440 ,n5354 ,n6369);
    xnor g1257(n6438 ,n6154 ,n6291);
    nor g1258(n6437 ,n5018 ,n6368);
    xnor g1259(n6436 ,n6290 ,n6065);
    xnor g1260(n6435 ,n5799 ,n6291);
    nor g1261(n6433 ,n5242 ,n6368);
    xnor g1262(n6432 ,n6068 ,n6335);
    xnor g1263(n6429 ,n6289 ,n6082);
    xnor g1264(n6427 ,n5960 ,n6292);
    or g1265(n6401 ,n5186 ,n6316);
    or g1266(n9[127] ,n4500 ,n6325);
    or g1267(n6400 ,n6054 ,n6302);
    or g1268(n6399 ,n4953 ,n6330);
    or g1269(n6398 ,n5192 ,n6329);
    or g1270(n9[111] ,n4493 ,n6327);
    or g1271(n6397 ,n4950 ,n6326);
    or g1272(n9[126] ,n5497 ,n6304);
    or g1273(n6396 ,n5505 ,n6299);
    or g1274(n6395 ,n5717 ,n6252);
    or g1275(n6394 ,n4725 ,n6324);
    or g1276(n6393 ,n5711 ,n6282);
    or g1277(n6392 ,n5724 ,n6323);
    or g1278(n9[101] ,n4479 ,n6322);
    or g1279(n9[100] ,n4719 ,n6320);
    or g1280(n6391 ,n5392 ,n6277);
    or g1281(n6390 ,n5187 ,n6319);
    or g1282(n9[23] ,n6018 ,n6318);
    or g1283(n6389 ,n6028 ,n6332);
    or g1284(n9[118] ,n5845 ,n6273);
    or g1285(n9[15] ,n6315 ,n6274);
    or g1286(n6388 ,n4711 ,n6313);
    or g1287(n6387 ,n4952 ,n6310);
    or g1288(n6386 ,n5487 ,n6272);
    or g1289(n9[86] ,n6108 ,n6331);
    nor g1290(n6385 ,n6170 ,n6307);
    or g1291(n9[78] ,n6104 ,n6328);
    or g1292(n9[36] ,n5761 ,n6321);
    or g1293(n9[21] ,n5738 ,n6317);
    or g1294(n9[13] ,n5754 ,n6314);
    or g1295(n9[117] ,n6305 ,n6333);
    or g1296(n9[6] ,n6093 ,n6312);
    or g1297(n9[5] ,n5769 ,n6311);
    nor g1298(n6384 ,n2365 ,n1009);
    or g1299(n6383 ,n6295 ,n6296);
    nor g1300(n6382 ,n2365 ,n6269);
    not g1301(n6381 ,n6380);
    not g1302(n6379 ,n6378);
    not g1303(n6377 ,n6376);
    not g1304(n6375 ,n6374);
    not g1305(n6373 ,n6372);
    not g1306(n6371 ,n6370);
    not g1307(n6365 ,n6366);
    not g1308(n6361 ,n6362);
    nor g1309(n6359 ,n1035 ,n6294);
    nor g1310(n6358 ,n1045 ,n6267);
    nor g1311(n6357 ,n3939 ,n6306);
    nor g1312(n6356 ,n4085 ,n6309);
    nor g1313(n6355 ,n1045 ,n6266);
    nor g1314(n6354 ,n2364 ,n6263);
    nor g1315(n6353 ,n1035 ,n6262);
    nor g1316(n6352 ,n1035 ,n6261);
    nor g1317(n6351 ,n1036 ,n6260);
    nor g1318(n6350 ,n1035 ,n6259);
    nor g1319(n6349 ,n1036 ,n6258);
    nor g1320(n6348 ,n1035 ,n6257);
    nor g1321(n6347 ,n1038 ,n6255);
    nor g1322(n6346 ,n2364 ,n6256);
    nor g1323(n6345 ,n1035 ,n6254);
    nor g1324(n6344 ,n1036 ,n6265);
    nor g1325(n6343 ,n1036 ,n6264);
    nor g1326(n6342 ,n1038 ,n6287);
    nor g1327(n6341 ,n2365 ,n6268);
    nor g1328(n6340 ,n2364 ,n6253);
    nor g1329(n6339 ,n1034 ,n6270);
    xnor g1330(n6380 ,n6148 ,n6058);
    xnor g1331(n6338 ,n6062 ,n6085);
    xnor g1332(n6378 ,n6149 ,n6081);
    xnor g1333(n6376 ,n6154 ,n6059);
    xnor g1334(n6374 ,n6152 ,n6077);
    xnor g1335(n6372 ,n6153 ,n6062);
    xnor g1336(n6370 ,n6150 ,n5959);
    nor g1337(n6369 ,n1029 ,n6291);
    nor g1338(n6368 ,n1029 ,n6290);
    nor g1339(n6367 ,n5017 ,n6337);
    nor g1340(n6366 ,n4645 ,n6337);
    nor g1341(n6364 ,n5125 ,n6336);
    nor g1342(n6363 ,n5120 ,n6336);
    nor g1343(n6362 ,n4523 ,n6336);
    nor g1344(n6360 ,n5243 ,n6337);
    nor g1345(n6334 ,n3930 ,n6164);
    or g1346(n9[119] ,n4906 ,n6202);
    or g1347(n6333 ,n4708 ,n6174);
    or g1348(n6332 ,n4892 ,n6146);
    or g1349(n6331 ,n5836 ,n6225);
    or g1350(n6330 ,n5874 ,n6106);
    or g1351(n6329 ,n5716 ,n6183);
    or g1352(n6328 ,n6224 ,n6138);
    or g1353(n6327 ,n3003 ,n6223);
    or g1354(n9[110] ,n5793 ,n6222);
    or g1355(n6326 ,n5882 ,n6103);
    or g1356(n6325 ,n3673 ,n6214);
    or g1357(n9[62] ,n5774 ,n6219);
    or g1358(n9[61] ,n5773 ,n6218);
    or g1359(n9[54] ,n5772 ,n6217);
    or g1360(n9[53] ,n5771 ,n6216);
    or g1361(n9[52] ,n5770 ,n6215);
    or g1362(n9[47] ,n5744 ,n6180);
    or g1363(n9[45] ,n5766 ,n6179);
    or g1364(n6324 ,n5723 ,n6102);
    or g1365(n9[39] ,n5743 ,n6178);
    or g1366(n6323 ,n3875 ,n6101);
    or g1367(n9[38] ,n6213 ,n6100);
    or g1368(n9[37] ,n6211 ,n6099);
    or g1369(n6322 ,n2680 ,n6212);
    or g1370(n6321 ,n6210 ,n5822);
    or g1371(n6320 ,n2723 ,n6209);
    or g1372(n9[31] ,n6208 ,n6098);
    or g1373(n9[30] ,n5759 ,n6207);
    or g1374(n9[29] ,n6206 ,n6118);
    or g1375(n9[28] ,n6205 ,n6097);
    or g1376(n6319 ,n5870 ,n6177);
    or g1377(n9[22] ,n5757 ,n6204);
    or g1378(n6318 ,n5871 ,n6117);
    or g1379(n6317 ,n6203 ,n5951);
    or g1380(n9[20] ,n5756 ,n6201);
    or g1381(n6316 ,n5716 ,n6176);
    or g1382(n6315 ,n5841 ,n6200);
    or g1383(n9[14] ,n5755 ,n6198);
    or g1384(n6314 ,n6197 ,n5829);
    or g1385(n9[12] ,n5753 ,n6196);
    or g1386(n6313 ,n5454 ,n6094);
    or g1387(n9[7] ,n5752 ,n6195);
    or g1388(n6312 ,n5831 ,n6194);
    or g1389(n6311 ,n6193 ,n5833);
    or g1390(n9[4] ,n5751 ,n6192);
    or g1391(n6310 ,n5457 ,n6092);
    nor g1392(n6309 ,n2366 ,n6147);
    or g1393(n9[63] ,n5502 ,n6220);
    nor g1394(n6308 ,n4078 ,n6126);
    or g1395(n6307 ,n2365 ,n6185);
    nor g1396(n6306 ,n2366 ,n6148);
    nor g1397(n6305 ,n1046 ,n6145);
    or g1398(n6304 ,n6105 ,n6128);
    nor g1399(n6303 ,n3931 ,n6109);
    or g1400(n6302 ,n4162 ,n6143);
    nor g1401(n6301 ,n4079 ,n6165);
    or g1402(n6300 ,n6190 ,n6182);
    or g1403(n6299 ,n4669 ,n6181);
    nor g1404(n6298 ,n3932 ,n6127);
    nor g1405(n6337 ,n1029 ,n6149);
    nor g1406(n6336 ,n1029 ,n6148);
    nor g1407(n6335 ,n5024 ,n6226);
    not g1408(n6297 ,n6296);
    not g1409(n6295 ,n6294);
    xnor g1410(n6287 ,n5902 ,n2136);
    nor g1411(n6286 ,n3926 ,n6125);
    nor g1412(n6285 ,n4074 ,n6163);
    nor g1413(n6284 ,n4072 ,n6124);
    nor g1414(n6283 ,n3924 ,n6166);
    or g1415(n6282 ,n6172 ,n6129);
    nor g1416(n6281 ,n3919 ,n6121);
    nor g1417(n6280 ,n4069 ,n6184);
    nor g1418(n6279 ,n4082 ,n6120);
    nor g1419(n6278 ,n3918 ,n6167);
    or g1420(n6277 ,n6171 ,n6140);
    nor g1421(n6276 ,n3915 ,n6119);
    nor g1422(n6275 ,n4066 ,n6168);
    or g1423(n6274 ,n5826 ,n6096);
    or g1424(n6273 ,n6095 ,n6113);
    or g1425(n6272 ,n4659 ,n6175);
    nor g1426(n6271 ,n4061 ,n6169);
    xnor g1427(n6270 ,n5885 ,n2128);
    xnor g1428(n6269 ,n5696 ,n5965);
    xnor g1429(n6268 ,n5690 ,n5963);
    xnor g1430(n6267 ,n5577 ,n5971);
    xnor g1431(n6266 ,n5693 ,n5976);
    xnor g1432(n6265 ,n5896 ,n5897);
    xnor g1433(n6264 ,n5898 ,n5899);
    xnor g1434(n6263 ,n1819 ,n5900);
    xnor g1435(n6262 ,n5895 ,n2125);
    xnor g1436(n6261 ,n5894 ,n2126);
    xnor g1437(n6260 ,n5893 ,n2127);
    xnor g1438(n6259 ,n5892 ,n2099);
    xnor g1439(n6258 ,n5891 ,n2078);
    xnor g1440(n6257 ,n5890 ,n2043);
    xnor g1441(n6256 ,n5888 ,n2108);
    xnor g1442(n6255 ,n5889 ,n2115);
    xnor g1443(n6254 ,n3219 ,n5976);
    xnor g1444(n6253 ,n5887 ,n2130);
    or g1445(n6252 ,n6173 ,n6090);
    xnor g1446(n6251 ,n5966 ,n2477);
    xnor g1447(n6250 ,n5965 ,n2478);
    xnor g1448(n6249 ,n5963 ,n2473);
    xnor g1449(n6248 ,n5971 ,n2120);
    xor g1450(n6247 ,n6058 ,n5960);
    xnor g1451(n6246 ,n2402 ,n5973);
    xor g1452(n6245 ,n6065 ,n0[8]);
    xnor g1453(n6244 ,n6077 ,n5800);
    xnor g1454(n6243 ,n2471 ,n5975);
    xnor g1455(n6296 ,n5578 ,n5962);
    xnor g1456(n6242 ,n0[1] ,n6068);
    xnor g1457(n6241 ,n6075 ,n6072);
    xnor g1458(n6294 ,n2371 ,n5901);
    xnor g1459(n6240 ,n5797 ,n5959);
    xnor g1460(n6239 ,n2110 ,n5980);
    xnor g1461(n6238 ,n6071 ,n6060);
    xnor g1462(n6237 ,n2152 ,n5886);
    xnor g1463(n6236 ,n6078 ,n3207);
    xor g1464(n6235 ,n6057 ,n3165);
    xnor g1465(n6293 ,n6067 ,n6080);
    nor g1466(n6292 ,n5076 ,n6226);
    xnor g1467(n6291 ,n5987 ,n4631);
    xnor g1468(n6290 ,n5988 ,n4875);
    nor g1469(n6289 ,n5019 ,n6226);
    nor g1470(n6288 ,n5665 ,n6226);
    not g1471(n6233 ,n6232);
    not g1472(n6230 ,n6229);
    or g1473(n6225 ,n5141 ,n6027);
    or g1474(n6224 ,n4510 ,n6026);
    or g1475(n6223 ,n5729 ,n5993);
    or g1476(n6222 ,n4740 ,n6025);
    or g1477(n6221 ,n4737 ,n6024);
    or g1478(n9[108] ,n5862 ,n5989);
    or g1479(n6220 ,n4288 ,n5990);
    or g1480(n6219 ,n5501 ,n5991);
    or g1481(n6218 ,n5500 ,n5992);
    or g1482(n6217 ,n5855 ,n6023);
    or g1483(n6216 ,n5853 ,n6022);
    or g1484(n6215 ,n5852 ,n5994);
    or g1485(n6214 ,n5396 ,n5995);
    or g1486(n9[46] ,n4483 ,n6021);
    or g1487(n6213 ,n5815 ,n6020);
    or g1488(n6212 ,n5726 ,n6000);
    or g1489(n6211 ,n5814 ,n6019);
    or g1490(n6210 ,n4444 ,n6039);
    or g1491(n6209 ,n5727 ,n6030);
    or g1492(n6208 ,n5679 ,n5913);
    or g1493(n6207 ,n5678 ,n5956);
    or g1494(n6206 ,n5677 ,n5955);
    or g1495(n6205 ,n5676 ,n5954);
    or g1496(n6204 ,n6038 ,n5953);
    or g1497(n6203 ,n4485 ,n6017);
    or g1498(n6202 ,n5728 ,n5948);
    or g1499(n6201 ,n6037 ,n5950);
    or g1500(n6200 ,n4466 ,n6016);
    or g1501(n6199 ,n4714 ,n6015);
    or g1502(n6198 ,n6036 ,n5947);
    or g1503(n6197 ,n4464 ,n6056);
    or g1504(n6196 ,n6035 ,n5946);
    or g1505(n6195 ,n6032 ,n5945);
    or g1506(n6194 ,n4577 ,n6013);
    or g1507(n6193 ,n4461 ,n6012);
    or g1508(n6192 ,n4902 ,n6011);
    nor g1509(n6191 ,n5811 ,n5973);
    nor g1510(n6190 ,n5809 ,n5975);
    nor g1511(n6189 ,n5806 ,n5980);
    nor g1512(n6188 ,n5809 ,n5965);
    nor g1513(n6187 ,n5806 ,n5966);
    nor g1514(n6186 ,n5811 ,n5971);
    nor g1515(n6185 ,n5686 ,n5966);
    nor g1516(n6184 ,n1046 ,n6083);
    nor g1517(n6183 ,n5807 ,n5972);
    nor g1518(n6182 ,n5808 ,n5974);
    nor g1519(n6181 ,n5810 ,n5979);
    or g1520(n9[55] ,n5418 ,n6043);
    or g1521(n6180 ,n6042 ,n5767);
    or g1522(n6179 ,n6041 ,n5817);
    or g1523(n6178 ,n6040 ,n5764);
    nor g1524(n6177 ,n5808 ,n5964);
    nor g1525(n6176 ,n5810 ,n5967);
    nor g1526(n6175 ,n5807 ,n5970);
    or g1527(n6174 ,n5620 ,n5943);
    nor g1528(n6173 ,n5996 ,n5982);
    nor g1529(n6172 ,n5998 ,n5984);
    nor g1530(n6171 ,n6005 ,n5986);
    nor g1531(n6170 ,n5685 ,n5967);
    nor g1532(n6169 ,n1046 ,n5968);
    nor g1533(n6168 ,n1045 ,n5961);
    nor g1534(n6167 ,n2365 ,n6070);
    nor g1535(n6166 ,n1046 ,n6074);
    nor g1536(n6165 ,n1046 ,n6066);
    nor g1537(n6164 ,n1046 ,n6065);
    nor g1538(n6163 ,n1045 ,n6069);
    or g1539(n6234 ,n1045 ,n6079);
    nor g1540(n6232 ,n2366 ,n5958);
    or g1541(n6231 ,n1045 ,n6076);
    nor g1542(n6229 ,n2366 ,n6063);
    nor g1543(n6228 ,n1045 ,n6061);
    nor g1544(n6227 ,n1045 ,n6073);
    nor g1545(n6226 ,n1029 ,n5911);
    not g1546(n6158 ,n6157);
    not g1547(n6156 ,n6155);
    not g1548(n6151 ,n6152);
    not g1549(n6147 ,n6148);
    nor g1550(n6146 ,n1034 ,n5905);
    nor g1551(n6145 ,n5944 ,n6007);
    nor g1552(n6144 ,n1046 ,n5931);
    nor g1553(n6143 ,n1045 ,n5930);
    nor g1554(n6142 ,n1045 ,n5929);
    nor g1555(n6141 ,n2365 ,n5926);
    nor g1556(n6140 ,n6006 ,n5985);
    nor g1557(n6139 ,n2365 ,n5928);
    nor g1558(n6138 ,n1045 ,n5927);
    nor g1559(n6137 ,n1045 ,n5914);
    nor g1560(n6136 ,n2365 ,n5925);
    nor g1561(n6135 ,n4062 ,n6008);
    nor g1562(n6134 ,n1045 ,n5957);
    nor g1563(n6133 ,n1046 ,n5924);
    nor g1564(n6132 ,n2365 ,n5923);
    nor g1565(n6131 ,n2365 ,n5921);
    nor g1566(n6130 ,n3917 ,n6001);
    nor g1567(n6129 ,n5999 ,n5983);
    nor g1568(n6128 ,n1045 ,n5922);
    nor g1569(n6127 ,n2365 ,n6067);
    nor g1570(n6126 ,n1045 ,n6064);
    nor g1571(n6125 ,n1045 ,n6068);
    nor g1572(n6124 ,n1045 ,n6075);
    nor g1573(n6123 ,n2365 ,n5920);
    nor g1574(n6122 ,n2365 ,n5933);
    nor g1575(n6121 ,n1045 ,n6082);
    nor g1576(n6120 ,n2365 ,n6071);
    nor g1577(n6119 ,n2365 ,n5960);
    nor g1578(n6118 ,n1045 ,n5940);
    nor g1579(n6117 ,n1046 ,n5912);
    nor g1580(n6116 ,n1045 ,n5932);
    nor g1581(n6115 ,n1045 ,n5919);
    nor g1582(n6114 ,n2366 ,n5917);
    nor g1583(n6113 ,n1045 ,n5918);
    nor g1584(n6112 ,n1046 ,n5916);
    nor g1585(n6111 ,n4070 ,n6009);
    nor g1586(n6110 ,n1046 ,n5915);
    nor g1587(n6109 ,n1046 ,n5969);
    nor g1588(n6108 ,n1036 ,n5906);
    nor g1589(n6107 ,n1036 ,n5907);
    nor g1590(n6106 ,n1036 ,n5908);
    nor g1591(n6105 ,n1035 ,n5904);
    nor g1592(n6104 ,n1036 ,n5909);
    nor g1593(n6103 ,n1034 ,n5910);
    nor g1594(n6102 ,n2364 ,n5934);
    nor g1595(n6101 ,n1038 ,n5903);
    nor g1596(n6100 ,n1035 ,n5935);
    nor g1597(n6099 ,n2364 ,n5936);
    nor g1598(n6098 ,n1035 ,n5937);
    nor g1599(n6097 ,n1036 ,n5938);
    nor g1600(n6096 ,n1035 ,n5939);
    nor g1601(n6095 ,n2364 ,n5941);
    nor g1602(n6094 ,n2364 ,n5942);
    nor g1603(n6093 ,n1035 ,n5949);
    nor g1604(n6092 ,n1038 ,n5952);
    nor g1605(n6091 ,n3921 ,n6002);
    nor g1606(n6090 ,n5997 ,n5981);
    nor g1607(n6089 ,n3933 ,n6004);
    nor g1608(n6088 ,n4080 ,n6010);
    nor g1609(n6087 ,n3928 ,n6003);
    nor g1610(n6086 ,n4076 ,n6029);
    nor g1611(n6162 ,n2366 ,n6060);
    nor g1612(n6161 ,n2365 ,n6072);
    or g1613(n6160 ,n2365 ,n6078);
    or g1614(n6159 ,n2365 ,n6077);
    nor g1615(n6157 ,n2366 ,n6062);
    xnor g1616(n6085 ,n5799 ,n2425);
    nor g1617(n6155 ,n1045 ,n5959);
    nor g1618(n6154 ,n4922 ,n6084);
    nor g1619(n6153 ,n5349 ,n6084);
    nor g1620(n6152 ,n4447 ,n6084);
    nor g1621(n6150 ,n4909 ,n6084);
    xnor g1622(n6149 ,n5813 ,n4877);
    xnor g1623(n6148 ,n5730 ,n5429);
    not g1624(n6083 ,n6082);
    not g1625(n6079 ,n6078);
    not g1626(n6076 ,n6077);
    not g1627(n6074 ,n6075);
    not g1628(n6073 ,n6072);
    not g1629(n6070 ,n6071);
    not g1630(n6069 ,n6068);
    not g1631(n6066 ,n6067);
    not g1632(n6065 ,n6064);
    not g1633(n6063 ,n6062);
    not g1634(n6061 ,n6060);
    or g1635(n6056 ,n4132 ,n5877);
    or g1636(n6055 ,n4497 ,n5835);
    or g1637(n6054 ,n4954 ,n5873);
    or g1638(n6053 ,n4496 ,n5834);
    or g1639(n6052 ,n4442 ,n5875);
    or g1640(n6051 ,n4495 ,n5832);
    or g1641(n6050 ,n4509 ,n5877);
    or g1642(n6049 ,n4508 ,n5878);
    or g1643(n6048 ,n4686 ,n5828);
    or g1644(n6047 ,n5191 ,n5880);
    or g1645(n6046 ,n4739 ,n5881);
    or g1646(n6045 ,n4735 ,n5884);
    or g1647(n9[60] ,n5407 ,n5860);
    or g1648(n6044 ,n4727 ,n5820);
    or g1649(n6043 ,n5856 ,n5728);
    or g1650(n6042 ,n4484 ,n5819);
    or g1651(n6041 ,n4724 ,n5818);
    or g1652(n9[44] ,n4915 ,n5848);
    or g1653(n6040 ,n4480 ,n5816);
    or g1654(n6039 ,n2560 ,n5821);
    or g1655(n6038 ,n4715 ,n5872);
    or g1656(n6037 ,n4468 ,n5874);
    or g1657(n6036 ,n4580 ,n5876);
    or g1658(n6035 ,n4713 ,n5878);
    or g1659(n6034 ,n4712 ,n5879);
    or g1660(n6033 ,n4903 ,n5830);
    or g1661(n6032 ,n4733 ,n5881);
    or g1662(n6031 ,n5185 ,n5870);
    or g1663(n6030 ,n5789 ,n5779);
    nor g1664(n6029 ,n2365 ,n5803);
    or g1665(n6028 ,n4164 ,n5871);
    or g1666(n6027 ,n5843 ,n5872);
    or g1667(n6026 ,n4126 ,n5876);
    or g1668(n6025 ,n5703 ,n5732);
    or g1669(n6024 ,n5883 ,n5842);
    or g1670(n6023 ,n4561 ,n5747);
    or g1671(n6022 ,n4272 ,n5746);
    or g1672(n6021 ,n3654 ,n5849);
    or g1673(n6020 ,n4721 ,n5763);
    or g1674(n6019 ,n4477 ,n5762);
    or g1675(n6018 ,n4582 ,n5740);
    or g1676(n6017 ,n4135 ,n5873);
    or g1677(n6016 ,n4133 ,n5875);
    or g1678(n6015 ,n5456 ,n5840);
    or g1679(n6014 ,n4498 ,n5837);
    or g1680(n6013 ,n5882 ,n5839);
    or g1681(n6012 ,n4130 ,n5883);
    or g1682(n6011 ,n5884 ,n5733);
    nor g1683(n6010 ,n2365 ,n5801);
    nor g1684(n6009 ,n1045 ,n5796);
    nor g1685(n6008 ,n2365 ,n5798);
    nor g1686(n6007 ,n4798 ,n5812);
    nor g1687(n6006 ,n4067 ,n5781);
    nor g1688(n6005 ,n3916 ,n5760);
    nor g1689(n6004 ,n2365 ,n5800);
    nor g1690(n6003 ,n2365 ,n5802);
    nor g1691(n6002 ,n2365 ,n5797);
    nor g1692(n6001 ,n1046 ,n5799);
    or g1693(n6000 ,n5790 ,n5778);
    nor g1694(n5999 ,n4064 ,n5838);
    nor g1695(n5998 ,n3920 ,n5765);
    nor g1696(n5997 ,n4075 ,n5782);
    nor g1697(n5996 ,n3927 ,n5768);
    or g1698(n5995 ,n5791 ,n5777);
    or g1699(n5994 ,n3819 ,n5745);
    or g1700(n5993 ,n5794 ,n5731);
    or g1701(n5992 ,n3838 ,n5748);
    or g1702(n5991 ,n3844 ,n5749);
    or g1703(n5990 ,n5750 ,n5775);
    or g1704(n5989 ,n5792 ,n5776);
    nor g1705(n5988 ,n1029 ,n5784);
    nor g1706(n5987 ,n1029 ,n5785);
    nor g1707(n6084 ,n1029 ,n5786);
    nor g1708(n6082 ,n5124 ,n5867);
    nor g1709(n6081 ,n5137 ,n5868);
    or g1710(n6080 ,n4520 ,n5869);
    nor g1711(n6078 ,n5132 ,n5869);
    nor g1712(n6077 ,n4438 ,n5804);
    nor g1713(n6075 ,n4887 ,n5866);
    nor g1714(n6072 ,n5130 ,n5868);
    nor g1715(n6071 ,n5121 ,n5866);
    nor g1716(n6068 ,n4522 ,n5867);
    nor g1717(n6067 ,n5129 ,n5867);
    nor g1718(n6064 ,n5016 ,n5866);
    nor g1719(n6062 ,n5140 ,n5804);
    nor g1720(n6060 ,n5026 ,n5868);
    nor g1721(n6059 ,n4924 ,n5804);
    or g1722(n6058 ,n5139 ,n5869);
    or g1723(n6057 ,n4525 ,n5868);
    not g1724(n5986 ,n5985);
    not g1725(n5984 ,n5983);
    not g1726(n5982 ,n5981);
    not g1727(n5980 ,n5979);
    not g1728(n5975 ,n5974);
    not g1729(n5973 ,n5972);
    not g1730(n5971 ,n5970);
    not g1731(n5968 ,n5969);
    not g1732(n5966 ,n5967);
    not g1733(n5965 ,n5964);
    not g1734(n5963 ,n5962);
    not g1735(n5961 ,n5960);
    not g1736(n5958 ,n5959);
    xnor g1737(n5957 ,n4956 ,n5603);
    or g1738(n5956 ,n4140 ,n5742);
    or g1739(n5955 ,n4139 ,n5741);
    or g1740(n5954 ,n4138 ,n5758);
    or g1741(n5953 ,n4136 ,n5739);
    xnor g1742(n5952 ,n3210 ,n5591);
    nor g1743(n5951 ,n5788 ,n5780);
    or g1744(n5950 ,n4134 ,n5737);
    xnor g1745(n5949 ,n5519 ,n2060);
    or g1746(n5948 ,n5787 ,n5783);
    or g1747(n5947 ,n4120 ,n5736);
    or g1748(n5946 ,n4131 ,n5735);
    or g1749(n5945 ,n4137 ,n5734);
    nor g1750(n5944 ,n4799 ,n5805);
    nor g1751(n5943 ,n5812 ,n5805);
    xnor g1752(n5942 ,n3181 ,n5580);
    xnor g1753(n5941 ,n3180 ,n5583);
    xnor g1754(n5940 ,n5572 ,n4957);
    xnor g1755(n5939 ,n5513 ,n1800);
    xnor g1756(n5938 ,n2137 ,n5518);
    xnor g1757(n5937 ,n1787 ,n5517);
    xnor g1758(n5936 ,n5516 ,n2134);
    xnor g1759(n5935 ,n5515 ,n2111);
    xnor g1760(n5934 ,n3204 ,n5581);
    xnor g1761(n5933 ,n4815 ,n5573);
    xnor g1762(n5932 ,n4802 ,n5572);
    xnor g1763(n5931 ,n4971 ,n5582);
    xnor g1764(n5930 ,n4966 ,n5594);
    xnor g1765(n5929 ,n4967 ,n5595);
    xnor g1766(n5928 ,n4975 ,n5596);
    xnor g1767(n5927 ,n4988 ,n5584);
    xnor g1768(n5926 ,n4968 ,n5600);
    xnor g1769(n5925 ,n4987 ,n5599);
    xnor g1770(n5924 ,n4976 ,n5604);
    xnor g1771(n5923 ,n4972 ,n5605);
    xnor g1772(n5922 ,n4969 ,n5593);
    xnor g1773(n5921 ,n4989 ,n5606);
    xnor g1774(n5920 ,n4814 ,n5581);
    xnor g1775(n5919 ,n4961 ,n5580);
    xnor g1776(n5918 ,n4797 ,n5583);
    xnor g1777(n5917 ,n4796 ,n5592);
    xnor g1778(n5916 ,n4800 ,n5591);
    xnor g1779(n5915 ,n4812 ,n5598);
    xnor g1780(n5914 ,n4957 ,n5597);
    or g1781(n5913 ,n4141 ,n5795);
    xnor g1782(n5912 ,n4956 ,n5601);
    xor g1783(n5911 ,n5514 ,n5426);
    xnor g1784(n5910 ,n3231 ,n5604);
    xnor g1785(n5909 ,n3238 ,n5584);
    xnor g1786(n5908 ,n3244 ,n5595);
    xnor g1787(n5907 ,n3246 ,n5594);
    xnor g1788(n5906 ,n3248 ,n5589);
    xnor g1789(n5905 ,n3249 ,n5582);
    xnor g1790(n5904 ,n3251 ,n5593);
    xnor g1791(n5903 ,n5573 ,n3202);
    xnor g1792(n5902 ,n2180 ,n5607);
    xnor g1793(n5901 ,n5687 ,n2198);
    xnor g1794(n5900 ,n2386 ,n5598);
    xnor g1795(n5899 ,n5694 ,n3170);
    xnor g1796(n5898 ,n0[2] ,n5689);
    xnor g1797(n5897 ,n5683 ,n3226);
    xnor g1798(n5896 ,n0[10] ,n5693);
    xnor g1799(n5895 ,n2031 ,n5596);
    xnor g1800(n5894 ,n2034 ,n5597);
    xnor g1801(n5893 ,n2033 ,n5599);
    xnor g1802(n5892 ,n2046 ,n5603);
    xnor g1803(n5891 ,n2122 ,n5587);
    xnor g1804(n5890 ,n2124 ,n5605);
    xnor g1805(n5889 ,n1796 ,n5606);
    xnor g1806(n5888 ,n2205 ,n5600);
    xnor g1807(n5887 ,n2188 ,n5592);
    xnor g1808(n5886 ,n5691 ,n5576);
    xnor g1809(n5985 ,n5690 ,n5694);
    xnor g1810(n5983 ,n5686 ,n5683);
    xnor g1811(n5981 ,n5696 ,n5691);
    xnor g1812(n5885 ,n5572 ,n2167);
    xnor g1813(n5979 ,n5577 ,n5699);
    nor g1814(n5978 ,n5117 ,n5866);
    xnor g1815(n5977 ,n5696 ,n5697);
    xnor g1816(n5976 ,n5577 ,n5578);
    xnor g1817(n5974 ,n5690 ,n5579);
    xnor g1818(n5972 ,n5686 ,n5687);
    xnor g1819(n5970 ,n5576 ,n5579);
    nor g1820(n5969 ,n5065 ,n5869);
    xnor g1821(n5967 ,n5689 ,n5697);
    xnor g1822(n5964 ,n5693 ,n5699);
    xnor g1823(n5962 ,n5687 ,n5700);
    nor g1824(n5960 ,n5119 ,n5867);
    nor g1825(n5959 ,n4901 ,n5804);
    or g1826(n5865 ,n4499 ,n5719);
    or g1827(n5864 ,n5485 ,n5725);
    or g1828(n5863 ,n4736 ,n5708);
    or g1829(n5862 ,n4949 ,n5709);
    or g1830(n5861 ,n4490 ,n5710);
    or g1831(n5860 ,n4730 ,n5664);
    or g1832(n5859 ,n5377 ,n5622);
    or g1833(n5858 ,n5188 ,n5711);
    or g1834(n5857 ,n4702 ,n5705);
    or g1835(n5856 ,n4704 ,n5522);
    or g1836(n5855 ,n4607 ,n5621);
    or g1837(n5854 ,n4488 ,n5712);
    or g1838(n5853 ,n4605 ,n5620);
    or g1839(n5852 ,n4573 ,n5702);
    or g1840(n5851 ,n4486 ,n5720);
    or g1841(n5850 ,n5498 ,n5722);
    or g1842(n5849 ,n5703 ,n5569);
    or g1843(n5848 ,n5709 ,n5568);
    or g1844(n5847 ,n4947 ,n5615);
    or g1845(n5846 ,n4907 ,n5725);
    or g1846(n5845 ,n4734 ,n5621);
    or g1847(n5844 ,n4945 ,n5702);
    nor g1848(n5843 ,n5094 ,n5590);
    nor g1849(n5842 ,n5090 ,n5588);
    nor g1850(n5841 ,n5105 ,n5586);
    nor g1851(n5840 ,n5105 ,n5608);
    nor g1852(n5839 ,n5094 ,n5574);
    or g1853(n10[18] ,n5064 ,n5634);
    or g1854(n10[19] ,n5179 ,n5635);
    or g1855(n10[20] ,n5177 ,n5636);
    or g1856(n10[21] ,n5176 ,n5637);
    or g1857(n10[22] ,n5174 ,n5639);
    nor g1858(n5838 ,n1046 ,n5701);
    or g1859(n10[8] ,n5127 ,n5669);
    or g1860(n10[7] ,n5022 ,n5668);
    or g1861(n10[6] ,n5015 ,n5667);
    or g1862(n10[5] ,n5021 ,n5666);
    or g1863(n10[4] ,n5025 ,n5659);
    or g1864(n5837 ,n4453 ,n5721);
    or g1865(n10[23] ,n5172 ,n5640);
    nor g1866(n5836 ,n5093 ,n5589);
    or g1867(n10[24] ,n5060 ,n5641);
    or g1868(n10[25] ,n5061 ,n5642);
    or g1869(n5835 ,n4220 ,n5717);
    or g1870(n10[26] ,n5063 ,n5643);
    or g1871(n5834 ,n4556 ,n5715);
    or g1872(n10[27] ,n5062 ,n5644);
    nor g1873(n5833 ,n5481 ,n5648);
    or g1874(n5832 ,n4671 ,n5707);
    nor g1875(n5831 ,n5093 ,n5573);
    or g1876(n5830 ,n4660 ,n5706);
    nor g1877(n5829 ,n5482 ,n5647);
    or g1878(n5828 ,n3910 ,n5706);
    or g1879(n5827 ,n4492 ,n5671);
    nor g1880(n5826 ,n5088 ,n5585);
    nor g1881(n5825 ,n5088 ,n5607);
    or g1882(n5824 ,n5670 ,n5494);
    nor g1883(n5823 ,n5111 ,n5587);
    nor g1884(n5822 ,n5483 ,n5646);
    or g1885(n5821 ,n3646 ,n5727);
    or g1886(n5820 ,n4668 ,n5719);
    or g1887(n5819 ,n3814 ,n5729);
    or g1888(n5818 ,n3809 ,n5708);
    nor g1889(n5817 ,n5464 ,n5645);
    or g1890(n5816 ,n3802 ,n5723);
    or g1891(n5815 ,n3801 ,n5724);
    or g1892(n5814 ,n3798 ,n5726);
    or g1893(n5884 ,n3859 ,n5663);
    or g1894(n5883 ,n3863 ,n5662);
    or g1895(n5882 ,n3866 ,n5661);
    or g1896(n5881 ,n3869 ,n5660);
    or g1897(n5880 ,n3874 ,n5658);
    or g1898(n5879 ,n3877 ,n5657);
    or g1899(n5878 ,n3881 ,n5656);
    or g1900(n5877 ,n3883 ,n5655);
    or g1901(n5876 ,n3884 ,n5654);
    or g1902(n5875 ,n3886 ,n5653);
    or g1903(n5874 ,n3896 ,n5652);
    or g1904(n5873 ,n3899 ,n5651);
    or g1905(n5872 ,n3902 ,n5650);
    or g1906(n5871 ,n3906 ,n5649);
    nor g1907(n5813 ,n1029 ,n5557);
    or g1908(n5870 ,n3782 ,n5561);
    nor g1909(n5869 ,n1029 ,n5546);
    nor g1910(n5868 ,n1029 ,n5547);
    nor g1911(n5867 ,n1029 ,n5552);
    nor g1912(n5866 ,n1029 ,n5559);
    not g1913(n5803 ,n5802);
    not g1914(n5801 ,n5800);
    not g1915(n5798 ,n5799);
    not g1916(n5796 ,n5797);
    nor g1917(n5795 ,n1046 ,n5525);
    or g1918(n10[16] ,n5074 ,n5632);
    or g1919(n10[15] ,n5134 ,n5630);
    or g1920(n10[14] ,n5138 ,n5629);
    or g1921(n10[13] ,n5071 ,n5628);
    or g1922(n10[12] ,n5069 ,n5627);
    or g1923(n10[11] ,n5142 ,n5626);
    or g1924(n10[10] ,n5135 ,n5625);
    or g1925(n10[9] ,n5114 ,n5638);
    nor g1926(n5794 ,n5333 ,n5586);
    nor g1927(n5793 ,n5330 ,n5624);
    nor g1928(n5792 ,n5318 ,n5612);
    nor g1929(n5791 ,n5324 ,n5614);
    nor g1930(n5790 ,n5357 ,n5617);
    nor g1931(n5789 ,n5363 ,n5619);
    nor g1932(n5788 ,n5089 ,n5610);
    nor g1933(n5787 ,n5244 ,n5602);
    xnor g1934(n5786 ,n5403 ,n5010);
    xor g1935(n5785 ,n5402 ,n4853);
    xnor g1936(n5784 ,n5401 ,n4850);
    nor g1937(n5783 ,n5240 ,n5601);
    nor g1938(n5782 ,n1045 ,n5688);
    nor g1939(n5781 ,n1045 ,n5575);
    nor g1940(n5780 ,n5110 ,n5609);
    nor g1941(n5779 ,n5370 ,n5618);
    nor g1942(n5778 ,n5358 ,n5616);
    nor g1943(n5777 ,n5322 ,n5613);
    nor g1944(n5776 ,n5316 ,n5611);
    nor g1945(n5775 ,n2366 ,n5537);
    nor g1946(n5774 ,n2366 ,n5536);
    nor g1947(n5773 ,n2366 ,n5535);
    nor g1948(n5772 ,n1046 ,n5534);
    nor g1949(n5771 ,n1046 ,n5533);
    nor g1950(n5770 ,n1046 ,n5532);
    nor g1951(n5769 ,n1046 ,n5541);
    nor g1952(n5768 ,n1046 ,n5689);
    nor g1953(n5767 ,n1045 ,n5531);
    nor g1954(n5766 ,n1046 ,n5530);
    nor g1955(n5765 ,n2365 ,n5700);
    nor g1956(n5764 ,n2365 ,n5529);
    nor g1957(n5763 ,n1045 ,n5528);
    nor g1958(n5762 ,n2365 ,n5527);
    nor g1959(n5761 ,n1046 ,n5526);
    nor g1960(n5760 ,n1045 ,n5576);
    or g1961(n10[17] ,n5131 ,n5682);
    nor g1962(n5759 ,n1045 ,n5524);
    nor g1963(n5758 ,n1045 ,n5523);
    nor g1964(n5757 ,n1045 ,n5571);
    nor g1965(n5756 ,n1046 ,n5521);
    nor g1966(n5755 ,n1046 ,n5520);
    nor g1967(n5754 ,n2366 ,n5538);
    nor g1968(n5753 ,n2366 ,n5539);
    nor g1969(n5752 ,n1045 ,n5540);
    nor g1970(n5751 ,n1045 ,n5542);
    nor g1971(n5750 ,n1036 ,n5549);
    nor g1972(n5749 ,n1034 ,n5550);
    nor g1973(n5748 ,n1034 ,n5551);
    nor g1974(n5747 ,n1035 ,n5553);
    nor g1975(n5746 ,n1035 ,n5554);
    nor g1976(n5745 ,n1034 ,n5555);
    nor g1977(n5744 ,n1038 ,n5556);
    nor g1978(n5743 ,n1034 ,n5558);
    nor g1979(n5742 ,n1036 ,n5560);
    nor g1980(n5741 ,n1034 ,n5543);
    nor g1981(n5740 ,n1034 ,n5544);
    nor g1982(n5739 ,n1034 ,n5562);
    nor g1983(n5738 ,n1036 ,n5545);
    nor g1984(n5737 ,n1038 ,n5563);
    nor g1985(n5736 ,n1034 ,n5564);
    nor g1986(n5735 ,n1036 ,n5565);
    nor g1987(n5734 ,n1038 ,n5566);
    nor g1988(n5733 ,n1038 ,n5567);
    nor g1989(n5732 ,n5326 ,n5623);
    nor g1990(n5731 ,n5331 ,n5585);
    nor g1991(n5812 ,n3911 ,n5610);
    or g1992(n5811 ,n2365 ,n5692);
    or g1993(n5810 ,n2365 ,n5694);
    or g1994(n5809 ,n2365 ,n5684);
    or g1995(n5808 ,n1046 ,n5683);
    or g1996(n5807 ,n1046 ,n5691);
    or g1997(n5806 ,n2366 ,n5695);
    nor g1998(n5805 ,n4065 ,n5609);
    nor g1999(n5730 ,n1029 ,n5548);
    nor g2000(n5804 ,n1029 ,n5570);
    nor g2001(n5802 ,n4446 ,n5698);
    nor g2002(n5800 ,n4914 ,n5698);
    nor g2003(n5799 ,n4910 ,n5698);
    nor g2004(n5797 ,n4921 ,n5698);
    not g2005(n5701 ,n5700);
    not g2006(n5695 ,n5694);
    not g2007(n5692 ,n5691);
    not g2008(n5688 ,n5689);
    not g2009(n5685 ,n5686);
    not g2010(n5684 ,n5683);
    or g2011(n5682 ,n5075 ,n5437);
    or g2012(n5681 ,n4427 ,n5406);
    or g2013(n5680 ,n5405 ,n5391);
    or g2014(n5679 ,n4475 ,n5456);
    or g2015(n5678 ,n4738 ,n5454);
    or g2016(n5677 ,n4717 ,n5458);
    or g2017(n5676 ,n4473 ,n5457);
    or g2018(n5675 ,n5493 ,n5303);
    or g2019(n5674 ,n4399 ,n5404);
    or g2020(n5673 ,n4946 ,n5458);
    or g2021(n5672 ,n4236 ,n5408);
    nor g2022(n5671 ,n1060 ,n5430);
    nor g2023(n5670 ,n1060 ,n5427);
    or g2024(n5669 ,n5115 ,n5452);
    or g2025(n5668 ,n5147 ,n5444);
    or g2026(n5667 ,n5146 ,n5443);
    or g2027(n5666 ,n5145 ,n5442);
    nor g2028(n5665 ,n1030 ,n5426);
    or g2029(n5664 ,n5425 ,n5416);
    or g2030(n5663 ,n5104 ,n5441);
    or g2031(n5662 ,n5106 ,n5442);
    or g2032(n5661 ,n5107 ,n5443);
    or g2033(n5660 ,n5108 ,n5444);
    or g2034(n5659 ,n5136 ,n5441);
    or g2035(n5658 ,n5203 ,n5451);
    or g2036(n5657 ,n5201 ,n5447);
    or g2037(n5656 ,n5200 ,n5446);
    or g2038(n5655 ,n5199 ,n5445);
    or g2039(n5654 ,n5198 ,n5440);
    or g2040(n5653 ,n5197 ,n5439);
    or g2041(n5652 ,n5193 ,n5434);
    or g2042(n5651 ,n5207 ,n5433);
    or g2043(n5650 ,n5206 ,n5432);
    or g2044(n5649 ,n5205 ,n5459);
    or g2045(n5648 ,n2364 ,n5423);
    or g2046(n5647 ,n2364 ,n5417);
    or g2047(n5646 ,n2364 ,n5422);
    or g2048(n5645 ,n2364 ,n5420);
    or g2049(n5644 ,n5169 ,n5450);
    or g2050(n5643 ,n5128 ,n5449);
    or g2051(n5642 ,n5170 ,n5431);
    or g2052(n5641 ,n5171 ,n5455);
    or g2053(n5640 ,n5173 ,n5459);
    or g2054(n5639 ,n5175 ,n5432);
    or g2055(n5638 ,n5066 ,n5451);
    or g2056(n5637 ,n5118 ,n5433);
    or g2057(n5636 ,n5178 ,n5434);
    or g2058(n5635 ,n5180 ,n5435);
    or g2059(n5634 ,n5014 ,n5436);
    or g2060(n5633 ,n5503 ,n5400);
    or g2061(n5632 ,n5073 ,n5438);
    or g2062(n5631 ,n5148 ,n5484);
    or g2063(n5630 ,n5123 ,n5439);
    or g2064(n5629 ,n5072 ,n5440);
    or g2065(n5628 ,n5070 ,n5445);
    or g2066(n5627 ,n5068 ,n5446);
    or g2067(n5626 ,n5116 ,n5447);
    or g2068(n5625 ,n5067 ,n5448);
    or g2069(n5729 ,n5378 ,n5476);
    or g2070(n5728 ,n5236 ,n5468);
    or g2071(n5727 ,n5362 ,n5415);
    or g2072(n5726 ,n5356 ,n5414);
    or g2073(n5725 ,n5102 ,n5455);
    or g2074(n5724 ,n5352 ,n5413);
    or g2075(n5723 ,n5336 ,n5412);
    or g2076(n5722 ,n5334 ,n5460);
    or g2077(n5721 ,n5342 ,n5480);
    or g2078(n5720 ,n5323 ,n5469);
    or g2079(n5719 ,n5341 ,n5463);
    or g2080(n5718 ,n5208 ,n5435);
    or g2081(n5717 ,n5340 ,n5479);
    or g2082(n5716 ,n5194 ,n5436);
    or g2083(n5715 ,n5339 ,n5478);
    or g2084(n5714 ,n5195 ,n5437);
    or g2085(n5713 ,n5196 ,n5438);
    or g2086(n5712 ,n5319 ,n5470);
    or g2087(n5711 ,n5311 ,n5471);
    or g2088(n5710 ,n5314 ,n5472);
    or g2089(n5709 ,n5321 ,n5473);
    or g2090(n5708 ,n5325 ,n5474);
    or g2091(n5707 ,n5337 ,n5477);
    or g2092(n5706 ,n5202 ,n5448);
    or g2093(n5705 ,n5327 ,n5462);
    or g2094(n5704 ,n5204 ,n5452);
    or g2095(n5703 ,n5328 ,n5475);
    or g2096(n5702 ,n5233 ,n5465);
    nor g2097(n5700 ,n4705 ,n5512);
    nor g2098(n5699 ,n4521 ,n5511);
    nor g2099(n5698 ,n1029 ,n5424);
    nor g2100(n5697 ,n4524 ,n5511);
    nor g2101(n5696 ,n4648 ,n5510);
    nor g2102(n5694 ,n4642 ,n5428);
    nor g2103(n5693 ,n4646 ,n5512);
    nor g2104(n5691 ,n4647 ,n5428);
    nor g2105(n5690 ,n4703 ,n5510);
    nor g2106(n5689 ,n3894 ,n5512);
    nor g2107(n5687 ,n4559 ,n5511);
    nor g2108(n5686 ,n3895 ,n5510);
    nor g2109(n5683 ,n3876 ,n5428);
    not g2110(n5624 ,n5623);
    not g2111(n5619 ,n5618);
    not g2112(n5617 ,n5616);
    not g2113(n5614 ,n5613);
    not g2114(n5612 ,n5611);
    not g2115(n5610 ,n5609);
    not g2116(n5608 ,n5607);
    not g2117(n5602 ,n5601);
    not g2118(n5590 ,n5589);
    not g2119(n5588 ,n5587);
    not g2120(n5586 ,n5585);
    not g2121(n5575 ,n5576);
    not g2122(n5574 ,n5573);
    xnor g2123(n5571 ,n5246 ,n5251);
    xnor g2124(n5570 ,n5211 ,n5013);
    or g2125(n5569 ,n5410 ,n5419);
    or g2126(n5568 ,n5411 ,n5421);
    xnor g2127(n5567 ,n3254 ,n5272);
    xnor g2128(n5566 ,n3199 ,n5275);
    xnor g2129(n5565 ,n3182 ,n5276);
    xnor g2130(n5564 ,n3184 ,n5249);
    xnor g2131(n5563 ,n3191 ,n5250);
    xnor g2132(n5562 ,n3193 ,n5251);
    or g2133(n5561 ,n5101 ,n5449);
    xnor g2134(n5560 ,n3201 ,n5253);
    xor g2135(n5559 ,n5212 ,n5213);
    xnor g2136(n5558 ,n3253 ,n5259);
    xor g2137(n5557 ,n5214 ,n5081);
    xnor g2138(n5556 ,n3209 ,n5261);
    xnor g2139(n5555 ,n3212 ,n5262);
    xnor g2140(n5554 ,n3213 ,n5263);
    xnor g2141(n5553 ,n3215 ,n5264);
    xor g2142(n5552 ,n5217 ,n5216);
    xnor g2143(n5551 ,n3221 ,n5267);
    xnor g2144(n5550 ,n3223 ,n5268);
    xnor g2145(n5549 ,n3225 ,n5269);
    xnor g2146(n5548 ,n5218 ,n4996);
    xor g2147(n5547 ,n5220 ,n5221);
    xor g2148(n5546 ,n5219 ,n5222);
    xnor g2149(n5545 ,n5227 ,n5225);
    xnor g2150(n5544 ,n5209 ,n5226);
    xnor g2151(n5543 ,n5210 ,n5223);
    xnor g2152(n5542 ,n5382 ,n5272);
    xnor g2153(n5541 ,n5386 ,n5273);
    xnor g2154(n5540 ,n5380 ,n5275);
    xnor g2155(n5539 ,n5387 ,n5276);
    xnor g2156(n5538 ,n5379 ,n5247);
    xnor g2157(n5537 ,n4977 ,n5269);
    xnor g2158(n5536 ,n4960 ,n5268);
    xnor g2159(n5535 ,n4808 ,n5267);
    xnor g2160(n5534 ,n4795 ,n5264);
    xnor g2161(n5533 ,n4801 ,n5263);
    xnor g2162(n5532 ,n4803 ,n5262);
    xnor g2163(n5531 ,n4982 ,n5261);
    xnor g2164(n5530 ,n4970 ,n5271);
    xnor g2165(n5529 ,n4816 ,n5259);
    xnor g2166(n5528 ,n4813 ,n5258);
    xnor g2167(n5527 ,n4809 ,n5257);
    xnor g2168(n5526 ,n4817 ,n5255);
    xnor g2169(n5525 ,n5384 ,n5254);
    xnor g2170(n5524 ,n5385 ,n5253);
    xnor g2171(n5523 ,n5383 ,n5252);
    or g2172(n5522 ,n3823 ,n5409);
    xnor g2173(n5521 ,n5388 ,n5250);
    xnor g2174(n5520 ,n5381 ,n5249);
    xnor g2175(n5623 ,n4978 ,n5381);
    or g2176(n5622 ,n5103 ,n5461);
    xnor g2177(n5519 ,n2190 ,n5228);
    or g2178(n5621 ,n5206 ,n5467);
    or g2179(n5620 ,n5207 ,n5466);
    xnor g2180(n5618 ,n4817 ,n5382);
    xnor g2181(n5616 ,n4809 ,n5386);
    or g2182(n5615 ,n5103 ,n5450);
    xnor g2183(n5518 ,n2073 ,n5252);
    xnor g2184(n5613 ,n4977 ,n5384);
    xnor g2185(n5517 ,n2068 ,n5254);
    xnor g2186(n5516 ,n1803 ,n5257);
    xnor g2187(n5515 ,n1813 ,n5258);
    xnor g2188(n5514 ,n5215 ,n4834);
    xnor g2189(n5513 ,n4789 ,n5224);
    xnor g2190(n5611 ,n4962 ,n5387);
    xnor g2191(n5609 ,n4801 ,n5265);
    xnor g2192(n5607 ,n4805 ,n5260);
    xnor g2193(n5606 ,n4970 ,n5379);
    xnor g2194(n5605 ,n4807 ,n5383);
    xnor g2195(n5604 ,n4815 ,n5385);
    xnor g2196(n5603 ,n4814 ,n5384);
    xnor g2197(n5601 ,n4793 ,n5260);
    xnor g2198(n5600 ,n4985 ,n5383);
    xnor g2199(n5599 ,n4965 ,n5382);
    xnor g2200(n5598 ,n4803 ,n5388);
    xnor g2201(n5597 ,n4989 ,n5386);
    xnor g2202(n5596 ,n4984 ,n5380);
    xnor g2203(n5595 ,n4812 ,n5387);
    xnor g2204(n5594 ,n4799 ,n5379);
    xnor g2205(n5593 ,n4960 ,n5385);
    xnor g2206(n5592 ,n4802 ,n5265);
    xnor g2207(n5591 ,n4968 ,n5388);
    xnor g2208(n5589 ,n4797 ,n5381);
    xnor g2209(n5587 ,n4811 ,n5266);
    xnor g2210(n5585 ,n4982 ,n5389);
    xnor g2211(n5584 ,n4981 ,n5390);
    xnor g2212(n5583 ,n4795 ,n5246);
    xnor g2213(n5582 ,n4792 ,n5389);
    xnor g2214(n5581 ,n4816 ,n5380);
    xnor g2215(n5580 ,n4969 ,n5246);
    nor g2216(n5579 ,n4564 ,n5511);
    nor g2217(n5578 ,n4575 ,n5428);
    nor g2218(n5577 ,n4584 ,n5510);
    nor g2219(n5576 ,n4583 ,n5512);
    xnor g2220(n5573 ,n4813 ,n5390);
    xnor g2221(n5572 ,n4808 ,n5266);
    or g2222(n5509 ,n4707 ,n5398);
    or g2223(n10[3] ,n4932 ,n5345);
    or g2224(n10[2] ,n4931 ,n5344);
    or g2225(n10[1] ,n4930 ,n5343);
    or g2226(n5508 ,n4511 ,n5369);
    or g2227(n5507 ,n4440 ,n5368);
    or g2228(n5506 ,n4439 ,n5367);
    or g2229(n5505 ,n5189 ,n5399);
    or g2230(n5504 ,n3532 ,n5365);
    or g2231(n5503 ,n4428 ,n5364);
    or g2232(n5502 ,n4491 ,n5396);
    or g2233(n5501 ,n4732 ,n5393);
    or g2234(n5500 ,n4731 ,n5395);
    or g2235(n5499 ,n4728 ,n5395);
    or g2236(n5498 ,n3602 ,n5361);
    or g2237(n5497 ,n4723 ,n5393);
    or g2238(n5496 ,n4474 ,n5394);
    or g2239(n5495 ,n4472 ,n5392);
    or g2240(n5494 ,n4585 ,n1016);
    or g2241(n5493 ,n5355 ,n4905);
    or g2242(n5492 ,n4487 ,n5391);
    or g2243(n5491 ,n4247 ,n5353);
    or g2244(n5490 ,n4243 ,n5351);
    or g2245(n5489 ,n4478 ,n5237);
    or g2246(n5488 ,n4240 ,n5350);
    or g2247(n5487 ,n5112 ,n5399);
    or g2248(n5486 ,n4458 ,n5235);
    or g2249(n10[28] ,n4897 ,n5234);
    or g2250(n5485 ,n4450 ,n5371);
    or g2251(n5484 ,n4456 ,n1016);
    nor g2252(n5483 ,n3433 ,n5256);
    nor g2253(n5482 ,n3415 ,n5248);
    nor g2254(n5481 ,n3411 ,n5274);
    nor g2255(n5480 ,n7313 ,n5307);
    nor g2256(n5479 ,n7313 ,n5304);
    nor g2257(n5478 ,n7313 ,n5305);
    nor g2258(n5477 ,n7313 ,n5300);
    nor g2259(n5476 ,n7313 ,n5297);
    nor g2260(n5475 ,n7313 ,n5296);
    nor g2261(n5474 ,n7313 ,n5294);
    nor g2262(n5473 ,n7313 ,n5293);
    nor g2263(n5472 ,n7313 ,n5292);
    nor g2264(n5471 ,n7313 ,n5291);
    nor g2265(n5470 ,n7313 ,n5290);
    nor g2266(n5469 ,n7313 ,n5289);
    nor g2267(n5468 ,n7313 ,n5282);
    nor g2268(n5467 ,n7313 ,n5281);
    nor g2269(n5466 ,n7313 ,n5280);
    nor g2270(n5465 ,n7313 ,n5277);
    nor g2271(n5464 ,n3447 ,n5270);
    nor g2272(n5463 ,n7313 ,n5306);
    nor g2273(n5462 ,n7313 ,n5295);
    nor g2274(n5461 ,n7313 ,n5288);
    nor g2275(n5460 ,n7313 ,n5286);
    nor g2276(n5512 ,n1029 ,n5231);
    nor g2277(n5511 ,n1029 ,n5230);
    nor g2278(n5510 ,n1029 ,n5232);
    not g2279(n5430 ,n5429);
    not g2280(n5427 ,n5426);
    nor g2281(n5425 ,n5313 ,n5302);
    xnor g2282(n5424 ,n5012 ,n5011);
    nor g2283(n5423 ,n3410 ,n5273);
    nor g2284(n5422 ,n3432 ,n5255);
    nor g2285(n5421 ,n5346 ,n5308);
    nor g2286(n5420 ,n3446 ,n5271);
    nor g2287(n5419 ,n5332 ,n5278);
    nor g2288(n5418 ,n5310 ,n5298);
    nor g2289(n5417 ,n3414 ,n5247);
    nor g2290(n5416 ,n5312 ,n5301);
    nor g2291(n5415 ,n7313 ,n5283);
    nor g2292(n5414 ,n7313 ,n5284);
    nor g2293(n5413 ,n7313 ,n5285);
    nor g2294(n5412 ,n7313 ,n5287);
    nor g2295(n5411 ,n5338 ,n5309);
    nor g2296(n5410 ,n5329 ,n5279);
    nor g2297(n5409 ,n5317 ,n5299);
    or g2298(n5408 ,n4457 ,n5347);
    or g2299(n5407 ,n3836 ,n5398);
    or g2300(n5406 ,n4190 ,n5373);
    or g2301(n5405 ,n3787 ,n5359);
    or g2302(n5404 ,n3727 ,n5241);
    nor g2303(n5459 ,n7398 ,n5282);
    or g2304(n5458 ,n3888 ,n5315);
    or g2305(n5457 ,n3856 ,n5245);
    or g2306(n5456 ,n3889 ,n5239);
    nor g2307(n5455 ,n7398 ,n5286);
    or g2308(n5454 ,n3858 ,n5238);
    or g2309(n5453 ,n3852 ,n5320);
    nor g2310(n5452 ,n7398 ,n5289);
    nor g2311(n5451 ,n7398 ,n5290);
    nor g2312(n5450 ,n7398 ,n5288);
    nor g2313(n5449 ,n7398 ,n5306);
    xnor g2314(n5403 ,n3946 ,n5084);
    nor g2315(n5448 ,n7398 ,n5291);
    nor g2316(n5447 ,n7398 ,n5292);
    nor g2317(n5446 ,n7398 ,n5293);
    nor g2318(n5445 ,n7398 ,n5294);
    xnor g2319(n5402 ,n5078 ,n4623);
    nor g2320(n5444 ,n7398 ,n5287);
    nor g2321(n5443 ,n7398 ,n5285);
    nor g2322(n5442 ,n7398 ,n5284);
    nor g2323(n5441 ,n7398 ,n5283);
    nor g2324(n5440 ,n7398 ,n5296);
    nor g2325(n5439 ,n7398 ,n5297);
    nor g2326(n5438 ,n7398 ,n5300);
    xnor g2327(n5401 ,n4868 ,n5077);
    nor g2328(n5437 ,n7398 ,n5305);
    nor g2329(n5436 ,n7398 ,n5304);
    nor g2330(n5435 ,n7398 ,n5307);
    nor g2331(n5434 ,n7398 ,n5277);
    nor g2332(n5433 ,n7398 ,n5280);
    nor g2333(n5432 ,n7398 ,n5281);
    nor g2334(n5431 ,n7398 ,n5295);
    nor g2335(n5429 ,n4693 ,n5366);
    nor g2336(n5428 ,n1029 ,n5229);
    nor g2337(n5426 ,n4606 ,n5374);
    or g2338(n5378 ,n3970 ,n5197);
    or g2339(n5377 ,n4729 ,n5020);
    or g2340(n5376 ,n4239 ,n5113);
    or g2341(n5375 ,n4393 ,n5165);
    nor g2342(n5374 ,n1025 ,n5099);
    nor g2343(n5373 ,n1060 ,n5085);
    nor g2344(n5372 ,n1060 ,n5079);
    or g2345(n5371 ,n4002 ,n5164);
    or g2346(n10[0] ,n5144 ,n5091);
    nor g2347(n5370 ,n4088 ,n5046);
    or g2348(n5369 ,n4214 ,n5163);
    or g2349(n5368 ,n4211 ,n5162);
    or g2350(n5367 ,n4210 ,n5044);
    nor g2351(n5366 ,n1022 ,n5099);
    or g2352(n5365 ,n4193 ,n5161);
    or g2353(n5364 ,n4192 ,n5043);
    nor g2354(n5363 ,n3914 ,n5028);
    or g2355(n5362 ,n3997 ,n5104);
    or g2356(n5361 ,n4185 ,n5157);
    or g2357(n5360 ,n5041 ,n4596);
    or g2358(n5359 ,n4147 ,n5040);
    nor g2359(n5358 ,n4068 ,n5047);
    nor g2360(n5357 ,n3913 ,n5029);
    or g2361(n5356 ,n3996 ,n5106);
    or g2362(n5355 ,n4174 ,n5153);
    nor g2363(n5354 ,n1028 ,n5079);
    or g2364(n5353 ,n4482 ,n5152);
    or g2365(n5352 ,n3993 ,n5107);
    or g2366(n5351 ,n4470 ,n5151);
    or g2367(n10[30] ,n5167 ,n5096);
    or g2368(n5350 ,n4463 ,n5038);
    nor g2369(n5349 ,n1030 ,n5085);
    or g2370(n10[31] ,n5166 ,n5092);
    or g2371(n10[29] ,n5168 ,n5098);
    nor g2372(n5348 ,n1058 ,n5081);
    nor g2373(n5347 ,n1057 ,n5077);
    nor g2374(n5346 ,n4089 ,n5048);
    or g2375(n5345 ,n4550 ,n5100);
    or g2376(n5344 ,n4549 ,n5097);
    or g2377(n5343 ,n4548 ,n5095);
    or g2378(n5342 ,n3980 ,n5208);
    or g2379(n5341 ,n3961 ,n5101);
    or g2380(n5340 ,n3963 ,n5194);
    or g2381(n5339 ,n3966 ,n5195);
    nor g2382(n5338 ,n3922 ,n5031);
    or g2383(n5337 ,n3969 ,n5196);
    or g2384(n5336 ,n3992 ,n5108);
    or g2385(n5335 ,n4430 ,n5133);
    or g2386(n5334 ,n3991 ,n5102);
    nor g2387(n5333 ,n3938 ,n5037);
    nor g2388(n5332 ,n4071 ,n5049);
    nor g2389(n5331 ,n4087 ,n5055);
    nor g2390(n5330 ,n3937 ,n5036);
    nor g2391(n5329 ,n3923 ,n5032);
    or g2392(n5328 ,n4001 ,n5198);
    or g2393(n5327 ,n3975 ,n5087);
    nor g2394(n5326 ,n4086 ,n5054);
    or g2395(n5325 ,n3976 ,n5199);
    nor g2396(n5324 ,n3925 ,n5030);
    or g2397(n5323 ,n3986 ,n5204);
    nor g2398(n5322 ,n4073 ,n5050);
    or g2399(n5321 ,n3978 ,n5200);
    or g2400(n5320 ,n4630 ,n5095);
    or g2401(n5319 ,n3985 ,n5203);
    nor g2402(n5318 ,n3935 ,n5035);
    nor g2403(n5317 ,n3929 ,n5033);
    nor g2404(n5316 ,n4083 ,n5053);
    or g2405(n5315 ,n4636 ,n5098);
    or g2406(n5314 ,n3981 ,n5201);
    nor g2407(n5313 ,n3934 ,n5034);
    nor g2408(n5312 ,n4081 ,n5052);
    or g2409(n5311 ,n3983 ,n5202);
    nor g2410(n5310 ,n4077 ,n5051);
    or g2411(n5400 ,n4634 ,n5091);
    or g2412(n5399 ,n3857 ,n5097);
    or g2413(n5398 ,n4891 ,n5059);
    or g2414(n5397 ,n4640 ,n5100);
    or g2415(n5396 ,n4783 ,n5058);
    or g2416(n5395 ,n4782 ,n5057);
    or g2417(n5394 ,n4764 ,n5184);
    or g2418(n5393 ,n4762 ,n5056);
    or g2419(n5392 ,n4759 ,n5183);
    or g2420(n5391 ,n4763 ,n5181);
    nor g2421(n5390 ,n2619 ,n5080);
    nor g2422(n5389 ,n2611 ,n5082);
    nor g2423(n5388 ,n2623 ,n5086);
    nor g2424(n5387 ,n2592 ,n5086);
    nor g2425(n5386 ,n2598 ,n5083);
    nor g2426(n5385 ,n2617 ,n5080);
    nor g2427(n5384 ,n2606 ,n5082);
    nor g2428(n5383 ,n2608 ,n5086);
    nor g2429(n5382 ,n2574 ,n5086);
    nor g2430(n5381 ,n2563 ,n5080);
    nor g2431(n5380 ,n2575 ,n5082);
    nor g2432(n5379 ,n2599 ,n5083);
    not g2433(n5309 ,n5308);
    not g2434(n5302 ,n5301);
    not g2435(n5299 ,n5298);
    not g2436(n5279 ,n5278);
    not g2437(n5274 ,n5273);
    not g2438(n5271 ,n5270);
    not g2439(n5256 ,n5255);
    not g2440(n5248 ,n5247);
    or g2441(n5245 ,n4635 ,n5109);
    nor g2442(n5244 ,n3912 ,n5027);
    nor g2443(n5243 ,n1030 ,n5081);
    nor g2444(n5242 ,n1026 ,n5077);
    or g2445(n5241 ,n3968 ,n5039);
    nor g2446(n5240 ,n4063 ,n5045);
    or g2447(n5239 ,n4637 ,n5092);
    or g2448(n5238 ,n4638 ,n5096);
    or g2449(n5237 ,n4110 ,n5150);
    or g2450(n5236 ,n3990 ,n5205);
    or g2451(n5235 ,n4108 ,n5149);
    or g2452(n5234 ,n4545 ,n5109);
    or g2453(n5233 ,n3982 ,n5193);
    xor g2454(n5232 ,n4751 ,n4752);
    xor g2455(n5231 ,n4757 ,n4756);
    xor g2456(n5230 ,n4754 ,n4755);
    xor g2457(n5229 ,n4758 ,n4753);
    xnor g2458(n5308 ,n4812 ,n4987);
    xnor g2459(n5228 ,n4958 ,n4813);
    xnor g2460(n5227 ,n0[5] ,n4801);
    xnor g2461(n5226 ,n4956 ,n3176);
    xnor g2462(n5225 ,n4973 ,n3211);
    xnor g2463(n5224 ,n4982 ,n2071);
    xnor g2464(n5223 ,n4957 ,n3205);
    xnor g2465(n5222 ,n4992 ,n5004);
    xnor g2466(n5221 ,n4990 ,n4512);
    xnor g2467(n5220 ,n5008 ,n4994);
    xnor g2468(n5219 ,n4864 ,n4334);
    xor g2469(n5307 ,n3355 ,n4830);
    xnor g2470(n5306 ,n3356 ,n1007);
    xor g2471(n5305 ,n3359 ,n4822);
    xor g2472(n5304 ,n3358 ,n4828);
    or g2473(n5303 ,n3994 ,n5182);
    xnor g2474(n5301 ,n4807 ,n4800);
    xor g2475(n5300 ,n3361 ,n4851);
    xnor g2476(n5298 ,n4805 ,n4971);
    xor g2477(n5297 ,n3363 ,n4857);
    xor g2478(n5296 ,n3364 ,n4859);
    xnor g2479(n5295 ,n3365 ,n1008);
    xor g2480(n5294 ,n3366 ,n4869);
    xnor g2481(n5218 ,n5000 ,n4327);
    xor g2482(n5293 ,n3367 ,n4820);
    xor g2483(n5292 ,n3369 ,n4824);
    xnor g2484(n5217 ,n4332 ,n5002);
    xnor g2485(n5216 ,n4998 ,n4866);
    xor g2486(n5291 ,n3370 ,n4826);
    xnor g2487(n5215 ,n4848 ,n4871);
    xor g2488(n5290 ,n3371 ,n4832);
    xor g2489(n5289 ,n3386 ,n4836);
    xnor g2490(n5288 ,n3368 ,n1005);
    xnor g2491(n5287 ,n3384 ,n4847);
    xnor g2492(n5286 ,n3374 ,n1006);
    xnor g2493(n5214 ,n4861 ,n4347);
    xnor g2494(n5285 ,n3375 ,n4846);
    xnor g2495(n5284 ,n3376 ,n4845);
    xnor g2496(n5213 ,n4873 ,n4818);
    xnor g2497(n5212 ,n4862 ,n4617);
    xnor g2498(n5283 ,n3377 ,n4842);
    xor g2499(n5282 ,n3382 ,n4840);
    xor g2500(n5281 ,n3362 ,n4843);
    xor g2501(n5280 ,n3360 ,n4855);
    xnor g2502(n5211 ,n5006 ,n4626);
    xnor g2503(n5278 ,n4797 ,n4988);
    xor g2504(n5277 ,n3379 ,n4838);
    xnor g2505(n5210 ,n0[13] ,n4808);
    xnor g2506(n5209 ,n0[7] ,n4793);
    xnor g2507(n5276 ,n4800 ,n4962);
    xnor g2508(n5275 ,n4971 ,n4816);
    xnor g2509(n5273 ,n4966 ,n4809);
    xnor g2510(n5272 ,n4967 ,n4817);
    xnor g2511(n5270 ,n4957 ,n4798);
    xnor g2512(n5269 ,n4814 ,n4789);
    xnor g2513(n5268 ,n4815 ,n4961);
    xnor g2514(n5267 ,n4811 ,n4796);
    nor g2515(n5266 ,n2603 ,n5083);
    nor g2516(n5265 ,n2590 ,n5083);
    xnor g2517(n5264 ,n4969 ,n4958);
    xnor g2518(n5263 ,n4802 ,n4966);
    xnor g2519(n5262 ,n4968 ,n4967);
    xnor g2520(n5261 ,n4792 ,n4975);
    nor g2521(n5260 ,n2582 ,n5082);
    xnor g2522(n5259 ,n4984 ,n4956);
    xnor g2523(n5258 ,n4981 ,n4976);
    xnor g2524(n5257 ,n4989 ,n4973);
    xnor g2525(n5255 ,n4965 ,n4972);
    xnor g2526(n5254 ,n4975 ,n4977);
    xnor g2527(n5253 ,n4988 ,n4960);
    xnor g2528(n5252 ,n4987 ,n4985);
    xnor g2529(n5251 ,n4795 ,n4976);
    xnor g2530(n5250 ,n4803 ,n4972);
    xnor g2531(n5249 ,n4961 ,n4978);
    xnor g2532(n5247 ,n4796 ,n4970);
    nor g2533(n5246 ,n2613 ,n5080);
    or g2534(n5192 ,n4928 ,n4441);
    or g2535(n5191 ,n3558 ,n4927);
    or g2536(n5190 ,n4926 ,n4436);
    or g2537(n5189 ,n3535 ,n4923);
    or g2538(n5188 ,n3511 ,n4919);
    or g2539(n5187 ,n4471 ,n4760);
    or g2540(n5186 ,n4244 ,n4904);
    or g2541(n5185 ,n3259 ,n4896);
    nor g2542(n5184 ,n7313 ,n4886);
    nor g2543(n5183 ,n7313 ,n4882);
    nor g2544(n5182 ,n7313 ,n4880);
    nor g2545(n5181 ,n7313 ,n4881);
    or g2546(n5180 ,n1691 ,n4772);
    nor g2547(n5179 ,n1061 ,n4831);
    or g2548(n5178 ,n1714 ,n4771);
    nor g2549(n5177 ,n1061 ,n4839);
    nor g2550(n5176 ,n1061 ,n4856);
    or g2551(n5175 ,n1695 ,n4770);
    nor g2552(n5174 ,n1061 ,n4844);
    or g2553(n5173 ,n1643 ,n4769);
    nor g2554(n5172 ,n1061 ,n4841);
    or g2555(n5171 ,n1622 ,n4768);
    or g2556(n5170 ,n1667 ,n4767);
    or g2557(n5169 ,n1709 ,n4765);
    or g2558(n5168 ,n4576 ,n4898);
    or g2559(n5167 ,n4656 ,n4899);
    or g2560(n5166 ,n4594 ,n4900);
    or g2561(n5165 ,n4199 ,n4933);
    nor g2562(n5164 ,n1060 ,n4995);
    nor g2563(n5163 ,n1060 ,n5007);
    nor g2564(n5162 ,n1057 ,n4993);
    nor g2565(n5161 ,n1060 ,n5005);
    nor g2566(n5160 ,n1058 ,n5003);
    nor g2567(n5159 ,n1060 ,n4863);
    nor g2568(n5158 ,n1058 ,n5001);
    nor g2569(n5157 ,n1057 ,n4878);
    nor g2570(n5156 ,n1057 ,n4999);
    nor g2571(n5155 ,n1060 ,n4867);
    nor g2572(n5154 ,n1058 ,n4876);
    nor g2573(n5153 ,n1058 ,n4997);
    nor g2574(n5152 ,n1060 ,n4854);
    nor g2575(n5151 ,n1058 ,n4872);
    nor g2576(n5150 ,n1058 ,n4835);
    nor g2577(n5149 ,n1060 ,n4849);
    nor g2578(n5148 ,n1057 ,n4865);
    or g2579(n5147 ,n1693 ,n4894);
    or g2580(n5146 ,n1629 ,n4893);
    or g2581(n5145 ,n1626 ,n4784);
    or g2582(n5144 ,n4591 ,n4929);
    nor g2583(n5143 ,n1030 ,n4854);
    nor g2584(n5142 ,n1061 ,n4825);
    or g2585(n5141 ,n4163 ,n4955);
    nor g2586(n5140 ,n1030 ,n5007);
    nor g2587(n5139 ,n1026 ,n4993);
    nor g2588(n5138 ,n1061 ,n4860);
    nor g2589(n5137 ,n1027 ,n4991);
    or g2590(n5136 ,n1680 ,n4889);
    nor g2591(n5135 ,n1061 ,n4827);
    nor g2592(n5134 ,n1061 ,n4858);
    or g2593(n5133 ,n4195 ,n4942);
    nor g2594(n5132 ,n1026 ,n5005);
    nor g2595(n5131 ,n1061 ,n4823);
    nor g2596(n5130 ,n1030 ,n5009);
    nor g2597(n5129 ,n1030 ,n5003);
    or g2598(n5128 ,n1689 ,n4766);
    nor g2599(n5127 ,n1061 ,n4837);
    or g2600(n5126 ,n4270 ,n4948);
    nor g2601(n5125 ,n1028 ,n5001);
    nor g2602(n5124 ,n1030 ,n4999);
    or g2603(n5123 ,n1682 ,n4775);
    or g2604(n5122 ,n4939 ,n4600);
    nor g2605(n5121 ,n1030 ,n4874);
    nor g2606(n5120 ,n1028 ,n4997);
    nor g2607(n5119 ,n1028 ,n4867);
    or g2608(n5118 ,n1697 ,n4890);
    nor g2609(n5117 ,n1026 ,n4819);
    or g2610(n5116 ,n1685 ,n4779);
    or g2611(n5115 ,n1656 ,n4895);
    nor g2612(n5114 ,n1061 ,n4833);
    or g2613(n5113 ,n4460 ,n4934);
    or g2614(n5112 ,n4119 ,n4925);
    nor g2615(n5208 ,n2369 ,n4831);
    nor g2616(n5207 ,n2369 ,n4856);
    nor g2617(n5206 ,n2369 ,n4844);
    nor g2618(n5205 ,n2369 ,n4841);
    nor g2619(n5204 ,n2369 ,n4837);
    nor g2620(n5203 ,n2369 ,n4833);
    nor g2621(n5202 ,n2369 ,n4827);
    nor g2622(n5201 ,n2369 ,n4825);
    nor g2623(n5200 ,n2369 ,n4821);
    nor g2624(n5199 ,n2369 ,n4870);
    nor g2625(n5198 ,n2369 ,n4860);
    nor g2626(n5197 ,n2369 ,n4858);
    nor g2627(n5196 ,n2369 ,n4852);
    nor g2628(n5195 ,n2369 ,n4823);
    nor g2629(n5194 ,n2369 ,n4829);
    nor g2630(n5193 ,n2369 ,n4839);
    not g2631(n5111 ,n5110);
    not g2632(n5090 ,n5089);
    not g2633(n5085 ,n5084);
    not g2634(n5079 ,n5078);
    nor g2635(n5076 ,n1030 ,n4848);
    or g2636(n5075 ,n1687 ,n4774);
    nor g2637(n5074 ,n1061 ,n4852);
    or g2638(n5073 ,n1710 ,n4788);
    or g2639(n5072 ,n1702 ,n4776);
    nor g2640(n5071 ,n1061 ,n4870);
    or g2641(n5070 ,n1639 ,n4777);
    nor g2642(n5069 ,n1061 ,n4821);
    or g2643(n5068 ,n1653 ,n4778);
    or g2644(n5067 ,n1704 ,n4780);
    or g2645(n5066 ,n1669 ,n4761);
    nor g2646(n5065 ,n1028 ,n4865);
    nor g2647(n5064 ,n1061 ,n4829);
    nor g2648(n5063 ,n1061 ,n1007);
    nor g2649(n5062 ,n1061 ,n1005);
    nor g2650(n5061 ,n1061 ,n1008);
    nor g2651(n5060 ,n1061 ,n1006);
    nor g2652(n5059 ,n7313 ,n4885);
    nor g2653(n5058 ,n7313 ,n4884);
    nor g2654(n5057 ,n7313 ,n4883);
    nor g2655(n5056 ,n7313 ,n4879);
    nor g2656(n5055 ,n1046 ,n4983);
    nor g2657(n5054 ,n1046 ,n4980);
    nor g2658(n5053 ,n1046 ,n4964);
    nor g2659(n5052 ,n1046 ,n4986);
    nor g2660(n5051 ,n1045 ,n4794);
    nor g2661(n5050 ,n1045 ,n4804);
    nor g2662(n5049 ,n1045 ,n4979);
    nor g2663(n5048 ,n2366 ,n4963);
    nor g2664(n5047 ,n1046 ,n4810);
    nor g2665(n5046 ,n2365 ,n4806);
    nor g2666(n5045 ,n1045 ,n4791);
    nor g2667(n5044 ,n1058 ,n4990);
    nor g2668(n5043 ,n1058 ,n5008);
    nor g2669(n5042 ,n1058 ,n4861);
    nor g2670(n5041 ,n1060 ,n4873);
    nor g2671(n5040 ,n1057 ,n4818);
    nor g2672(n5039 ,n1058 ,n4850);
    nor g2673(n5038 ,n1057 ,n4868);
    nor g2674(n5037 ,n2365 ,n4984);
    nor g2675(n5036 ,n2366 ,n4981);
    nor g2676(n5035 ,n1046 ,n4965);
    nor g2677(n5034 ,n1046 ,n4985);
    nor g2678(n5033 ,n1045 ,n4793);
    nor g2679(n5032 ,n1045 ,n4978);
    nor g2680(n5031 ,n2365 ,n4962);
    nor g2681(n5030 ,n2365 ,n4805);
    nor g2682(n5029 ,n1045 ,n4811);
    nor g2683(n5028 ,n2366 ,n4807);
    nor g2684(n5027 ,n1046 ,n4792);
    nor g2685(n5026 ,n1030 ,n4994);
    nor g2686(n5025 ,n1061 ,n4842);
    nor g2687(n5024 ,n1028 ,n4871);
    nor g2688(n5023 ,n1026 ,n4850);
    nor g2689(n5022 ,n1061 ,n4847);
    nor g2690(n5021 ,n1061 ,n4845);
    or g2691(n5020 ,n4280 ,n4940);
    nor g2692(n5019 ,n1028 ,n4834);
    nor g2693(n5018 ,n1030 ,n4868);
    nor g2694(n5017 ,n1030 ,n4861);
    nor g2695(n5016 ,n1028 ,n4862);
    nor g2696(n5015 ,n1061 ,n4846);
    or g2697(n5014 ,n1699 ,n4773);
    nor g2698(n5110 ,n2365 ,n4974);
    xnor g2699(n5013 ,n3942 ,n4613);
    xnor g2700(n5012 ,n4615 ,n4619);
    xnor g2701(n5011 ,n3944 ,n4621);
    nor g2702(n5109 ,n7398 ,n4885);
    nor g2703(n5108 ,n2369 ,n4847);
    nor g2704(n5107 ,n2369 ,n4846);
    nor g2705(n5106 ,n2369 ,n4845);
    or g2706(n5105 ,n1045 ,n4789);
    nor g2707(n5104 ,n2369 ,n4842);
    xnor g2708(n5010 ,n4609 ,n4611);
    nor g2709(n5103 ,n2369 ,n1005);
    nor g2710(n5102 ,n2369 ,n1006);
    nor g2711(n5101 ,n2369 ,n1007);
    nor g2712(n5100 ,n7398 ,n4886);
    or g2713(n5099 ,n1373 ,n4888);
    nor g2714(n5098 ,n7398 ,n4883);
    nor g2715(n5097 ,n7398 ,n4882);
    nor g2716(n5096 ,n7398 ,n4879);
    nor g2717(n5095 ,n7398 ,n4880);
    or g2718(n5094 ,n2365 ,n4958);
    or g2719(n5093 ,n2365 ,n4959);
    nor g2720(n5092 ,n7398 ,n4884);
    nor g2721(n5091 ,n7398 ,n4881);
    nor g2722(n5089 ,n1046 ,n4973);
    or g2723(n5088 ,n1046 ,n4790);
    nor g2724(n5087 ,n2369 ,n1008);
    nor g2725(n5086 ,n1029 ,n4785);
    nor g2726(n5084 ,n4918 ,n4390);
    nor g2727(n5083 ,n1029 ,n4787);
    nor g2728(n5082 ,n1029 ,n4786);
    nor g2729(n5081 ,n4597 ,n4944);
    nor g2730(n5080 ,n1029 ,n4781);
    nor g2731(n5078 ,n4943 ,n4246);
    nor g2732(n5077 ,n4675 ,n4908);
    not g2733(n5009 ,n5008);
    not g2734(n5007 ,n5006);
    not g2735(n5005 ,n5004);
    not g2736(n5003 ,n5002);
    not g2737(n5001 ,n5000);
    not g2738(n4999 ,n4998);
    not g2739(n4997 ,n4996);
    not g2740(n4995 ,n4994);
    not g2741(n4993 ,n4992);
    not g2742(n4991 ,n4990);
    not g2743(n4986 ,n4985);
    not g2744(n4983 ,n4984);
    not g2745(n4980 ,n4981);
    not g2746(n4979 ,n4978);
    not g2747(n4974 ,n4973);
    not g2748(n4964 ,n4965);
    not g2749(n4963 ,n4962);
    not g2750(n4959 ,n4958);
    or g2751(n4955 ,n7366 ,n4651);
    or g2752(n4954 ,n7354 ,n4650);
    or g2753(n4953 ,n3606 ,n4649);
    or g2754(n4952 ,n3546 ,n4578);
    or g2755(n4951 ,n3566 ,n4644);
    or g2756(n4950 ,n3545 ,n4643);
    or g2757(n4949 ,n3533 ,n4641);
    or g2758(n4948 ,n2556 ,n4562);
    or g2759(n4947 ,n4029 ,n4587);
    or g2760(n4946 ,n3273 ,n4579);
    or g2761(n4945 ,n4505 ,n4563);
    nor g2762(n4944 ,n1021 ,n4633);
    nor g2763(n4943 ,n1021 ,n4639);
    nor g2764(n4942 ,n1057 ,n4614);
    nor g2765(n4941 ,n1060 ,n4610);
    nor g2766(n4940 ,n1057 ,n4620);
    nor g2767(n4939 ,n1060 ,n4618);
    nor g2768(n4938 ,n1057 ,n4616);
    nor g2769(n4937 ,n1057 ,n4622);
    nor g2770(n4936 ,n1057 ,n4612);
    nor g2771(n4935 ,n1057 ,n4624);
    nor g2772(n4934 ,n1057 ,n4632);
    nor g2773(n4933 ,n1057 ,n4627);
    or g2774(n4932 ,n4417 ,n4568);
    or g2775(n4931 ,n4406 ,n4567);
    or g2776(n4930 ,n4407 ,n4566);
    or g2777(n4929 ,n4279 ,n4565);
    or g2778(n4928 ,n4213 ,n4672);
    or g2779(n4927 ,n4204 ,n4555);
    or g2780(n4926 ,n4203 ,n4670);
    or g2781(n4925 ,n4459 ,n4629);
    nor g2782(n4924 ,n1027 ,n4614);
    or g2783(n4923 ,n4194 ,n4629);
    nor g2784(n4922 ,n1028 ,n4610);
    nor g2785(n4921 ,n1028 ,n4616);
    nor g2786(n4920 ,n1030 ,n4624);
    or g2787(n4919 ,n4189 ,n4667);
    nor g2788(n4918 ,n1022 ,n4639);
    or g2789(n4917 ,n3941 ,n4726);
    or g2790(n4916 ,n4554 ,n4601);
    or g2791(n4915 ,n3807 ,n4722);
    nor g2792(n4914 ,n1026 ,n4620);
    or g2793(n4913 ,n4142 ,n4598);
    or g2794(n4912 ,n3794 ,n4720);
    or g2795(n4911 ,n4718 ,n4630);
    nor g2796(n4910 ,n1026 ,n4622);
    nor g2797(n4909 ,n1027 ,n4612);
    nor g2798(n4908 ,n1022 ,n4633);
    or g2799(n4907 ,n3789 ,n4716);
    or g2800(n4906 ,n4454 ,n4581);
    or g2801(n4905 ,n3301 ,n4630);
    or g2802(n4904 ,n4661 ,n4467);
    or g2803(n4903 ,n3850 ,n4710);
    or g2804(n4902 ,n3824 ,n4709);
    nor g2805(n4901 ,n1026 ,n4627);
    or g2806(n4900 ,n4295 ,n4570);
    or g2807(n4899 ,n4234 ,n4571);
    or g2808(n4898 ,n4233 ,n4572);
    or g2809(n4897 ,n4268 ,n4560);
    or g2810(n4896 ,n4175 ,n4665);
    or g2811(n4895 ,n3986 ,n4553);
    or g2812(n4894 ,n3992 ,n4543);
    or g2813(n4893 ,n3993 ,n4547);
    or g2814(n4892 ,n7324 ,n4652);
    or g2815(n4891 ,n3962 ,n4635);
    or g2816(n4890 ,n3950 ,n4534);
    or g2817(n4889 ,n3997 ,n4551);
    nor g2818(n4888 ,n2972 ,n4558);
    nor g2819(n4887 ,n1028 ,n4617);
    nor g2820(n5008 ,n4695 ,n4653);
    nor g2821(n5006 ,n4294 ,n4557);
    nor g2822(n5004 ,n4677 ,n4657);
    nor g2823(n5002 ,n4690 ,n4700);
    nor g2824(n5000 ,n4691 ,n4699);
    nor g2825(n4998 ,n4689 ,n4701);
    nor g2826(n4996 ,n4692 ,n4698);
    nor g2827(n4994 ,n4697 ,n4655);
    nor g2828(n4992 ,n4694 ,n4658);
    nor g2829(n4990 ,n4654 ,n4696);
    nor g2830(n4989 ,n2601 ,n4608);
    nor g2831(n4988 ,n1459 ,n4748);
    nor g2832(n4987 ,n1465 ,n4742);
    nor g2833(n4985 ,n2616 ,n4744);
    nor g2834(n4984 ,n2614 ,n4745);
    nor g2835(n4982 ,n2612 ,n4743);
    nor g2836(n4981 ,n2610 ,n4628);
    nor g2837(n4978 ,n2609 ,n4750);
    nor g2838(n4977 ,n2632 ,n4743);
    nor g2839(n4976 ,n2607 ,n4748);
    nor g2840(n4975 ,n1456 ,n4747);
    nor g2841(n4973 ,n2605 ,n4749);
    nor g2842(n4972 ,n2602 ,n4742);
    nor g2843(n4971 ,n2631 ,n4747);
    nor g2844(n4970 ,n2600 ,n4746);
    nor g2845(n4969 ,n2597 ,n4628);
    nor g2846(n4968 ,n2621 ,n4625);
    nor g2847(n4967 ,n2627 ,n4742);
    nor g2848(n4966 ,n2628 ,n4749);
    nor g2849(n4965 ,n2594 ,n4625);
    nor g2850(n4962 ,n2593 ,n4744);
    nor g2851(n4961 ,n2569 ,n4748);
    nor g2852(n4960 ,n2629 ,n4750);
    nor g2853(n4958 ,n2630 ,n4748);
    nor g2854(n4957 ,n1458 ,n4749);
    nor g2855(n4956 ,n2596 ,n4747);
    not g2856(n4878 ,n4877);
    not g2857(n4876 ,n4875);
    not g2858(n4874 ,n4873);
    not g2859(n4872 ,n4871);
    not g2860(n4870 ,n4869);
    not g2861(n4867 ,n4866);
    not g2862(n4865 ,n4864);
    not g2863(n4863 ,n4862);
    not g2864(n4860 ,n4859);
    not g2865(n4858 ,n4857);
    not g2866(n4856 ,n4855);
    not g2867(n4854 ,n4853);
    not g2868(n4852 ,n4851);
    not g2869(n4849 ,n4848);
    not g2870(n4844 ,n4843);
    not g2871(n4841 ,n4840);
    not g2872(n4839 ,n4838);
    not g2873(n4837 ,n4836);
    not g2874(n4835 ,n4834);
    not g2875(n4833 ,n4832);
    not g2876(n4831 ,n4830);
    not g2877(n4829 ,n4828);
    not g2878(n4827 ,n4826);
    not g2879(n4825 ,n4824);
    not g2880(n4823 ,n4822);
    not g2881(n4821 ,n4820);
    not g2882(n4819 ,n4818);
    not g2883(n4810 ,n4811);
    not g2884(n4806 ,n4807);
    not g2885(n4804 ,n4805);
    not g2886(n4798 ,n4799);
    not g2887(n4794 ,n4793);
    not g2888(n4791 ,n4792);
    not g2889(n4790 ,n4789);
    or g2890(n4788 ,n3969 ,n4530);
    xnor g2891(n4787 ,n4222 ,n2393);
    xnor g2892(n4786 ,n4223 ,n2398);
    xnor g2893(n4785 ,n4224 ,n2414);
    or g2894(n4784 ,n3996 ,n4542);
    or g2895(n4783 ,n3989 ,n4637);
    or g2896(n4782 ,n3988 ,n4636);
    xnor g2897(n4781 ,n4221 ,n2381);
    or g2898(n4780 ,n3983 ,n4546);
    or g2899(n4779 ,n3981 ,n4526);
    or g2900(n4778 ,n3978 ,n4527);
    or g2901(n4777 ,n3976 ,n4528);
    or g2902(n4776 ,n4001 ,n4529);
    or g2903(n4775 ,n3970 ,n4544);
    or g2904(n4774 ,n3966 ,n4531);
    or g2905(n4773 ,n3963 ,n4552);
    or g2906(n4772 ,n3980 ,n4532);
    or g2907(n4771 ,n3982 ,n4533);
    or g2908(n4770 ,n3948 ,n4540);
    or g2909(n4769 ,n3990 ,n4535);
    or g2910(n4768 ,n3991 ,n4539);
    or g2911(n4767 ,n3975 ,n4536);
    or g2912(n4766 ,n3961 ,n4537);
    or g2913(n4765 ,n3949 ,n4538);
    or g2914(n4764 ,n4000 ,n4640);
    or g2915(n4763 ,n3987 ,n4634);
    or g2916(n4762 ,n3995 ,n4638);
    or g2917(n4761 ,n3985 ,n4541);
    or g2918(n4760 ,n4114 ,n4663);
    or g2919(n4759 ,n3974 ,n4629);
    xnor g2920(n4886 ,n4313 ,n3372);
    xnor g2921(n4758 ,n4335 ,n4323);
    xnor g2922(n4757 ,n4354 ,n4343);
    xnor g2923(n4756 ,n4345 ,n3766);
    xnor g2924(n4755 ,n4341 ,n4319);
    xnor g2925(n4754 ,n4339 ,n4337);
    xnor g2926(n4885 ,n4308 ,n3357);
    xnor g2927(n4884 ,n4307 ,n3385);
    xnor g2928(n4883 ,n4318 ,n3373);
    xnor g2929(n4753 ,n4321 ,n3765);
    xnor g2930(n4882 ,n4315 ,n3378);
    xnor g2931(n4881 ,n4311 ,n3383);
    xnor g2932(n4880 ,n4317 ,n3409);
    xnor g2933(n4879 ,n4309 ,n3380);
    xnor g2934(n4752 ,n4350 ,n3764);
    xnor g2935(n4751 ,n4514 ,n4330);
    nor g2936(n4877 ,n4599 ,n4684);
    nor g2937(n4875 ,n4683 ,n4589);
    nor g2938(n4873 ,n4680 ,n4592);
    nor g2939(n4871 ,n4602 ,n4685);
    xnor g2940(n4869 ,n3395 ,n4325);
    nor g2941(n4868 ,n4676 ,n4586);
    nor g2942(n4866 ,n4688 ,n4706);
    nor g2943(n4864 ,n4674 ,n4574);
    nor g2944(n4862 ,n4681 ,n4593);
    nor g2945(n4861 ,n4682 ,n4595);
    xnor g2946(n4859 ,n3394 ,n4329);
    xnor g2947(n4857 ,n3392 ,n4328);
    xnor g2948(n4855 ,n3388 ,n4352);
    nor g2949(n4853 ,n4384 ,n4569);
    xnor g2950(n4851 ,n3404 ,n4349);
    nor g2951(n4850 ,n4678 ,n4588);
    nor g2952(n4848 ,n4603 ,n4741);
    xnor g2953(n4847 ,n4312 ,n3391);
    xnor g2954(n4846 ,n4314 ,n3354);
    xnor g2955(n4845 ,n4316 ,n3396);
    xnor g2956(n4843 ,n3397 ,n4326);
    xnor g2957(n4842 ,n4310 ,n3393);
    xnor g2958(n4840 ,n3390 ,n4333);
    xnor g2959(n4838 ,n3387 ,n4349);
    xnor g2960(n4836 ,n3400 ,n4353);
    nor g2961(n4834 ,n4687 ,n4604);
    xnor g2962(n4832 ,n3399 ,n4325);
    xnor g2963(n4830 ,n3381 ,n4333);
    xnor g2964(n4828 ,n3407 ,n4326);
    xnor g2965(n4826 ,n3402 ,n4329);
    xnor g2966(n4824 ,n3403 ,n4328);
    xnor g2967(n4822 ,n3405 ,n4352);
    xnor g2968(n4820 ,n3389 ,n4353);
    nor g2969(n4818 ,n4679 ,n4590);
    nor g2970(n4817 ,n2553 ,n4744);
    nor g2971(n4816 ,n2576 ,n4743);
    nor g2972(n4815 ,n2570 ,n4628);
    nor g2973(n4814 ,n2552 ,n4745);
    nor g2974(n4813 ,n2568 ,n4750);
    nor g2975(n4812 ,n1486 ,n4625);
    nor g2976(n4811 ,n2558 ,n4608);
    nor g2977(n4809 ,n2557 ,n4746);
    nor g2978(n4808 ,n2615 ,n4746);
    nor g2979(n4807 ,n2547 ,n4625);
    nor g2980(n4805 ,n2548 ,n4745);
    nor g2981(n4803 ,n1565 ,n4744);
    nor g2982(n4802 ,n2549 ,n4608);
    nor g2983(n4801 ,n1566 ,n4746);
    nor g2984(n4800 ,n2586 ,n4742);
    nor g2985(n4799 ,n1455 ,n4608);
    nor g2986(n4797 ,n1451 ,n4628);
    nor g2987(n4796 ,n2584 ,n4749);
    nor g2988(n4795 ,n1585 ,n4750);
    nor g2989(n4793 ,n1569 ,n4743);
    nor g2990(n4792 ,n1433 ,n4745);
    nor g2991(n4789 ,n2626 ,n4747);
    nor g2992(n4741 ,n1025 ,n4359);
    or g2993(n4740 ,n3551 ,n4435);
    or g2994(n4739 ,n3871 ,n4434);
    or g2995(n4738 ,n3577 ,n4404);
    or g2996(n4737 ,n3864 ,n4433);
    or g2997(n4736 ,n4432 ,n3862);
    or g2998(n4735 ,n3861 ,n4431);
    or g2999(n4734 ,n4145 ,n4242);
    or g3000(n4733 ,n3585 ,n4429);
    or g3001(n4732 ,n4426 ,n4287);
    or g3002(n4731 ,n4425 ,n4285);
    or g3003(n4730 ,n4424 ,n4283);
    or g3004(n4729 ,n2591 ,n4281);
    or g3005(n4728 ,n3505 ,n4420);
    or g3006(n4727 ,n4043 ,n4277);
    or g3007(n4726 ,n4040 ,n4267);
    or g3008(n4725 ,n4416 ,n3808);
    or g3009(n4724 ,n2573 ,n4415);
    or g3010(n4723 ,n4414 ,n3793);
    or g3011(n4722 ,n2572 ,n4413);
    or g3012(n4721 ,n2554 ,n4408);
    or g3013(n4720 ,n2559 ,n4258);
    or g3014(n4719 ,n3328 ,n4504);
    or g3015(n4718 ,n4046 ,n4257);
    or g3016(n4717 ,n3318 ,n4403);
    or g3017(n4716 ,n3797 ,n4402);
    or g3018(n4715 ,n3300 ,n4401);
    or g3019(n4714 ,n3882 ,n4396);
    or g3020(n4713 ,n3281 ,n4398);
    or g3021(n4712 ,n4021 ,n4241);
    or g3022(n4711 ,n3780 ,n4397);
    or g3023(n4710 ,n3853 ,n4395);
    or g3024(n4709 ,n4394 ,n3887);
    or g3025(n4708 ,n4144 ,n4237);
    or g3026(n4707 ,n3256 ,n4449);
    nor g3027(n4706 ,n1022 ,n4365);
    nor g3028(n4705 ,n1026 ,n4346);
    or g3029(n4704 ,n4123 ,n4422);
    nor g3030(n4703 ,n1026 ,n4331);
    or g3031(n4702 ,n3721 ,n4275);
    nor g3032(n4701 ,n1022 ,n4363);
    nor g3033(n4700 ,n1024 ,n4361);
    nor g3034(n4699 ,n1024 ,n4359);
    nor g3035(n4698 ,n1022 ,n4358);
    nor g3036(n4697 ,n1025 ,n4517);
    nor g3037(n4696 ,n1021 ,n4376);
    nor g3038(n4695 ,n1025 ,n4374);
    nor g3039(n4694 ,n1021 ,n4366);
    nor g3040(n4693 ,n1021 ,n4356);
    nor g3041(n4692 ,n1021 ,n4357);
    nor g3042(n4691 ,n1025 ,n4358);
    nor g3043(n4690 ,n1021 ,n4360);
    nor g3044(n4689 ,n1021 ,n4362);
    nor g3045(n4688 ,n1021 ,n4364);
    nor g3046(n4687 ,n1021 ,n4363);
    or g3047(n4686 ,n3561 ,n4437);
    nor g3048(n4685 ,n1021 ,n4367);
    nor g3049(n4684 ,n1025 ,n4519);
    nor g3050(n4683 ,n1021 ,n4377);
    nor g3051(n4682 ,n1021 ,n4368);
    nor g3052(n4681 ,n1021 ,n4518);
    nor g3053(n4680 ,n1021 ,n4370);
    nor g3054(n4679 ,n1021 ,n4372);
    nor g3055(n4678 ,n1021 ,n4375);
    nor g3056(n4677 ,n1021 ,n4365);
    nor g3057(n4676 ,n1025 ,n4371);
    nor g3058(n4675 ,n1021 ,n4369);
    nor g3059(n4674 ,n1025 ,n4361);
    nor g3060(n4673 ,n1060 ,n4515);
    nor g3061(n4672 ,n1058 ,n4322);
    nor g3062(n4671 ,n1057 ,n4348);
    nor g3063(n4670 ,n1058 ,n4513);
    nor g3064(n4669 ,n1058 ,n4324);
    nor g3065(n4668 ,n1060 ,n4355);
    nor g3066(n4667 ,n1057 ,n4331);
    nor g3067(n4666 ,n1058 ,n4346);
    nor g3068(n4665 ,n1060 ,n4336);
    nor g3069(n4664 ,n1057 ,n4344);
    nor g3070(n4663 ,n1060 ,n4342);
    nor g3071(n4662 ,n1057 ,n4351);
    nor g3072(n4661 ,n1058 ,n4320);
    nor g3073(n4660 ,n1057 ,n4340);
    nor g3074(n4659 ,n1057 ,n4338);
    nor g3075(n4658 ,n1022 ,n4367);
    nor g3076(n4657 ,n1022 ,n4364);
    nor g3077(n4656 ,n3908 ,n4379);
    nor g3078(n4655 ,n1022 ,n4518);
    nor g3079(n4654 ,n1022 ,n4375);
    nor g3080(n4653 ,n1022 ,n4372);
    or g3081(n4652 ,n3681 ,n4448);
    or g3082(n4651 ,n2886 ,n4445);
    or g3083(n4650 ,n3678 ,n4443);
    or g3084(n4649 ,n2753 ,n4489);
    nor g3085(n4648 ,n1026 ,n4515);
    nor g3086(n4647 ,n1028 ,n4322);
    nor g3087(n4646 ,n1026 ,n4355);
    nor g3088(n4645 ,n1026 ,n4348);
    or g3089(n4644 ,n4207 ,n4452);
    or g3090(n4643 ,n2722 ,n4507);
    nor g3091(n4642 ,n1030 ,n4324);
    or g3092(n4641 ,n3060 ,n4506);
    nor g3093(n4750 ,n1029 ,n4225);
    nor g3094(n4749 ,n1029 ,n4255);
    nor g3095(n4748 ,n1029 ,n4253);
    nor g3096(n4747 ,n1029 ,n4252);
    nor g3097(n4746 ,n1029 ,n4251);
    nor g3098(n4745 ,n1029 ,n4249);
    nor g3099(n4744 ,n1029 ,n4230);
    nor g3100(n4743 ,n1029 ,n4226);
    nor g3101(n4742 ,n1029 ,n4256);
    not g3102(n4632 ,n4631);
    not g3103(n4627 ,n4626);
    not g3104(n4624 ,n4623);
    not g3105(n4622 ,n4621);
    not g3106(n4620 ,n4619);
    not g3107(n4618 ,n4617);
    not g3108(n4616 ,n4615);
    not g3109(n4614 ,n4613);
    not g3110(n4612 ,n4611);
    not g3111(n4610 ,n4609);
    or g3112(n4607 ,n3719 ,n4421);
    nor g3113(n4606 ,n1022 ,n4356);
    or g3114(n4605 ,n4157 ,n4419);
    nor g3115(n4604 ,n1022 ,n4362);
    nor g3116(n4603 ,n1022 ,n4357);
    nor g3117(n4602 ,n1022 ,n4366);
    or g3118(n4601 ,n3716 ,n4266);
    or g3119(n4600 ,n3715 ,n4265);
    nor g3120(n4599 ,n1022 ,n4377);
    or g3121(n4598 ,n3713 ,n4412);
    nor g3122(n4597 ,n1022 ,n4368);
    or g3123(n4596 ,n3712 ,n4261);
    nor g3124(n4595 ,n1022 ,n4369);
    nor g3125(n4594 ,n3907 ,n4380);
    nor g3126(n4593 ,n1022 ,n4517);
    nor g3127(n4592 ,n1024 ,n4371);
    nor g3128(n4591 ,n3909 ,n4381);
    nor g3129(n4590 ,n1024 ,n4374);
    nor g3130(n4589 ,n1022 ,n4519);
    nor g3131(n4588 ,n1022 ,n4376);
    or g3132(n4587 ,n3705 ,n4250);
    nor g3133(n4586 ,n1022 ,n4370);
    or g3134(n4585 ,n4107 ,n4494);
    nor g3135(n4584 ,n1028 ,n4351);
    nor g3136(n4583 ,n1027 ,n4344);
    or g3137(n4582 ,n4028 ,n4469);
    or g3138(n4581 ,n2757 ,n4400);
    or g3139(n4580 ,n3692 ,n4465);
    or g3140(n4579 ,n2659 ,n4503);
    or g3141(n4578 ,n2730 ,n4502);
    or g3142(n4577 ,n4129 ,n4462);
    nor g3143(n4576 ,n3898 ,n4378);
    nor g3144(n4575 ,n1026 ,n4336);
    nor g3145(n4574 ,n1022 ,n4360);
    or g3146(n4573 ,n4152 ,n4418);
    nor g3147(n4572 ,n1061 ,n4318);
    nor g3148(n4571 ,n1061 ,n4309);
    nor g3149(n4570 ,n1061 ,n4307);
    nor g3150(n4569 ,n1024 ,n4373);
    nor g3151(n4568 ,n1061 ,n4313);
    nor g3152(n4567 ,n1061 ,n4315);
    nor g3153(n4566 ,n1061 ,n4317);
    nor g3154(n4565 ,n1061 ,n4311);
    nor g3155(n4564 ,n1028 ,n4337);
    or g3156(n4563 ,n3056 ,n4455);
    or g3157(n4562 ,n2702 ,n4451);
    or g3158(n4561 ,n4143 ,n4501);
    nor g3159(n4560 ,n1061 ,n4308);
    nor g3160(n4559 ,n1028 ,n4339);
    nor g3161(n4558 ,n2440 ,n4516);
    nor g3162(n4557 ,n1025 ,n4373);
    nor g3163(n4556 ,n1060 ,n4327);
    nor g3164(n4555 ,n1058 ,n4334);
    nor g3165(n4554 ,n1057 ,n4332);
    nor g3166(n4553 ,n1044 ,n4298);
    nor g3167(n4552 ,n1042 ,n4269);
    nor g3168(n4551 ,n1041 ,n4292);
    nor g3169(n4550 ,n1041 ,n4276);
    nor g3170(n4549 ,n1041 ,n4278);
    nor g3171(n4548 ,n1042 ,n4297);
    nor g3172(n4547 ,n1039 ,n4289);
    nor g3173(n4546 ,n1044 ,n4306);
    nor g3174(n4545 ,n1042 ,n4299);
    nor g3175(n4544 ,n1039 ,n4286);
    nor g3176(n4543 ,n1044 ,n4290);
    nor g3177(n4542 ,n1042 ,n4274);
    nor g3178(n4541 ,n1041 ,n4273);
    nor g3179(n4540 ,n1044 ,n4260);
    nor g3180(n4539 ,n1039 ,n4301);
    nor g3181(n4538 ,n1044 ,n4284);
    nor g3182(n4537 ,n1042 ,n4300);
    nor g3183(n4536 ,n1040 ,n4291);
    nor g3184(n4535 ,n1041 ,n4262);
    nor g3185(n4534 ,n1040 ,n4264);
    nor g3186(n4533 ,n1044 ,n4302);
    nor g3187(n4532 ,n1039 ,n4259);
    nor g3188(n4531 ,n1039 ,n4282);
    nor g3189(n4530 ,n1044 ,n4271);
    nor g3190(n4529 ,n1039 ,n4303);
    nor g3191(n4528 ,n1041 ,n4304);
    nor g3192(n4527 ,n1040 ,n4305);
    nor g3193(n4526 ,n1044 ,n4293);
    nor g3194(n4525 ,n1030 ,n4512);
    nor g3195(n4524 ,n1028 ,n4319);
    nor g3196(n4523 ,n1030 ,n4327);
    nor g3197(n4522 ,n1028 ,n4332);
    nor g3198(n4521 ,n1030 ,n4341);
    nor g3199(n4520 ,n1026 ,n4334);
    nor g3200(n4640 ,n2369 ,n4313);
    or g3201(n4639 ,n3734 ,n4516);
    nor g3202(n4638 ,n2369 ,n4309);
    nor g3203(n4637 ,n2369 ,n4307);
    nor g3204(n4636 ,n2369 ,n4318);
    nor g3205(n4635 ,n2369 ,n4308);
    nor g3206(n4634 ,n2369 ,n4311);
    or g3207(n4633 ,n1371 ,n4481);
    nor g3208(n4631 ,n4385 ,n4296);
    nor g3209(n4630 ,n2369 ,n4317);
    nor g3210(n4629 ,n2369 ,n4315);
    nor g3211(n4628 ,n1029 ,n4231);
    nor g3212(n4626 ,n4383 ,n4235);
    nor g3213(n4625 ,n1029 ,n4227);
    nor g3214(n4623 ,n4389 ,n4238);
    nor g3215(n4621 ,n4388 ,n4254);
    nor g3216(n4619 ,n4392 ,n4263);
    nor g3217(n4617 ,n1442 ,n4476);
    nor g3218(n4615 ,n4387 ,n4248);
    nor g3219(n4613 ,n4391 ,n4232);
    nor g3220(n4611 ,n4382 ,n4228);
    nor g3221(n4609 ,n4386 ,n4229);
    nor g3222(n4608 ,n1029 ,n4245);
    not g3223(n4515 ,n4514);
    not g3224(n4513 ,n4512);
    or g3225(n4511 ,n3603 ,n3964);
    or g3226(n4510 ,n7340 ,n4054);
    or g3227(n4509 ,n7343 ,n4052);
    or g3228(n4508 ,n7329 ,n4050);
    or g3229(n4507 ,n7357 ,n3867);
    or g3230(n4506 ,n7325 ,n3855);
    or g3231(n4505 ,n7349 ,n3865);
    or g3232(n4504 ,n7339 ,n3791);
    or g3233(n4503 ,n7314 ,n3872);
    or g3234(n4502 ,n7315 ,n3891);
    nor g3235(n4501 ,n1150 ,n4016);
    or g3236(n4500 ,n4177 ,n3613);
    or g3237(n4499 ,n3618 ,n4218);
    or g3238(n4498 ,n3626 ,n4219);
    or g3239(n4497 ,n3615 ,n4215);
    or g3240(n4496 ,n3597 ,n4212);
    or g3241(n4495 ,n3583 ,n4209);
    or g3242(n4494 ,n3304 ,n3788);
    or g3243(n4493 ,n4208 ,n3880);
    or g3244(n4492 ,n3556 ,n4202);
    or g3245(n4491 ,n2595 ,n3849);
    or g3246(n4490 ,n3521 ,n4191);
    or g3247(n4489 ,n7345 ,n3897);
    or g3248(n4488 ,n3491 ,n4188);
    or g3249(n4487 ,n3294 ,n4179);
    or g3250(n4486 ,n3590 ,n4186);
    or g3251(n4485 ,n3813 ,n4026);
    or g3252(n4484 ,n2581 ,n4035);
    or g3253(n4483 ,n2579 ,n4034);
    or g3254(n4482 ,n3292 ,n3816);
    nor g3255(n4481 ,n3092 ,n3841);
    or g3256(n4480 ,n2564 ,n4032);
    or g3257(n4479 ,n4216 ,n3799);
    or g3258(n4478 ,n3303 ,n3860);
    or g3259(n4477 ,n2561 ,n4031);
    nor g3260(n4476 ,n3093 ,n3792);
    or g3261(n4475 ,n3786 ,n4030);
    or g3262(n4474 ,n3322 ,n4181);
    or g3263(n4473 ,n3873 ,n4045);
    or g3264(n4472 ,n3308 ,n4180);
    or g3265(n4471 ,n3306 ,n3784);
    or g3266(n4470 ,n3290 ,n3827);
    or g3267(n4469 ,n2577 ,n4027);
    or g3268(n4468 ,n3815 ,n4025);
    or g3269(n4467 ,n3331 ,n3822);
    or g3270(n4466 ,n3830 ,n4023);
    or g3271(n4465 ,n3834 ,n3286);
    or g3272(n4464 ,n3839 ,n4022);
    or g3273(n4463 ,n3271 ,n3868);
    or g3274(n4462 ,n3879 ,n4019);
    or g3275(n4461 ,n3803 ,n4018);
    or g3276(n4460 ,n3267 ,n3890);
    or g3277(n4459 ,n3265 ,n3892);
    or g3278(n4458 ,n3264 ,n3893);
    or g3279(n4457 ,n3555 ,n3900);
    or g3280(n4456 ,n4206 ,n3536);
    nor g3281(n4455 ,n1270 ,n4014);
    nor g3282(n4454 ,n1096 ,n4015);
    nor g3283(n4453 ,n1057 ,n3947);
    nor g3284(n4452 ,n1057 ,n3943);
    nor g3285(n4451 ,n1057 ,n3945);
    or g3286(n4450 ,n3627 ,n3999);
    or g3287(n4449 ,n4217 ,n3680);
    or g3288(n4448 ,n3730 ,n3905);
    nor g3289(n4447 ,n1030 ,n3947);
    nor g3290(n4446 ,n1030 ,n3945);
    or g3291(n4445 ,n3729 ,n3903);
    or g3292(n4444 ,n3796 ,n3330);
    or g3293(n4443 ,n3728 ,n3901);
    or g3294(n4442 ,n7337 ,n4056);
    or g3295(n4441 ,n3594 ,n3965);
    or g3296(n4440 ,n3592 ,n3967);
    or g3297(n4439 ,n3588 ,n3968);
    nor g3298(n4438 ,n1026 ,n3943);
    or g3299(n4437 ,n4205 ,n3971);
    or g3300(n4436 ,n3553 ,n3973);
    or g3301(n4435 ,n3671 ,n4200);
    or g3302(n4434 ,n2724 ,n4201);
    or g3303(n4433 ,n2721 ,n4198);
    or g3304(n4432 ,n2803 ,n4197);
    or g3305(n4431 ,n2719 ,n4196);
    or g3306(n4430 ,n3539 ,n3977);
    or g3307(n4429 ,n3703 ,n3781);
    or g3308(n4428 ,n3528 ,n3979);
    or g3309(n4427 ,n3565 ,n3949);
    or g3310(n4426 ,n1670 ,n3845);
    or g3311(n4425 ,n1620 ,n3840);
    or g3312(n4424 ,n1655 ,n3835);
    or g3313(n4423 ,n3829 ,n4150);
    or g3314(n4422 ,n4153 ,n3496);
    or g3315(n4421 ,n3492 ,n3948);
    or g3316(n4420 ,n4187 ,n3656);
    or g3317(n4419 ,n3544 ,n3950);
    or g3318(n4418 ,n3257 ,n4155);
    or g3319(n4417 ,n1701 ,n4000);
    or g3320(n4416 ,n2689 ,n4184);
    or g3321(n4415 ,n3037 ,n3810);
    or g3322(n4414 ,n3038 ,n4183);
    or g3323(n4413 ,n2777 ,n3805);
    or g3324(n4412 ,n4116 ,n3346);
    or g3325(n4411 ,n3804 ,n4149);
    or g3326(n4410 ,n2674 ,n4182);
    or g3327(n4409 ,n3811 ,n4148);
    or g3328(n4408 ,n2820 ,n3800);
    or g3329(n4407 ,n1706 ,n3994);
    or g3330(n4406 ,n1703 ,n3974);
    or g3331(n4405 ,n3848 ,n4151);
    or g3332(n4404 ,n3708 ,n3785);
    or g3333(n4403 ,n3707 ,n3783);
    or g3334(n4402 ,n2546 ,n3999);
    or g3335(n4401 ,n3701 ,n3806);
    or g3336(n4400 ,n3065 ,n4173);
    or g3337(n4399 ,n4103 ,n4024);
    or g3338(n4398 ,n3691 ,n3843);
    or g3339(n4397 ,n2651 ,n4176);
    or g3340(n4396 ,n2634 ,n4178);
    or g3341(n4395 ,n2544 ,n3971);
    or g3342(n4394 ,n1690 ,n3885);
    or g3343(n4393 ,n3262 ,n3984);
    nor g3344(n4392 ,n1021 ,n3957);
    nor g3345(n4391 ,n1025 ,n3954);
    nor g3346(n4390 ,n1025 ,n3958);
    nor g3347(n4389 ,n1021 ,n3952);
    nor g3348(n4388 ,n1021 ,n3955);
    nor g3349(n4387 ,n1025 ,n3953);
    nor g3350(n4386 ,n1021 ,n3959);
    nor g3351(n4385 ,n1021 ,n3951);
    nor g3352(n4384 ,n1025 ,n3972);
    nor g3353(n4383 ,n1025 ,n3956);
    nor g3354(n4382 ,n1021 ,n3960);
    or g3355(n4381 ,n1042 ,n4171);
    or g3356(n4380 ,n1042 ,n4170);
    or g3357(n4379 ,n1042 ,n4172);
    or g3358(n4378 ,n1042 ,n4169);
    or g3359(n4519 ,n3040 ,n3812);
    or g3360(n4518 ,n3041 ,n3795);
    or g3361(n4517 ,n3039 ,n3820);
    nor g3362(n4516 ,n1368 ,n3826);
    nor g3363(n4514 ,n4102 ,n4060);
    nor g3364(n4512 ,n2633 ,n4013);
    not g3365(n4355 ,n4354);
    not g3366(n4351 ,n4350);
    not g3367(n4348 ,n4347);
    not g3368(n4346 ,n4345);
    not g3369(n4344 ,n4343);
    not g3370(n4342 ,n4341);
    not g3371(n4340 ,n4339);
    not g3372(n4338 ,n4337);
    not g3373(n4336 ,n4335);
    not g3374(n4331 ,n4330);
    not g3375(n4324 ,n4323);
    not g3376(n4322 ,n4321);
    not g3377(n4320 ,n4319);
    not g3378(n4317 ,n4316);
    not g3379(n4315 ,n4314);
    not g3380(n4313 ,n4312);
    not g3381(n4311 ,n4310);
    xnor g3382(n4306 ,n1[74] ,n3217);
    xnor g3383(n4305 ,n1[76] ,n3252);
    xnor g3384(n4304 ,n1[77] ,n3190);
    xnor g3385(n4303 ,n1[78] ,n3250);
    xnor g3386(n4302 ,n1[84] ,n3174);
    xnor g3387(n4301 ,n1[88] ,n3172);
    xnor g3388(n4300 ,n1[90] ,n3236);
    xnor g3389(n4299 ,n1[92] ,n3234);
    xnor g3390(n4298 ,n1[72] ,n3222);
    xnor g3391(n4297 ,n1[65] ,n3166);
    nor g3392(n4296 ,n1024 ,n3960);
    or g3393(n4295 ,n1665 ,n3989);
    nor g3394(n4294 ,n1022 ,n3972);
    xnor g3395(n4293 ,n1[75] ,n3198);
    xnor g3396(n4292 ,n1[68] ,n3229);
    xnor g3397(n4291 ,n1[89] ,n3237);
    xnor g3398(n4290 ,n1[71] ,n3185);
    xnor g3399(n4289 ,n1[70] ,n3195);
    or g3400(n4288 ,n3847 ,n4161);
    or g3401(n4287 ,n2710 ,n4160);
    xnor g3402(n4286 ,n1[79] ,n3194);
    or g3403(n4285 ,n2708 ,n4159);
    xnor g3404(n4284 ,n1[91] ,n3247);
    or g3405(n4283 ,n2759 ,n4158);
    xnor g3406(n4282 ,n1[81] ,n3192);
    or g3407(n4281 ,n2707 ,n3949);
    nor g3408(n4280 ,n4044 ,n4168);
    or g3409(n4279 ,n1621 ,n3987);
    xnor g3410(n4278 ,n1[66] ,n3189);
    or g3411(n4277 ,n3005 ,n3833);
    xnor g3412(n4276 ,n1[67] ,n3196);
    nor g3413(n4275 ,n4042 ,n4167);
    xnor g3414(n4274 ,n1[69] ,n3218);
    xnor g3415(n4273 ,n1[73] ,n3203);
    or g3416(n4272 ,n3821 ,n4156);
    xnor g3417(n4271 ,n1[80] ,n3245);
    nor g3418(n4270 ,n4041 ,n4166);
    xnor g3419(n4269 ,n1[82] ,n3241);
    or g3420(n4268 ,n1658 ,n3962);
    or g3421(n4267 ,n3032 ,n3817);
    nor g3422(n4266 ,n4039 ,n4038);
    nor g3423(n4265 ,n4037 ,n4036);
    xnor g3424(n4264 ,n1[85] ,n3230);
    nor g3425(n4263 ,n1022 ,n3956);
    xnor g3426(n4262 ,n1[87] ,n3173);
    nor g3427(n4261 ,n4033 ,n4165);
    xnor g3428(n4260 ,n1[86] ,n3224);
    xnor g3429(n4259 ,n1[83] ,n3214);
    or g3430(n4258 ,n2678 ,n4154);
    or g3431(n4257 ,n2813 ,n3790);
    xor g3432(n4256 ,n3178 ,n3156);
    xor g3433(n4255 ,n3179 ,n3157);
    nor g3434(n4254 ,n1022 ,n3954);
    xor g3435(n4253 ,n3183 ,n3155);
    xor g3436(n4252 ,n3187 ,n3152);
    xor g3437(n4251 ,n3188 ,n3171);
    or g3438(n4250 ,n4115 ,n3984);
    xor g3439(n4249 ,n3227 ,n3160);
    nor g3440(n4248 ,n1022 ,n3952);
    or g3441(n4247 ,n4113 ,n3964);
    nor g3442(n4246 ,n1022 ,n3958);
    xnor g3443(n4245 ,n3153 ,n3161);
    or g3444(n4244 ,n4112 ,n3965);
    or g3445(n4243 ,n4111 ,n3967);
    or g3446(n4242 ,n4122 ,n3948);
    or g3447(n4241 ,n3696 ,n4104);
    or g3448(n4240 ,n4106 ,n3973);
    or g3449(n4239 ,n4109 ,n3977);
    nor g3450(n4238 ,n1022 ,n3953);
    or g3451(n4237 ,n4121 ,n3950);
    or g3452(n4236 ,n4105 ,n3979);
    nor g3453(n4235 ,n1022 ,n3957);
    or g3454(n4234 ,n1624 ,n3995);
    or g3455(n4233 ,n1686 ,n3988);
    nor g3456(n4232 ,n1022 ,n3955);
    xnor g3457(n4231 ,n3154 ,n3163);
    xor g3458(n4230 ,n3233 ,n3169);
    nor g3459(n4229 ,n1024 ,n3951);
    nor g3460(n4228 ,n1024 ,n3959);
    xnor g3461(n4227 ,n3235 ,n2409);
    xor g3462(n4226 ,n3240 ,n3168);
    xor g3463(n4225 ,n3242 ,n3175);
    or g3464(n4377 ,n2971 ,n4012);
    xnor g3465(n4224 ,n3228 ,n2396);
    xnor g3466(n4223 ,n3220 ,n2404);
    or g3467(n4376 ,n1370 ,n4146);
    or g3468(n4375 ,n2620 ,n4004);
    or g3469(n4374 ,n2550 ,n4005);
    xnor g3470(n4373 ,n2538 ,n3486);
    or g3471(n4372 ,n2571 ,n4006);
    xnor g3472(n4222 ,n3186 ,n2430);
    or g3473(n4371 ,n2545 ,n4007);
    or g3474(n4370 ,n2624 ,n4008);
    or g3475(n4369 ,n2562 ,n4009);
    or g3476(n4368 ,n2551 ,n4011);
    xnor g3477(n4221 ,n3232 ,n2405);
    or g3478(n4367 ,n1419 ,n3818);
    or g3479(n4366 ,n3683 ,n4117);
    or g3480(n4365 ,n1452 ,n3825);
    or g3481(n4364 ,n1461 ,n3828);
    or g3482(n4363 ,n1460 ,n3831);
    or g3483(n4362 ,n1411 ,n3832);
    or g3484(n4361 ,n1431 ,n3837);
    or g3485(n4360 ,n1379 ,n3842);
    or g3486(n4359 ,n1424 ,n3846);
    or g3487(n4358 ,n1406 ,n3854);
    or g3488(n4357 ,n2922 ,n4118);
    or g3489(n4356 ,n1387 ,n3870);
    nor g3490(n4354 ,n4099 ,n4057);
    xnor g3491(n4353 ,n3393 ,n3404);
    xnor g3492(n4352 ,n3408 ,n3395);
    nor g3493(n4350 ,n4101 ,n4059);
    xnor g3494(n4349 ,n3401 ,n3389);
    nor g3495(n4347 ,n2565 ,n4010);
    nor g3496(n4345 ,n4098 ,n4055);
    nor g3497(n4343 ,n4097 ,n4053);
    nor g3498(n4341 ,n4096 ,n4049);
    nor g3499(n4339 ,n4095 ,n4048);
    nor g3500(n4337 ,n4094 ,n4047);
    nor g3501(n4335 ,n4092 ,n4020);
    nor g3502(n4334 ,n1415 ,n3904);
    xnor g3503(n4333 ,n3398 ,n3392);
    nor g3504(n4332 ,n2917 ,n4128);
    nor g3505(n4330 ,n4100 ,n4058);
    xnor g3506(n4329 ,n3354 ,n3407);
    xnor g3507(n4328 ,n3391 ,n3381);
    nor g3508(n4327 ,n1416 ,n3851);
    xnor g3509(n4326 ,n3406 ,n3394);
    xnor g3510(n4325 ,n3396 ,n3405);
    nor g3511(n4323 ,n4091 ,n4051);
    nor g3512(n4321 ,n4003 ,n4017);
    nor g3513(n4319 ,n4093 ,n3878);
    xnor g3514(n4318 ,n3164 ,n3388);
    xnor g3515(n4316 ,n1863 ,n3399);
    xnor g3516(n4314 ,n1825 ,n3402);
    xnor g3517(n4312 ,n1872 ,n3403);
    xnor g3518(n4310 ,n1839 ,n3400);
    xnor g3519(n4309 ,n3162 ,n3397);
    xnor g3520(n4308 ,n3159 ,n3387);
    xnor g3521(n4307 ,n3158 ,n3390);
    nor g3522(n4220 ,n1058 ,n3764);
    or g3523(n4219 ,n7352 ,n3589);
    or g3524(n4218 ,n7327 ,n3625);
    or g3525(n4217 ,n7320 ,n3623);
    or g3526(n4216 ,n7326 ,n3336);
    or g3527(n4215 ,n7358 ,n3612);
    or g3528(n4214 ,n7331 ,n3601);
    or g3529(n4213 ,n7333 ,n3596);
    or g3530(n4212 ,n7377 ,n3595);
    or g3531(n4211 ,n7328 ,n3591);
    or g3532(n4210 ,n7335 ,n3586);
    or g3533(n4209 ,n7365 ,n3579);
    or g3534(n4208 ,n7371 ,n3567);
    or g3535(n4207 ,n7346 ,n3564);
    or g3536(n4206 ,n7321 ,n3569);
    or g3537(n4205 ,n7348 ,n3560);
    or g3538(n4204 ,n7350 ,n3557);
    or g3539(n4203 ,n7351 ,n3554);
    or g3540(n4202 ,n7330 ,n3552);
    or g3541(n4201 ,n7353 ,n3550);
    or g3542(n4200 ,n7376 ,n3549);
    or g3543(n4199 ,n7317 ,n3562);
    or g3544(n4198 ,n7359 ,n3542);
    or g3545(n4197 ,n7318 ,n3541);
    or g3546(n4196 ,n7360 ,n3540);
    or g3547(n4195 ,n7362 ,n3538);
    or g3548(n4194 ,n7364 ,n3534);
    or g3549(n4193 ,n7367 ,n3531);
    or g3550(n4192 ,n7370 ,n3527);
    or g3551(n4191 ,n7332 ,n3518);
    or g3552(n4190 ,n7323 ,n3509);
    or g3553(n4189 ,n7338 ,n3507);
    or g3554(n4188 ,n7347 ,n3489);
    or g3555(n4187 ,n7316 ,n3581);
    or g3556(n4186 ,n7355 ,n3593);
    or g3557(n4185 ,n7334 ,n3604);
    or g3558(n4184 ,n7363 ,n3351);
    or g3559(n4183 ,n7374 ,n3543);
    or g3560(n4182 ,n7368 ,n3335);
    or g3561(n4181 ,n7356 ,n3320);
    or g3562(n4180 ,n7369 ,n3305);
    or g3563(n4179 ,n7372 ,n3291);
    or g3564(n4178 ,n7375 ,n3285);
    or g3565(n4177 ,n7373 ,n3497);
    or g3566(n4176 ,n7361 ,n3619);
    or g3567(n4175 ,n7319 ,n3258);
    or g3568(n4174 ,n7342 ,n3607);
    or g3569(n4173 ,n7336 ,n3757);
    nor g3570(n4172 ,n1156 ,n3435);
    nor g3571(n4171 ,n1158 ,n3425);
    nor g3572(n4170 ,n1307 ,n3471);
    nor g3573(n4169 ,n1155 ,n3477);
    nor g3574(n4168 ,n1136 ,n3620);
    nor g3575(n4167 ,n1135 ,n3313);
    nor g3576(n4166 ,n1297 ,n3578);
    nor g3577(n4165 ,n1133 ,n3341);
    nor g3578(n4164 ,n1131 ,n3621);
    nor g3579(n4163 ,n1126 ,n3616);
    nor g3580(n4162 ,n1299 ,n3609);
    nor g3581(n4161 ,n1293 ,n3523);
    nor g3582(n4160 ,n1290 ,n3520);
    nor g3583(n4159 ,n1300 ,n3516);
    nor g3584(n4158 ,n1140 ,n3513);
    nor g3585(n4157 ,n1138 ,n3353);
    nor g3586(n4156 ,n1294 ,n3502);
    nor g3587(n4155 ,n1295 ,n3573);
    nor g3588(n4154 ,n1146 ,n3329);
    nor g3589(n4153 ,n1289 ,n3353);
    nor g3590(n4152 ,n1291 ,n3353);
    or g3591(n4151 ,n2622 ,n3547);
    or g3592(n4150 ,n2588 ,n3500);
    or g3593(n4149 ,n2580 ,n3344);
    or g3594(n4148 ,n2567 ,n3343);
    or g3595(n4147 ,n2604 ,n3324);
    nor g3596(n4146 ,n3094 ,n3307);
    or g3597(n4145 ,n3682 ,n3287);
    or g3598(n4144 ,n3762 ,n3266);
    nor g3599(n4143 ,n1122 ,n3490);
    nor g3600(n4142 ,n1267 ,n3348);
    nor g3601(n4141 ,n1109 ,n3276);
    nor g3602(n4140 ,n1115 ,n3321);
    nor g3603(n4139 ,n1108 ,n3317);
    nor g3604(n4138 ,n1124 ,n3319);
    nor g3605(n4137 ,n1276 ,n3614);
    nor g3606(n4136 ,n1274 ,n3571);
    nor g3607(n4135 ,n1121 ,n3297);
    nor g3608(n4134 ,n1271 ,n3295);
    nor g3609(n4133 ,n1123 ,n3600);
    nor g3610(n4132 ,n1117 ,n3282);
    nor g3611(n4131 ,n1281 ,n3279);
    nor g3612(n4130 ,n1282 ,n3270);
    nor g3613(n4129 ,n1284 ,n3350);
    nor g3614(n4128 ,n1103 ,n3723);
    nor g3615(n4127 ,n1254 ,n3353);
    nor g3616(n4126 ,n1259 ,n3353);
    nor g3617(n4125 ,n1263 ,n3353);
    nor g3618(n4124 ,n1261 ,n3353);
    nor g3619(n4123 ,n1265 ,n3617);
    nor g3620(n4122 ,n1257 ,n3353);
    nor g3621(n4121 ,n1106 ,n3353);
    nor g3622(n4120 ,n1246 ,n3530);
    nor g3623(n4119 ,n1249 ,n3316);
    nor g3624(n4118 ,n1088 ,n3725);
    nor g3625(n4117 ,n1091 ,n3718);
    nor g3626(n4116 ,n1082 ,n3347);
    nor g3627(n4115 ,n1089 ,n3309);
    nor g3628(n4114 ,n1084 ,n3277);
    nor g3629(n4113 ,n1092 ,n3293);
    nor g3630(n4112 ,n1242 ,n3575);
    nor g3631(n4111 ,n1091 ,n3283);
    nor g3632(n4110 ,n1243 ,n3274);
    nor g3633(n4109 ,n1087 ,n3610);
    nor g3634(n4108 ,n1088 ,n3263);
    nor g3635(n4107 ,n1076 ,n3559);
    nor g3636(n4106 ,n1080 ,n3272);
    nor g3637(n4105 ,n1237 ,n3260);
    nor g3638(n4104 ,n1075 ,n3261);
    nor g3639(n4103 ,n1227 ,n3508);
    nor g3640(n4102 ,n1021 ,n3768);
    nor g3641(n4101 ,n1025 ,n3770);
    nor g3642(n4100 ,n1021 ,n3771);
    nor g3643(n4099 ,n1025 ,n3773);
    nor g3644(n4098 ,n1025 ,n3775);
    nor g3645(n4097 ,n1025 ,n3777);
    nor g3646(n4096 ,n1025 ,n3769);
    nor g3647(n4095 ,n1025 ,n3776);
    nor g3648(n4094 ,n1021 ,n3772);
    nor g3649(n4093 ,n1021 ,n3779);
    nor g3650(n4092 ,n1021 ,n3774);
    nor g3651(n4091 ,n1021 ,n3778);
    nor g3652(n4090 ,n2364 ,n3481);
    nor g3653(n4089 ,n2364 ,n3445);
    nor g3654(n4088 ,n2364 ,n3421);
    nor g3655(n4087 ,n1038 ,n3475);
    nor g3656(n4086 ,n1038 ,n3473);
    nor g3657(n4085 ,n1036 ,n3469);
    nor g3658(n4084 ,n2364 ,n3467);
    nor g3659(n4083 ,n1035 ,n3465);
    nor g3660(n4082 ,n1035 ,n3437);
    nor g3661(n4081 ,n1035 ,n3463);
    nor g3662(n4080 ,n1035 ,n3483);
    nor g3663(n4079 ,n1035 ,n3461);
    nor g3664(n4078 ,n1035 ,n3485);
    nor g3665(n4077 ,n1034 ,n3459);
    nor g3666(n4076 ,n1036 ,n3457);
    nor g3667(n4075 ,n1038 ,n3455);
    nor g3668(n4074 ,n1035 ,n3453);
    nor g3669(n4073 ,n1035 ,n3413);
    nor g3670(n4072 ,n2364 ,n3451);
    nor g3671(n4071 ,n1035 ,n3449);
    nor g3672(n4070 ,n1038 ,n3419);
    nor g3673(n4069 ,n1034 ,n3441);
    nor g3674(n4068 ,n1038 ,n3431);
    nor g3675(n4067 ,n1036 ,n3427);
    nor g3676(n4066 ,n1038 ,n3423);
    nor g3677(n4065 ,n1036 ,n3479);
    nor g3678(n4064 ,n1038 ,n3443);
    nor g3679(n4063 ,n1038 ,n3417);
    nor g3680(n4062 ,n1034 ,n3429);
    nor g3681(n4061 ,n1036 ,n3439);
    nor g3682(n4060 ,n1022 ,n3769);
    nor g3683(n4059 ,n1022 ,n3771);
    nor g3684(n4058 ,n1022 ,n3772);
    nor g3685(n4057 ,n1022 ,n3774);
    or g3686(n4056 ,n2744 ,n3582);
    nor g3687(n4055 ,n1022 ,n3776);
    or g3688(n4054 ,n2741 ,n3576);
    nor g3689(n4053 ,n1022 ,n3778);
    or g3690(n4052 ,n2740 ,n3572);
    nor g3691(n4051 ,n1022 ,n3777);
    or g3692(n4050 ,n2738 ,n3568);
    nor g3693(n4049 ,n1022 ,n3768);
    nor g3694(n4048 ,n1022 ,n3775);
    nor g3695(n4047 ,n1022 ,n3770);
    or g3696(n4046 ,n2555 ,n3710);
    or g3697(n4045 ,n3724 ,n3315);
    nor g3698(n4044 ,n1[59] ,n3510);
    or g3699(n4043 ,n2618 ,n3722);
    nor g3700(n4042 ,n3014 ,n3504);
    nor g3701(n4041 ,n1[51] ,n3340);
    or g3702(n4040 ,n2585 ,n3717);
    nor g3703(n4039 ,n1[49] ,n3598);
    nor g3704(n4038 ,n3033 ,n3754);
    nor g3705(n4037 ,n1[48] ,n3299);
    nor g3706(n4036 ,n2764 ,n3753);
    or g3707(n4035 ,n3655 ,n3275);
    or g3708(n4034 ,n3714 ,n3763);
    nor g3709(n4033 ,n2989 ,n3563);
    or g3710(n4032 ,n3650 ,n3537);
    or g3711(n4031 ,n3647 ,n3608);
    or g3712(n4030 ,n3709 ,n3323);
    or g3713(n4029 ,n3706 ,n3311);
    nor g3714(n4028 ,n3017 ,n3629);
    or g3715(n4027 ,n3658 ,n3302);
    or g3716(n4026 ,n3700 ,n3298);
    or g3717(n4025 ,n3699 ,n3296);
    or g3718(n4024 ,n3694 ,n3289);
    or g3719(n4023 ,n3693 ,n3288);
    or g3720(n4022 ,n3711 ,n3284);
    or g3721(n4021 ,n1649 ,n3278);
    nor g3722(n4020 ,n1022 ,n3773);
    or g3723(n4019 ,n3688 ,n3269);
    or g3724(n4018 ,n3687 ,n3268);
    nor g3725(n4017 ,n1022 ,n3779);
    nor g3726(n4016 ,n3028 ,n3352);
    nor g3727(n4015 ,n2792 ,n3352);
    nor g3728(n4014 ,n2762 ,n3352);
    nor g3729(n4013 ,n1064 ,n3624);
    nor g3730(n4012 ,n1064 ,n3255);
    nor g3731(n4011 ,n1064 ,n3342);
    nor g3732(n4010 ,n1064 ,n3339);
    nor g3733(n4009 ,n1064 ,n3334);
    nor g3734(n4008 ,n1064 ,n3326);
    nor g3735(n4007 ,n1064 ,n3580);
    nor g3736(n4006 ,n1020 ,n3349);
    nor g3737(n4005 ,n1064 ,n3498);
    nor g3738(n4004 ,n1064 ,n3312);
    nor g3739(n4003 ,n1021 ,n3767);
    or g3740(n4002 ,n7322 ,n3599);
    not g3741(n3947 ,n3946);
    not g3742(n3945 ,n3944);
    not g3743(n3943 ,n3942);
    nor g3744(n3941 ,n1058 ,n3766);
    nor g3745(n3940 ,n2364 ,n3480);
    nor g3746(n3939 ,n2364 ,n3468);
    nor g3747(n3938 ,n1035 ,n3474);
    nor g3748(n3937 ,n2364 ,n3472);
    nor g3749(n3936 ,n1035 ,n3466);
    nor g3750(n3935 ,n1035 ,n3464);
    nor g3751(n3934 ,n2364 ,n3462);
    nor g3752(n3933 ,n1036 ,n3482);
    nor g3753(n3932 ,n1036 ,n3460);
    nor g3754(n3931 ,n1035 ,n3438);
    nor g3755(n3930 ,n2364 ,n3484);
    nor g3756(n3929 ,n1034 ,n3458);
    nor g3757(n3928 ,n1038 ,n3456);
    nor g3758(n3927 ,n1038 ,n3454);
    nor g3759(n3926 ,n1034 ,n3452);
    nor g3760(n3925 ,n2364 ,n3412);
    nor g3761(n3924 ,n1035 ,n3450);
    nor g3762(n3923 ,n1035 ,n3448);
    nor g3763(n3922 ,n2364 ,n3444);
    nor g3764(n3921 ,n1035 ,n3418);
    nor g3765(n3920 ,n1038 ,n3442);
    nor g3766(n3919 ,n1034 ,n3440);
    nor g3767(n3918 ,n1036 ,n3436);
    nor g3768(n3917 ,n1036 ,n3428);
    nor g3769(n3916 ,n1036 ,n3426);
    nor g3770(n3915 ,n1038 ,n3422);
    nor g3771(n3914 ,n1034 ,n3420);
    nor g3772(n3913 ,n1036 ,n3430);
    nor g3773(n3912 ,n1034 ,n3416);
    nor g3774(n3911 ,n1038 ,n3478);
    nor g3775(n3910 ,n1060 ,n3765);
    nor g3776(n3909 ,n1[64] ,n3424);
    nor g3777(n3908 ,n1[94] ,n3434);
    nor g3778(n3907 ,n1[95] ,n3470);
    nor g3779(n3906 ,n1033 ,n3382);
    or g3780(n3905 ,n3761 ,n2887);
    nor g3781(n3904 ,n2987 ,n3501);
    or g3782(n3903 ,n3760 ,n3679);
    nor g3783(n3902 ,n1033 ,n3362);
    or g3784(n3901 ,n3759 ,n2884);
    or g3785(n3900 ,n2734 ,n3684);
    nor g3786(n3899 ,n1033 ,n3360);
    nor g3787(n3898 ,n1[93] ,n3476);
    or g3788(n3897 ,n2334 ,n3677);
    nor g3789(n3896 ,n1033 ,n3379);
    nor g3790(n3895 ,n1030 ,n3764);
    nor g3791(n3894 ,n1026 ,n3766);
    or g3792(n3893 ,n2773 ,n3685);
    or g3793(n3892 ,n2774 ,n3726);
    or g3794(n3891 ,n2330 ,n3665);
    or g3795(n3890 ,n2641 ,n3686);
    nor g3796(n3889 ,n1033 ,n3385);
    nor g3797(n3888 ,n1033 ,n3373);
    or g3798(n3887 ,n2643 ,n3737);
    nor g3799(n3886 ,n1033 ,n3363);
    or g3800(n3885 ,n2315 ,n3662);
    nor g3801(n3884 ,n1033 ,n3364);
    nor g3802(n3883 ,n1033 ,n3366);
    or g3803(n3882 ,n2844 ,n3632);
    nor g3804(n3881 ,n1033 ,n3367);
    or g3805(n3880 ,n2737 ,n3675);
    or g3806(n3879 ,n2635 ,n3633);
    nor g3807(n3878 ,n1022 ,n3767);
    nor g3808(n3877 ,n1033 ,n3369);
    nor g3809(n3876 ,n1026 ,n3765);
    or g3810(n3875 ,n2784 ,n3651);
    nor g3811(n3874 ,n1033 ,n3371);
    or g3812(n3873 ,n2646 ,n3657);
    or g3813(n3872 ,n2333 ,n3674);
    or g3814(n3871 ,n2866 ,n3672);
    nor g3815(n3870 ,n2984 ,n3548);
    nor g3816(n3869 ,n1033 ,n3384);
    or g3817(n3868 ,n2647 ,n3689);
    or g3818(n3867 ,n2329 ,n3670);
    nor g3819(n3866 ,n1033 ,n3375);
    or g3820(n3865 ,n3758 ,n2636);
    or g3821(n3864 ,n2858 ,n3669);
    nor g3822(n3863 ,n1033 ,n3376);
    or g3823(n3862 ,n2720 ,n3668);
    or g3824(n3861 ,n2864 ,n3667);
    or g3825(n3860 ,n2799 ,n3690);
    nor g3826(n3859 ,n1033 ,n3377);
    nor g3827(n3858 ,n1033 ,n3380);
    nor g3828(n3857 ,n1033 ,n3378);
    nor g3829(n3856 ,n1033 ,n3357);
    or g3830(n3855 ,n2336 ,n3663);
    nor g3831(n3854 ,n3012 ,n3529);
    or g3832(n3853 ,n2650 ,n3735);
    nor g3833(n3852 ,n1033 ,n3409);
    nor g3834(n3851 ,n2983 ,n3525);
    nor g3835(n3850 ,n2371 ,n3570);
    or g3836(n3849 ,n2712 ,n3664);
    nor g3837(n3848 ,n3488 ,n3745);
    nor g3838(n3847 ,n1[63] ,n3524);
    nor g3839(n3846 ,n2980 ,n3522);
    or g3840(n3845 ,n2341 ,n3661);
    nor g3841(n3844 ,n1[62] ,n3519);
    or g3842(n3843 ,n1678 ,n3666);
    nor g3843(n3842 ,n2997 ,n3517);
    or g3844(n3841 ,n2244 ,n3739);
    or g3845(n3840 ,n2340 ,n3660);
    or g3846(n3839 ,n2717 ,n3635);
    nor g3847(n3838 ,n1[61] ,n3515);
    nor g3848(n3837 ,n3018 ,n3512);
    nor g3849(n3836 ,n1[60] ,n3514);
    or g3850(n3835 ,n2342 ,n3659);
    or g3851(n3834 ,n1728 ,n3636);
    nor g3852(n3833 ,n3314 ,n3755);
    nor g3853(n3832 ,n2981 ,n3506);
    nor g3854(n3831 ,n2977 ,n3503);
    or g3855(n3830 ,n2658 ,n3637);
    nor g3856(n3829 ,n3332 ,n3733);
    nor g3857(n3828 ,n3010 ,n3499);
    or g3858(n3827 ,n2661 ,n3695);
    or g3859(n3826 ,n2520 ,n3720);
    nor g3860(n3825 ,n3009 ,n3493);
    nor g3861(n3824 ,n2002 ,n3495);
    nor g3862(n3823 ,n1[55] ,n3494);
    or g3863(n3822 ,n2638 ,n3697);
    nor g3864(n3821 ,n1[53] ,n3487);
    or g3865(n3820 ,n3088 ,n3742);
    nor g3866(n3819 ,n1[52] ,n3574);
    nor g3867(n3818 ,n2985 ,n3584);
    nor g3868(n3817 ,n3587 ,n3743);
    or g3869(n3816 ,n2662 ,n3698);
    or g3870(n3815 ,n2663 ,n3638);
    nor g3871(n3814 ,n3611 ,n3752);
    or g3872(n3813 ,n2664 ,n3639);
    or g3873(n3812 ,n3087 ,n3732);
    nor g3874(n3811 ,n3310 ,n3749);
    or g3875(n3810 ,n2688 ,n3653);
    nor g3876(n3809 ,n3526 ,n3751);
    or g3877(n3808 ,n2845 ,n3676);
    nor g3878(n3807 ,n3605 ,n3750);
    or g3879(n3806 ,n1632 ,n3640);
    or g3880(n3805 ,n2687 ,n3652);
    nor g3881(n3804 ,n3345 ,n3731);
    or g3882(n3803 ,n2640 ,n3631);
    nor g3883(n3802 ,n3338 ,n3748);
    nor g3884(n3801 ,n3337 ,n3747);
    or g3885(n3800 ,n2699 ,n3649);
    or g3886(n3799 ,n2795 ,n3648);
    nor g3887(n3798 ,n3333 ,n3746);
    or g3888(n3797 ,n2681 ,n3736);
    nor g3889(n3796 ,n3622 ,n3740);
    or g3890(n3795 ,n3089 ,n3738);
    nor g3891(n3794 ,n1[35] ,n3280);
    or g3892(n3793 ,n2709 ,n3641);
    or g3893(n3792 ,n2243 ,n3741);
    or g3894(n3791 ,n2324 ,n3645);
    nor g3895(n3790 ,n3327 ,n3756);
    nor g3896(n3789 ,n2373 ,n3628);
    or g3897(n3788 ,n2855 ,n3702);
    nor g3898(n3787 ,n3325 ,n3744);
    or g3899(n3786 ,n2652 ,n3644);
    or g3900(n3785 ,n1677 ,n3643);
    or g3901(n3784 ,n2767 ,n3704);
    or g3902(n3783 ,n1644 ,n3642);
    nor g3903(n3782 ,n1033 ,n3356);
    or g3904(n3781 ,n1675 ,n3630);
    or g3905(n3780 ,n2785 ,n3634);
    nor g3906(n4001 ,n7399 ,n3364);
    nor g3907(n4000 ,n7399 ,n3372);
    nor g3908(n3999 ,n1033 ,n3374);
    nor g3909(n3998 ,n1033 ,n3365);
    nor g3910(n3997 ,n7399 ,n3377);
    nor g3911(n3996 ,n7399 ,n3376);
    nor g3912(n3995 ,n7399 ,n3380);
    nor g3913(n3994 ,n7399 ,n3409);
    nor g3914(n3993 ,n7399 ,n3375);
    nor g3915(n3992 ,n7399 ,n3384);
    nor g3916(n3991 ,n7399 ,n3374);
    nor g3917(n3990 ,n7399 ,n3382);
    nor g3918(n3989 ,n7399 ,n3385);
    nor g3919(n3988 ,n7399 ,n3373);
    nor g3920(n3987 ,n7399 ,n3383);
    nor g3921(n3986 ,n7399 ,n3386);
    nor g3922(n3985 ,n7399 ,n3371);
    nor g3923(n3984 ,n1033 ,n3368);
    nor g3924(n3983 ,n7399 ,n3370);
    nor g3925(n3982 ,n7399 ,n3379);
    nor g3926(n3981 ,n7399 ,n3369);
    nor g3927(n3980 ,n7399 ,n3355);
    nor g3928(n3979 ,n1033 ,n3383);
    nor g3929(n3978 ,n7399 ,n3367);
    nor g3930(n3977 ,n1033 ,n3372);
    nor g3931(n3976 ,n7399 ,n3366);
    nor g3932(n3975 ,n7399 ,n3365);
    nor g3933(n3974 ,n7399 ,n3378);
    nor g3934(n3973 ,n1033 ,n3386);
    xnor g3935(n3972 ,n2528 ,n2837);
    nor g3936(n3971 ,n1033 ,n3370);
    nor g3937(n3970 ,n7399 ,n3363);
    nor g3938(n3969 ,n7399 ,n3361);
    nor g3939(n3968 ,n1033 ,n3361);
    nor g3940(n3967 ,n1033 ,n3359);
    nor g3941(n3966 ,n7399 ,n3359);
    nor g3942(n3965 ,n1033 ,n3358);
    nor g3943(n3964 ,n1033 ,n3355);
    nor g3944(n3963 ,n7399 ,n3358);
    nor g3945(n3962 ,n7399 ,n3357);
    nor g3946(n3961 ,n7399 ,n3356);
    xnor g3947(n3960 ,n2540 ,n2835);
    xnor g3948(n3959 ,n2534 ,n2825);
    xnor g3949(n3958 ,n2537 ,n2828);
    xnor g3950(n3957 ,n2542 ,n2829);
    xnor g3951(n3956 ,n2529 ,n2827);
    xnor g3952(n3955 ,n2530 ,n2832);
    xnor g3953(n3954 ,n2532 ,n2833);
    xnor g3954(n3953 ,n2539 ,n2834);
    xnor g3955(n3952 ,n2531 ,n2838);
    xnor g3956(n3951 ,n2536 ,n2836);
    nor g3957(n3950 ,n7399 ,n3360);
    nor g3958(n3949 ,n7399 ,n3368);
    nor g3959(n3948 ,n7399 ,n3362);
    xnor g3960(n3946 ,n2830 ,n2535);
    xnor g3961(n3944 ,n2831 ,n2541);
    xnor g3962(n3942 ,n2826 ,n2533);
    or g3963(n3763 ,n2763 ,n2846);
    or g3964(n3762 ,n7344 ,n2729);
    nor g3965(n3761 ,n1137 ,n2848);
    nor g3966(n3760 ,n1128 ,n2779);
    nor g3967(n3759 ,n1298 ,n2852);
    nor g3968(n3758 ,n1288 ,n2791);
    nor g3969(n3757 ,n1144 ,n3045);
    nor g3970(n3756 ,n1296 ,n3099);
    nor g3971(n3755 ,n1132 ,n3111);
    or g3972(n3754 ,n1125 ,n3132);
    or g3973(n3753 ,n1130 ,n3119);
    nor g3974(n3752 ,n1129 ,n3150);
    nor g3975(n3751 ,n1286 ,n3123);
    nor g3976(n3750 ,n1285 ,n3097);
    nor g3977(n3749 ,n1292 ,n3126);
    nor g3978(n3748 ,n1143 ,n3139);
    nor g3979(n3747 ,n1287 ,n3145);
    nor g3980(n3746 ,n1134 ,n3141);
    nor g3981(n3745 ,n1141 ,n3103);
    nor g3982(n3744 ,n1142 ,n3130);
    nor g3983(n3743 ,n1258 ,n3095);
    nor g3984(n3742 ,n1253 ,n2890);
    nor g3985(n3741 ,n1103 ,n3019);
    nor g3986(n3740 ,n1105 ,n3149);
    nor g3987(n3739 ,n1088 ,n2996);
    nor g3988(n3738 ,n1086 ,n2895);
    nor g3989(n3737 ,n2001 ,n3054);
    nor g3990(n3736 ,n2372 ,n3071);
    nor g3991(n3735 ,n2370 ,n3091);
    nor g3992(n3734 ,n1079 ,n2909);
    nor g3993(n3733 ,n1236 ,n3138);
    nor g3994(n3732 ,n1236 ,n2891);
    nor g3995(n3731 ,n1228 ,n3125);
    nor g3996(n3730 ,n1716 ,n2758);
    nor g3997(n3729 ,n1717 ,n2756);
    nor g3998(n3728 ,n1718 ,n2754);
    nor g3999(n3727 ,n2039 ,n3120);
    nor g4000(n3726 ,n2048 ,n3104);
    nor g4001(n3725 ,n1741 ,n3092);
    nor g4002(n3724 ,n2045 ,n3108);
    nor g4003(n3723 ,n1744 ,n3093);
    nor g4004(n3722 ,n1724 ,n2706);
    or g4005(n3721 ,n2589 ,n2637);
    nor g4006(n3720 ,n0[120] ,n2587);
    nor g4007(n3719 ,n1[54] ,n3067);
    nor g4008(n3718 ,n1598 ,n3094);
    nor g4009(n3717 ,n1719 ,n2696);
    or g4010(n3716 ,n2543 ,n2693);
    or g4011(n3715 ,n2583 ,n2691);
    nor g4012(n3714 ,n1722 ,n2690);
    nor g4013(n3713 ,n1[43] ,n3083);
    or g4014(n3712 ,n2566 ,n2683);
    nor g4015(n3711 ,n2023 ,n3124);
    nor g4016(n3710 ,n1720 ,n2677);
    nor g4017(n3709 ,n2005 ,n3102);
    nor g4018(n3708 ,n2019 ,n3144);
    nor g4019(n3707 ,n2059 ,n3106);
    nor g4020(n3706 ,n1721 ,n2694);
    nor g4021(n3705 ,n2053 ,n3110);
    nor g4022(n3704 ,n2042 ,n3112);
    nor g4023(n3703 ,n2025 ,n3140);
    nor g4024(n3702 ,n2051 ,n3114);
    nor g4025(n3701 ,n2062 ,n3122);
    nor g4026(n3700 ,n2009 ,n3116);
    nor g4027(n3699 ,n2011 ,n3129);
    nor g4028(n3698 ,n2013 ,n3118);
    nor g4029(n3697 ,n2082 ,n3096);
    nor g4030(n3696 ,n2077 ,n3135);
    nor g4031(n3695 ,n2015 ,n3133);
    nor g4032(n3694 ,n1723 ,n2660);
    nor g4033(n3693 ,n2021 ,n3151);
    nor g4034(n3692 ,n0[14] ,n2840);
    nor g4035(n3691 ,n2093 ,n3098);
    nor g4036(n3690 ,n2007 ,n3127);
    nor g4037(n3689 ,n2027 ,n3137);
    nor g4038(n3688 ,n2057 ,n3146);
    nor g4039(n3687 ,n2029 ,n3142);
    nor g4040(n3686 ,n2080 ,n3148);
    nor g4041(n3685 ,n2055 ,n3100);
    nor g4042(n3684 ,n2037 ,n3131);
    nor g4043(n3683 ,n1064 ,n2625);
    or g4044(n3682 ,n7341 ,n2656);
    nor g4045(n3681 ,n2419 ,n1060);
    nor g4046(n3680 ,n2409 ,n1060);
    nor g4047(n3679 ,n2390 ,n1060);
    nor g4048(n3678 ,n2391 ,n1060);
    nor g4049(n3677 ,n2420 ,n1060);
    nor g4050(n3676 ,n2408 ,n1057);
    nor g4051(n3675 ,n2412 ,n1060);
    nor g4052(n3674 ,n2428 ,n1057);
    nor g4053(n3673 ,n2432 ,n1057);
    nor g4054(n3672 ,n2433 ,n1060);
    nor g4055(n3671 ,n2511 ,n1060);
    nor g4056(n3670 ,n2424 ,n1057);
    nor g4057(n3669 ,n2407 ,n1057);
    nor g4058(n3668 ,n2509 ,n1058);
    nor g4059(n3667 ,n2421 ,n1058);
    nor g4060(n3666 ,n2396 ,n1060);
    nor g4061(n3665 ,n2382 ,n1060);
    nor g4062(n3664 ,n2395 ,n1057);
    nor g4063(n3663 ,n2490 ,n1058);
    nor g4064(n3662 ,n2397 ,n1060);
    nor g4065(n3661 ,n2417 ,n1060);
    nor g4066(n3660 ,n2406 ,n1060);
    nor g4067(n3659 ,n2380 ,n1058);
    nor g4068(n3658 ,n2399 ,n1057);
    nor g4069(n3657 ,n2388 ,n1057);
    nor g4070(n3656 ,n2411 ,n1058);
    nor g4071(n3655 ,n2431 ,n1057);
    nor g4072(n3654 ,n2429 ,n1060);
    nor g4073(n3653 ,n2423 ,n1060);
    nor g4074(n3652 ,n2387 ,n1060);
    nor g4075(n3651 ,n2502 ,n1058);
    nor g4076(n3650 ,n2377 ,n1057);
    nor g4077(n3649 ,n2403 ,n1060);
    nor g4078(n3648 ,n2496 ,n1058);
    nor g4079(n3647 ,n2379 ,n1058);
    nor g4080(n3646 ,n2384 ,n1060);
    nor g4081(n3645 ,n2495 ,n1060);
    nor g4082(n3644 ,n2394 ,n1057);
    nor g4083(n3643 ,n2434 ,n1057);
    nor g4084(n3642 ,n2393 ,n1057);
    nor g4085(n3641 ,n2427 ,n1058);
    nor g4086(n3640 ,n2392 ,n1058);
    nor g4087(n3639 ,n2400 ,n1057);
    nor g4088(n3638 ,n2414 ,n1058);
    nor g4089(n3637 ,n2398 ,n1060);
    nor g4090(n3636 ,n2381 ,n1058);
    nor g4091(n3635 ,n2426 ,n1058);
    nor g4092(n3634 ,n2389 ,n1060);
    nor g4093(n3633 ,n2405 ,n1060);
    nor g4094(n3632 ,n2418 ,n1057);
    nor g4095(n3631 ,n2430 ,n1060);
    nor g4096(n3630 ,n2404 ,n1060);
    or g4097(n3629 ,n1053 ,n2896);
    nor g4098(n3628 ,n1050 ,n3138);
    or g4099(n3627 ,n2860 ,n2697);
    or g4100(n3626 ,n3076 ,n2760);
    or g4101(n3625 ,n2281 ,n2788);
    nor g4102(n3624 ,n1538 ,n2986);
    or g4103(n3623 ,n2335 ,n3055);
    nor g4104(n3622 ,n0[4] ,n3053);
    nor g4105(n3621 ,n1031 ,n2847);
    or g4106(n3620 ,n3109 ,n3002);
    or g4107(n3619 ,n2337 ,n2841);
    or g4108(n3618 ,n3077 ,n2761);
    nor g4109(n3617 ,n2885 ,n2822);
    nor g4110(n3616 ,n1031 ,n2849);
    or g4111(n3615 ,n3073 ,n2755);
    nor g4112(n3614 ,n1031 ,n2966);
    or g4113(n3613 ,n2908 ,n2644);
    or g4114(n3612 ,n2279 ,n2851);
    nor g4115(n3611 ,n1[47] ,n3057);
    nor g4116(n3610 ,n1031 ,n2943);
    nor g4117(n3609 ,n1031 ,n2853);
    or g4118(n3608 ,n2819 ,n2642);
    or g4119(n3607 ,n2285 ,n3080);
    or g4120(n3606 ,n2883 ,n2857);
    nor g4121(n3605 ,n1[44] ,n3060);
    or g4122(n3604 ,n2250 ,n3034);
    or g4123(n3603 ,n2750 ,n2878);
    or g4124(n3602 ,n2991 ,n2692);
    or g4125(n3601 ,n2278 ,n2882);
    nor g4126(n3600 ,n1031 ,n2959);
    or g4127(n3599 ,n2287 ,n3000);
    or g4128(n3598 ,n3074 ,n3020);
    or g4129(n3597 ,n3074 ,n2749);
    or g4130(n3596 ,n2280 ,n2748);
    or g4131(n3595 ,n2290 ,n2881);
    or g4132(n3594 ,n2880 ,n2888);
    or g4133(n3593 ,n2275 ,n2815);
    or g4134(n3592 ,n2747 ,n2892);
    or g4135(n3591 ,n2289 ,n2879);
    or g4136(n3590 ,n3084 ,n2695);
    or g4137(n3589 ,n2271 ,n2901);
    or g4138(n3588 ,n2746 ,n2893);
    nor g4139(n3587 ,n1[50] ,n3073);
    or g4140(n3586 ,n2277 ,n2877);
    or g4141(n3585 ,n2736 ,n2821);
    nor g4142(n3584 ,n2453 ,n2912);
    or g4143(n3583 ,n3086 ,n2742);
    or g4144(n3582 ,n2876 ,n2894);
    or g4145(n3581 ,n2322 ,n3062);
    nor g4146(n3580 ,n1528 ,n3011);
    or g4147(n3579 ,n2276 ,n2897);
    or g4148(n3578 ,n3117 ,n3030);
    or g4149(n3577 ,n2810 ,n2733);
    or g4150(n3576 ,n2875 ,n2898);
    nor g4151(n3575 ,n1031 ,n2950);
    nor g4152(n3574 ,n3056 ,n3043);
    nor g4153(n3573 ,n3128 ,n2766);
    or g4154(n3572 ,n2874 ,n2900);
    nor g4155(n3571 ,n1031 ,n2970);
    nor g4156(n3570 ,n1050 ,n3125);
    or g4157(n3569 ,n2269 ,n2872);
    or g4158(n3568 ,n2871 ,n2902);
    or g4159(n3567 ,n2338 ,n3057);
    or g4160(n3566 ,n2870 ,n2735);
    or g4161(n3565 ,n2713 ,n2998);
    or g4162(n3564 ,n2274 ,n2903);
    or g4163(n3563 ,n1[40] ,n3084);
    or g4164(n3562 ,n2283 ,n2839);
    or g4165(n3561 ,n2869 ,n2731);
    or g4166(n3560 ,n2266 ,n2812);
    nor g4167(n3559 ,n1031 ,n2967);
    or g4168(n3558 ,n2868 ,n2728);
    or g4169(n3557 ,n2288 ,n2910);
    or g4170(n3556 ,n3081 ,n2727);
    or g4171(n3555 ,n1694 ,n2771);
    or g4172(n3554 ,n2273 ,n2867);
    or g4173(n3553 ,n2726 ,n2911);
    or g4174(n3552 ,n2256 ,n2913);
    or g4175(n3551 ,n3016 ,n2725);
    or g4176(n3550 ,n2332 ,n2918);
    or g4177(n3549 ,n2331 ,n2923);
    nor g4178(n3548 ,n2451 ,n3087);
    or g4179(n3547 ,n2823 ,n2751);
    or g4180(n3546 ,n2873 ,n3035);
    or g4181(n3545 ,n2865 ,n2934);
    or g4182(n3544 ,n1637 ,n2700);
    or g4183(n3543 ,n2319 ,n3064);
    or g4184(n3542 ,n2328 ,n2939);
    or g4185(n3541 ,n2327 ,n3059);
    or g4186(n3540 ,n2326 ,n2942);
    or g4187(n3539 ,n2856 ,n2718);
    or g4188(n3538 ,n2297 ,n2765);
    or g4189(n3537 ,n3026 ,n2682);
    or g4190(n3536 ,n2974 ,n2743);
    or g4191(n3535 ,n2716 ,n2992);
    or g4192(n3534 ,n2304 ,n2863);
    or g4193(n3533 ,n2715 ,n2993);
    or g4194(n3532 ,n2739 ,n2889);
    or g4195(n3531 ,n2317 ,n2862);
    nor g4196(n3530 ,n1031 ,n2947);
    nor g4197(n3529 ,n2448 ,n2921);
    or g4198(n3528 ,n2861 ,n2714);
    or g4199(n3527 ,n2303 ,n2899);
    nor g4200(n3526 ,n1[45] ,n3059);
    nor g4201(n3525 ,n2486 ,n2920);
    nor g4202(n3524 ,n3058 ,n3050);
    nor g4203(n3523 ,n3101 ,n2994);
    nor g4204(n3522 ,n2444 ,n2919);
    or g4205(n3521 ,n3082 ,n2685);
    nor g4206(n3520 ,n3143 ,n2800);
    nor g4207(n3519 ,n3064 ,n3049);
    or g4208(n3518 ,n2270 ,n2999);
    nor g4209(n3517 ,n2442 ,n3089);
    nor g4210(n3516 ,n3105 ,n2781);
    nor g4211(n3515 ,n3062 ,n3047);
    nor g4212(n3514 ,n3055 ,n3048);
    nor g4213(n3513 ,n3107 ,n3001);
    nor g4214(n3512 ,n2457 ,n3088);
    or g4215(n3511 ,n2976 ,n3004);
    or g4216(n3510 ,n3078 ,n3022);
    or g4217(n3509 ,n2272 ,n3078);
    nor g4218(n3508 ,n1031 ,n2948);
    or g4219(n3507 ,n2265 ,n2705);
    nor g4220(n3506 ,n2461 ,n2916);
    or g4221(n3505 ,n3015 ,n2732);
    or g4222(n3504 ,n1[57] ,n3081);
    nor g4223(n3503 ,n2446 ,n2907);
    nor g4224(n3502 ,n3115 ,n2818);
    nor g4225(n3501 ,n2463 ,n2904);
    or g4226(n3500 ,n2704 ,n3025);
    nor g4227(n3499 ,n2459 ,n2915);
    nor g4228(n3498 ,n1519 ,n3007);
    or g4229(n3497 ,n2320 ,n3058);
    or g4230(n3496 ,n1666 ,n2703);
    nor g4231(n3495 ,n1050 ,n3149);
    nor g4232(n3494 ,n3065 ,n3044);
    nor g4233(n3493 ,n2455 ,n2914);
    or g4234(n3492 ,n1631 ,n2701);
    or g4235(n3491 ,n3079 ,n2666);
    nor g4236(n3490 ,n3121 ,n3027);
    or g4237(n3489 ,n2284 ,n3029);
    nor g4238(n3488 ,n1[34] ,n3072);
    nor g4239(n3487 ,n3068 ,n3042);
    nor g4240(n3486 ,n1064 ,n2937);
    or g4241(n3779 ,n1389 ,n2925);
    or g4242(n3778 ,n1444 ,n2926);
    or g4243(n3777 ,n1429 ,n2927);
    or g4244(n3776 ,n1438 ,n2928);
    or g4245(n3775 ,n1372 ,n2929);
    or g4246(n3774 ,n1464 ,n2931);
    or g4247(n3773 ,n1407 ,n2932);
    or g4248(n3772 ,n1388 ,n2933);
    or g4249(n3771 ,n1435 ,n2935);
    or g4250(n3770 ,n1427 ,n2936);
    or g4251(n3769 ,n1391 ,n2940);
    or g4252(n3768 ,n1417 ,n2941);
    nor g4253(n3767 ,n1361 ,n2973);
    nor g4254(n3766 ,n1479 ,n2930);
    nor g4255(n3765 ,n1378 ,n2924);
    nor g4256(n3764 ,n1392 ,n2938);
    not g4257(n3485 ,n3484);
    not g4258(n3483 ,n3482);
    not g4259(n3481 ,n3480);
    not g4260(n3479 ,n3478);
    not g4261(n3477 ,n3476);
    not g4262(n3475 ,n3474);
    not g4263(n3473 ,n3472);
    not g4264(n3471 ,n3470);
    not g4265(n3469 ,n3468);
    not g4266(n3467 ,n3466);
    not g4267(n3465 ,n3464);
    not g4268(n3463 ,n3462);
    not g4269(n3461 ,n3460);
    not g4270(n3459 ,n3458);
    not g4271(n3457 ,n3456);
    not g4272(n3455 ,n3454);
    not g4273(n3453 ,n3452);
    not g4274(n3451 ,n3450);
    not g4275(n3449 ,n3448);
    not g4276(n3447 ,n3446);
    not g4277(n3445 ,n3444);
    not g4278(n3443 ,n3442);
    not g4279(n3441 ,n3440);
    not g4280(n3439 ,n3438);
    not g4281(n3437 ,n3436);
    not g4282(n3435 ,n3434);
    not g4283(n3433 ,n3432);
    not g4284(n3431 ,n3430);
    not g4285(n3429 ,n3428);
    not g4286(n3427 ,n3426);
    not g4287(n3425 ,n3424);
    not g4288(n3423 ,n3422);
    not g4289(n3421 ,n3420);
    not g4290(n3419 ,n3418);
    not g4291(n3417 ,n3416);
    not g4292(n3415 ,n3414);
    not g4293(n3413 ,n3412);
    not g4294(n3411 ,n3410);
    not g4295(n3352 ,n3353);
    or g4296(n3351 ,n2325 ,n3061);
    nor g4297(n3350 ,n1031 ,n2944);
    nor g4298(n3349 ,n1525 ,n3006);
    nor g4299(n3348 ,n3134 ,n2769);
    nor g4300(n3347 ,n1031 ,n2772);
    or g4301(n3346 ,n1661 ,n2686);
    nor g4302(n3345 ,n0[10] ,n3090);
    or g4303(n3344 ,n3046 ,n2684);
    or g4304(n3343 ,n3051 ,n2711);
    nor g4305(n3342 ,n1521 ,n3008);
    or g4306(n3341 ,n3136 ,n2824);
    or g4307(n3340 ,n3076 ,n3021);
    nor g4308(n3339 ,n1541 ,n2982);
    nor g4309(n3338 ,n1[39] ,n3061);
    nor g4310(n3337 ,n1[38] ,n3063);
    or g4311(n3336 ,n2305 ,n3069);
    or g4312(n3335 ,n2299 ,n3063);
    nor g4313(n3334 ,n1530 ,n2979);
    nor g4314(n3333 ,n1[37] ,n3069);
    nor g4315(n3332 ,n0[24] ,n3070);
    or g4316(n3331 ,n1636 ,n2797);
    or g4317(n3330 ,n2816 ,n2679);
    nor g4318(n3329 ,n3147 ,n2780);
    or g4319(n3328 ,n3023 ,n2814);
    nor g4320(n3327 ,n1[33] ,n3080);
    nor g4321(n3326 ,n1534 ,n2975);
    nor g4322(n3325 ,n1[32] ,n3085);
    or g4323(n3324 ,n2811 ,n2676);
    or g4324(n3323 ,n1652 ,n2770);
    or g4325(n3322 ,n3075 ,n2675);
    nor g4326(n3321 ,n1031 ,n2956);
    or g4327(n3320 ,n2298 ,n2786);
    nor g4328(n3319 ,n1031 ,n2969);
    or g4329(n3318 ,n2809 ,n2673);
    nor g4330(n3317 ,n1031 ,n2955);
    nor g4331(n3316 ,n1031 ,n2957);
    or g4332(n3315 ,n1700 ,n2906);
    nor g4333(n3314 ,n1[58] ,n3077);
    or g4334(n3313 ,n3113 ,n3024);
    nor g4335(n3312 ,n1552 ,n2978);
    or g4336(n3311 ,n1651 ,n2808);
    nor g4337(n3310 ,n1[41] ,n3079);
    nor g4338(n3309 ,n1031 ,n2965);
    or g4339(n3308 ,n3072 ,n2670);
    or g4340(n3307 ,n2241 ,n2995);
    or g4341(n3306 ,n1619 ,n2669);
    or g4342(n3305 ,n2296 ,n2807);
    or g4343(n3304 ,n1650 ,n2752);
    or g4344(n3303 ,n1640 ,n2649);
    or g4345(n3302 ,n2817 ,n2667);
    or g4346(n3301 ,n2645 ,n2805);
    or g4347(n3300 ,n2804 ,n2665);
    or g4348(n3299 ,n3086 ,n3013);
    or g4349(n3298 ,n1672 ,n2802);
    nor g4350(n3297 ,n1031 ,n2953);
    or g4351(n3296 ,n1641 ,n2801);
    nor g4352(n3295 ,n1031 ,n2952);
    or g4353(n3294 ,n3085 ,n2657);
    nor g4354(n3293 ,n1031 ,n2951);
    or g4355(n3292 ,n1674 ,n3031);
    or g4356(n3291 ,n2306 ,n2798);
    or g4357(n3290 ,n1707 ,n2905);
    or g4358(n3289 ,n1711 ,n2794);
    or g4359(n3288 ,n1708 ,n2793);
    or g4360(n3287 ,n3066 ,n2796);
    or g4361(n3286 ,n2790 ,n2655);
    or g4362(n3285 ,n2318 ,n2843);
    or g4363(n3284 ,n1671 ,n2789);
    nor g4364(n3283 ,n1031 ,n2949);
    nor g4365(n3282 ,n1031 ,n2958);
    or g4366(n3281 ,n2653 ,n2787);
    nor g4367(n3280 ,n3075 ,n2988);
    nor g4368(n3279 ,n1031 ,n2964);
    or g4369(n3278 ,n2990 ,n2668);
    nor g4370(n3277 ,n1031 ,n2954);
    nor g4371(n3276 ,n1031 ,n2945);
    or g4372(n3275 ,n3036 ,n2654);
    nor g4373(n3274 ,n1031 ,n2960);
    or g4374(n3273 ,n2842 ,n2783);
    nor g4375(n3272 ,n1031 ,n2946);
    or g4376(n3271 ,n1633 ,n2782);
    nor g4377(n3270 ,n1031 ,n2968);
    or g4378(n3269 ,n1630 ,n2778);
    or g4379(n3268 ,n1696 ,n2854);
    or g4380(n3267 ,n1688 ,n2776);
    or g4381(n3266 ,n3068 ,n2775);
    or g4382(n3265 ,n1663 ,n2672);
    or g4383(n3264 ,n1660 ,n2671);
    nor g4384(n3263 ,n1031 ,n2963);
    or g4385(n3262 ,n2639 ,n2806);
    nor g4386(n3261 ,n1031 ,n2961);
    nor g4387(n3260 ,n1031 ,n2962);
    or g4388(n3259 ,n2745 ,n2768);
    or g4389(n3258 ,n2286 ,n2850);
    or g4390(n3257 ,n1647 ,n2698);
    or g4391(n3256 ,n2859 ,n2648);
    nor g4392(n3255 ,n2245 ,n2578);
    xnor g4393(n3484 ,n2143 ,n2086);
    xnor g4394(n3254 ,n2002 ,n2204);
    xnor g4395(n3253 ,n1804 ,n2112);
    xnor g4396(n3482 ,n2164 ,n2087);
    xnor g4397(n3480 ,n2140 ,n2435);
    xnor g4398(n3252 ,n1[108] ,n2093);
    xnor g4399(n3251 ,n2199 ,n2095);
    xnor g4400(n3250 ,n1[110] ,n2016);
    xnor g4401(n3249 ,n2200 ,n2040);
    xnor g4402(n3248 ,n2202 ,n2030);
    xnor g4403(n3247 ,n1[123] ,n2053);
    xnor g4404(n3246 ,n2142 ,n2003);
    xnor g4405(n3245 ,n1[112] ,n2039);
    xnor g4406(n3244 ,n2203 ,n2129);
    xnor g4407(n3243 ,n2171 ,n2410);
    xnor g4408(n3478 ,n1759 ,n2135);
    xnor g4409(n3242 ,n2429 ,n2403);
    xnor g4410(n3241 ,n1[114] ,n2082);
    xnor g4411(n3240 ,n2431 ,n2377);
    xnor g4412(n3239 ,n2173 ,n2422);
    xnor g4413(n3238 ,n2032 ,n2094);
    xnor g4414(n3237 ,n1[121] ,n2051);
    xnor g4415(n3236 ,n1[122] ,n2042);
    xnor g4416(n3235 ,n2186 ,n2386);
    xnor g4417(n3234 ,n1[124] ,n2045);
    xnor g4418(n3476 ,n1[125] ,n2059);
    xnor g4419(n3474 ,n1799 ,n2131);
    xnor g4420(n3233 ,n2380 ,n2387);
    xnor g4421(n3472 ,n1793 ,n2097);
    xnor g4422(n3232 ,n2434 ,n2392);
    xnor g4423(n3470 ,n1[127] ,n2005);
    xnor g4424(n3231 ,n2035 ,n2101);
    xnor g4425(n3230 ,n1[117] ,n2009);
    xnor g4426(n3229 ,n1[100] ,n1861);
    xnor g4427(n3228 ,n2388 ,n2397);
    xnor g4428(n3468 ,n2169 ,n2480);
    xnor g4429(n3227 ,n2412 ,n2408);
    xnor g4430(n3226 ,n4[26] ,n2085);
    xnor g4431(n3466 ,n2104 ,n2089);
    xnor g4432(n3464 ,n1801 ,n2133);
    xnor g4433(n3225 ,n1775 ,n2031);
    xnor g4434(n3224 ,n1[118] ,n2062);
    xnor g4435(n3223 ,n1776 ,n2032);
    xnor g4436(n3222 ,n1[104] ,n2027);
    xnor g4437(n3221 ,n1777 ,n2034);
    xnor g4438(n3220 ,n2394 ,n2399);
    xnor g4439(n3462 ,n1778 ,n2033);
    xnor g4440(n3219 ,n2174 ,n2482);
    xnor g4441(n3460 ,n2183 ,n2091);
    xnor g4442(n3218 ,n1[101] ,n2029);
    xnor g4443(n3217 ,n1[106] ,n1859);
    xnor g4444(n3458 ,n2170 ,n2046);
    xnor g4445(n3216 ,n2159 ,n2098);
    xnor g4446(n3215 ,n1765 ,n2035);
    xnor g4447(n3214 ,n1[115] ,n2013);
    xnor g4448(n3213 ,n1779 ,n2078);
    xnor g4449(n3212 ,n1781 ,n2043);
    xnor g4450(n3211 ,n4[21] ,n2064);
    xnor g4451(n3210 ,n2191 ,n2100);
    xnor g4452(n3456 ,n2151 ,n2084);
    xnor g4453(n3454 ,n2141 ,n2066);
    xnor g4454(n3452 ,n2185 ,n2083);
    xnor g4455(n3450 ,n2175 ,n2089);
    xnor g4456(n3209 ,n2206 ,n2102);
    xnor g4457(n3208 ,n2192 ,n2468);
    xnor g4458(n3207 ,n4[17] ,n2378);
    xnor g4459(n3206 ,n2153 ,n2472);
    xnor g4460(n3448 ,n2207 ,n2107);
    xnor g4461(n3205 ,n4[29] ,n2072);
    xnor g4462(n3446 ,n2208 ,n2103);
    xnor g4463(n3444 ,n2209 ,n2105);
    xnor g4464(n3204 ,n2040 ,n2109);
    xnor g4465(n3442 ,n2162 ,n2466);
    xnor g4466(n3440 ,n2156 ,n2481);
    xnor g4467(n3203 ,n1[105] ,n2007);
    xnor g4468(n3438 ,n2163 ,n2470);
    xnor g4469(n3436 ,n1753 ,n2147);
    xnor g4470(n3202 ,n2030 ,n2118);
    xnor g4471(n3434 ,n1[126] ,n2019);
    xnor g4472(n3432 ,n2210 ,n2106);
    xnor g4473(n3430 ,n2117 ,n2003);
    xnor g4474(n3428 ,n1876 ,n2146);
    xnor g4475(n3426 ,n2201 ,n2485);
    xnor g4476(n3424 ,n1[96] ,n2037);
    xnor g4477(n3422 ,n2165 ,n2483);
    xnor g4478(n3420 ,n2138 ,n2096);
    xnor g4479(n3201 ,n1762 ,n2063);
    xnor g4480(n3200 ,n2119 ,n2410);
    xnor g4481(n3199 ,n2176 ,n2065);
    xnor g4482(n3198 ,n1[107] ,n2077);
    xnor g4483(n3197 ,n2166 ,n2401);
    xnor g4484(n3196 ,n1[99] ,n2080);
    xnor g4485(n3195 ,n1[102] ,n2057);
    xnor g4486(n3194 ,n1[111] ,n2021);
    xnor g4487(n3193 ,n1805 ,n2075);
    xnor g4488(n3192 ,n1[113] ,n2015);
    xnor g4489(n3191 ,n1772 ,n2074);
    xnor g4490(n3190 ,n1[109] ,n2023);
    xnor g4491(n3189 ,n1[98] ,n2048);
    xnor g4492(n3418 ,n2139 ,n2145);
    xnor g4493(n3416 ,n1869 ,n2160);
    xnor g4494(n3188 ,n2423 ,n2379);
    xnor g4495(n3187 ,n2419 ,n2433);
    xnor g4496(n3186 ,n2400 ,n2426);
    xnor g4497(n3185 ,n1[103] ,n2025);
    xnor g4498(n3184 ,n1808 ,n2088);
    xnor g4499(n3414 ,n1809 ,n2070);
    xnor g4500(n3183 ,n2390 ,n2424);
    xnor g4501(n3182 ,n1782 ,n2069);
    xnor g4502(n3412 ,n2158 ,n2114);
    xnor g4503(n3181 ,n2189 ,n2113);
    xnor g4504(n3180 ,n1761 ,n2123);
    xnor g4505(n3179 ,n2391 ,n2407);
    xnor g4506(n3178 ,n2420 ,n2421);
    xnor g4507(n3410 ,n2187 ,n2067);
    xnor g4508(n3177 ,n2168 ,n2383);
    xnor g4509(n3176 ,n4[23] ,n2000);
    xnor g4510(n3175 ,n0[54] ,n2417);
    xnor g4511(n3174 ,n1[116] ,n2011);
    xnor g4512(n3173 ,n1[119] ,n1766);
    xnor g4513(n3172 ,n1[120] ,n1774);
    xnor g4514(n3171 ,n0[53] ,n2406);
    xnor g4515(n3170 ,n4[18] ,n2049);
    xnor g4516(n3169 ,n0[52] ,n2384);
    xnor g4517(n3168 ,n0[55] ,n2395);
    xnor g4518(n3167 ,n0[104] ,n1752);
    xnor g4519(n3166 ,n1[97] ,n2055);
    xnor g4520(n3165 ,n4[24] ,n2373);
    xnor g4521(n3164 ,n0[125] ,n1828);
    xnor g4522(n3163 ,n0[102] ,n2155);
    xnor g4523(n3162 ,n0[126] ,n1833);
    xnor g4524(n3161 ,n0[101] ,n2177);
    xnor g4525(n3160 ,n0[119] ,n2432);
    xnor g4526(n3159 ,n0[124] ,n1834);
    xnor g4527(n3158 ,n0[127] ,n1835);
    xnor g4528(n3157 ,n0[77] ,n2428);
    xnor g4529(n3156 ,n0[76] ,n2382);
    xnor g4530(n3155 ,n0[78] ,n2389);
    xnor g4531(n3154 ,n0[118] ,n2427);
    xnor g4532(n3153 ,n0[117] ,n2411);
    xnor g4533(n3152 ,n0[79] ,n2418);
    xnor g4534(n3409 ,n1768 ,n1746);
    xnor g4535(n3408 ,n0[117] ,n1810);
    xnor g4536(n3407 ,n0[110] ,n1840);
    xnor g4537(n3406 ,n0[118] ,n1824);
    xnor g4538(n3405 ,n0[109] ,n1838);
    xnor g4539(n3404 ,n0[108] ,n1837);
    xnor g4540(n3403 ,n0[103] ,n1829);
    xnor g4541(n3402 ,n0[70] ,n1842);
    xnor g4542(n3401 ,n0[116] ,n1827);
    xnor g4543(n3400 ,n0[100] ,n1831);
    xnor g4544(n3399 ,n0[101] ,n1830);
    xnor g4545(n3398 ,n0[119] ,n1798);
    xnor g4546(n3397 ,n0[90] ,n1848);
    xnor g4547(n3396 ,n0[105] ,n1844);
    xnor g4548(n3395 ,n0[81] ,n1843);
    xnor g4549(n3394 ,n0[114] ,n1852);
    xnor g4550(n3393 ,n0[72] ,n1851);
    xnor g4551(n3392 ,n0[115] ,n1849);
    xnor g4552(n3391 ,n0[75] ,n1847);
    xnor g4553(n3390 ,n0[123] ,n1845);
    xnor g4554(n3389 ,n0[112] ,n1853);
    xnor g4555(n3388 ,n0[121] ,n1850);
    xnor g4556(n3387 ,n0[120] ,n1846);
    xnor g4557(n3386 ,n1879 ,n1855);
    xnor g4558(n3385 ,n1860 ,n1826);
    xnor g4559(n3384 ,n1817 ,n1816);
    xnor g4560(n3383 ,n1786 ,n1771);
    xnor g4561(n3382 ,n1878 ,n1747);
    xnor g4562(n3381 ,n0[111] ,n1841);
    xnor g4563(n3380 ,n1867 ,n1870);
    xnor g4564(n3379 ,n1749 ,n1751);
    xnor g4565(n3378 ,n1811 ,n1871);
    xnor g4566(n3377 ,n1836 ,n1832);
    xnor g4567(n3376 ,n1873 ,n1814);
    xnor g4568(n3375 ,n1821 ,n1854);
    xnor g4569(n3374 ,n1760 ,n1792);
    xnor g4570(n3373 ,n1818 ,n1857);
    xnor g4571(n3372 ,n1789 ,n1877);
    xnor g4572(n3371 ,n1815 ,n1820);
    xnor g4573(n3370 ,n1806 ,n1866);
    xnor g4574(n3369 ,n1797 ,n1868);
    xnor g4575(n3368 ,n1823 ,n1795);
    xnor g4576(n3367 ,n1865 ,n1858);
    xnor g4577(n3366 ,n1791 ,n1875);
    xnor g4578(n3365 ,n1874 ,n1784);
    xnor g4579(n3364 ,n1788 ,n1790);
    xnor g4580(n3363 ,n1783 ,n1780);
    xnor g4581(n3362 ,n1769 ,n1802);
    xnor g4582(n3361 ,n1773 ,n1864);
    xnor g4583(n3360 ,n1785 ,n1748);
    xnor g4584(n3359 ,n1770 ,n1807);
    xnor g4585(n3358 ,n1822 ,n1764);
    xnor g4586(n3357 ,n1767 ,n1763);
    xnor g4587(n3356 ,n1757 ,n1794);
    xnor g4588(n3355 ,n1856 ,n1862);
    xnor g4589(n3354 ,n7676 ,n2148);
    nor g4590(n3353 ,n1031 ,n1059);
    not g4591(n3151 ,n3150);
    not g4592(n3148 ,n3147);
    not g4593(n3146 ,n3145);
    not g4594(n3144 ,n3143);
    not g4595(n3142 ,n3141);
    not g4596(n3140 ,n3139);
    not g4597(n3137 ,n3136);
    not g4598(n3135 ,n3134);
    not g4599(n3133 ,n3132);
    not g4600(n3131 ,n3130);
    not g4601(n3129 ,n3128);
    not g4602(n3127 ,n3126);
    not g4603(n3124 ,n3123);
    not g4604(n3122 ,n3121);
    not g4605(n3120 ,n3119);
    not g4606(n3118 ,n3117);
    not g4607(n3116 ,n3115);
    not g4608(n3114 ,n3113);
    not g4609(n3112 ,n3111);
    not g4610(n3110 ,n3109);
    not g4611(n3108 ,n3107);
    not g4612(n3106 ,n3105);
    not g4613(n3104 ,n3103);
    not g4614(n3102 ,n3101);
    not g4615(n3100 ,n3099);
    not g4616(n3098 ,n3097);
    not g4617(n3096 ,n3095);
    not g4618(n3091 ,n3090);
    not g4619(n3083 ,n3082);
    not g4620(n3071 ,n3070);
    not g4621(n3067 ,n3066);
    not g4622(n3054 ,n3053);
    not g4623(n1061 ,n3052);
    not g4624(n1058 ,n1059);
    not g4625(n1057 ,n1059);
    not g4626(n1059 ,n1060);
    nor g4627(n3051 ,n1048 ,n2481);
    nor g4628(n3050 ,n1149 ,n2367);
    nor g4629(n3049 ,n1148 ,n1051);
    nor g4630(n3048 ,n1301 ,n2367);
    nor g4631(n3047 ,n1304 ,n1049);
    nor g4632(n3046 ,n1049 ,n2466);
    or g4633(n3045 ,n0[119] ,n2367);
    nor g4634(n3044 ,n1289 ,n1048);
    nor g4635(n3043 ,n1291 ,n1051);
    nor g4636(n3042 ,n1138 ,n1049);
    nor g4637(n3041 ,n1545 ,n2513);
    nor g4638(n3040 ,n1547 ,n2515);
    nor g4639(n3039 ,n1548 ,n2517);
    nor g4640(n3038 ,n1048 ,n2095);
    nor g4641(n3037 ,n1051 ,n2103);
    nor g4642(n3036 ,n1051 ,n2102);
    nor g4643(n3035 ,n1051 ,n2100);
    nor g4644(n3034 ,n2367 ,n2214);
    nor g4645(n3033 ,n0[49] ,n1049);
    nor g4646(n3032 ,n1051 ,n2225);
    nor g4647(n3031 ,n1049 ,n2374);
    nor g4648(n3030 ,n0[51] ,n2367);
    nor g4649(n3029 ,n2367 ,n2475);
    nor g4650(n3028 ,n1[54] ,n1051);
    nor g4651(n3027 ,n0[54] ,n1051);
    nor g4652(n3026 ,n1049 ,n2112);
    nor g4653(n3025 ,n1048 ,n2220);
    nor g4654(n3024 ,n0[57] ,n1051);
    nor g4655(n3023 ,n1105 ,n1052);
    nor g4656(n3022 ,n1104 ,n1051);
    nor g4657(n3021 ,n1262 ,n1048);
    nor g4658(n3020 ,n1103 ,n2367);
    nor g4659(n3019 ,n1262 ,n2523);
    nor g4660(n3018 ,n1253 ,n2516);
    nor g4661(n3017 ,n1265 ,n2000);
    nor g4662(n3016 ,n1246 ,n1053);
    nor g4663(n3015 ,n1049 ,n2128);
    nor g4664(n3014 ,n1098 ,n1051);
    nor g4665(n3013 ,n1095 ,n2367);
    nor g4666(n3012 ,n1245 ,n2293);
    nor g4667(n3011 ,n1094 ,n2217);
    nor g4668(n3010 ,n1250 ,n2295);
    nor g4669(n3009 ,n1252 ,n2294);
    nor g4670(n3008 ,n1251 ,n2221);
    nor g4671(n3007 ,n1101 ,n2219);
    nor g4672(n3006 ,n1097 ,n2224);
    nor g4673(n3005 ,n1049 ,n2482);
    nor g4674(n3004 ,n1049 ,n2473);
    nor g4675(n3003 ,n1048 ,n2131);
    nor g4676(n3002 ,n0[59] ,n1051);
    nor g4677(n3001 ,n0[60] ,n1049);
    nor g4678(n3000 ,n1049 ,n2435);
    nor g4679(n2999 ,n2367 ,n2467);
    nor g4680(n2998 ,n1048 ,n2472);
    nor g4681(n2997 ,n1086 ,n2512);
    nor g4682(n2996 ,n1087 ,n2510);
    nor g4683(n2995 ,n1091 ,n2282);
    nor g4684(n2994 ,n0[63] ,n1048);
    nor g4685(n2993 ,n1048 ,n2133);
    nor g4686(n2992 ,n2367 ,n2110);
    nor g4687(n2991 ,n1236 ,n1052);
    nor g4688(n2990 ,n2367 ,n2416);
    nor g4689(n2989 ,n1072 ,n1051);
    nor g4690(n2988 ,n1239 ,n1049);
    nor g4691(n2987 ,n1235 ,n2257);
    nor g4692(n2986 ,n1081 ,n2230);
    nor g4693(n2985 ,n1238 ,n2259);
    nor g4694(n2984 ,n1236 ,n2514);
    nor g4695(n2983 ,n1074 ,n2261);
    nor g4696(n2982 ,n1233 ,n2215);
    nor g4697(n2981 ,n1080 ,n2254);
    nor g4698(n2980 ,n1232 ,n2260);
    nor g4699(n2979 ,n1077 ,n2228);
    nor g4700(n2978 ,n1070 ,n2223);
    nor g4701(n2977 ,n1072 ,n2292);
    nor g4702(n2976 ,n1228 ,n1052);
    nor g4703(n2975 ,n1228 ,n2218);
    nor g4704(n2974 ,n1048 ,n2470);
    nor g4705(n2973 ,n1064 ,n2226);
    nor g4706(n2972 ,n1226 ,n2262);
    nor g4707(n2971 ,n1226 ,n2237);
    nor g4708(n2970 ,n1056 ,n2061);
    nor g4709(n2969 ,n1054 ,n2044);
    nor g4710(n2968 ,n1053 ,n2028);
    nor g4711(n2967 ,n1054 ,n2050);
    nor g4712(n2966 ,n1053 ,n2024);
    nor g4713(n2965 ,n1053 ,n2052);
    nor g4714(n2964 ,n1054 ,n2092);
    nor g4715(n2963 ,n1052 ,n2054);
    nor g4716(n2962 ,n1054 ,n2036);
    nor g4717(n2961 ,n1056 ,n2076);
    nor g4718(n2960 ,n1053 ,n2006);
    nor g4719(n2959 ,n1056 ,n2020);
    nor g4720(n2958 ,n1056 ,n2022);
    nor g4721(n2957 ,n1054 ,n2047);
    nor g4722(n2956 ,n1056 ,n2018);
    nor g4723(n2955 ,n1052 ,n2058);
    nor g4724(n2954 ,n1056 ,n2041);
    nor g4725(n2953 ,n1056 ,n2008);
    nor g4726(n2952 ,n1056 ,n2010);
    nor g4727(n2951 ,n1054 ,n2012);
    nor g4728(n2950 ,n1056 ,n2081);
    nor g4729(n2949 ,n1054 ,n2014);
    nor g4730(n2948 ,n1052 ,n2038);
    nor g4731(n2947 ,n1056 ,n2017);
    nor g4732(n2946 ,n1056 ,n2026);
    nor g4733(n2945 ,n1052 ,n2004);
    nor g4734(n2944 ,n1056 ,n2056);
    nor g4735(n2943 ,n1056 ,n2079);
    nor g4736(n2942 ,n1048 ,n2124);
    nor g4737(n2941 ,n1410 ,n2452);
    nor g4738(n2940 ,n1385 ,n2441);
    nor g4739(n2939 ,n1049 ,n2122);
    nor g4740(n2938 ,n1380 ,n2487);
    nor g4741(n2937 ,n1544 ,n2216);
    nor g4742(n2936 ,n1421 ,n2465);
    nor g4743(n2935 ,n1441 ,n2449);
    nor g4744(n2934 ,n1049 ,n2101);
    nor g4745(n2933 ,n1390 ,n2445);
    nor g4746(n2932 ,n1408 ,n2443);
    nor g4747(n2931 ,n1450 ,n2458);
    nor g4748(n2930 ,n1462 ,n2450);
    nor g4749(n2929 ,n1393 ,n2462);
    nor g4750(n2928 ,n1420 ,n2447);
    nor g4751(n2927 ,n1443 ,n2460);
    nor g4752(n2926 ,n1404 ,n2456);
    nor g4753(n2925 ,n1386 ,n2454);
    nor g4754(n2924 ,n1382 ,n2464);
    nor g4755(n2923 ,n1049 ,n2097);
    nor g4756(n2922 ,n2510 ,n2465);
    nor g4757(n2921 ,n0[99] ,n2494);
    nor g4758(n2920 ,n0[115] ,n2504);
    nor g4759(n2919 ,n0[107] ,n2501);
    nor g4760(n2918 ,n1048 ,n2099);
    nor g4761(n2917 ,n2523 ,n2450);
    nor g4762(n2916 ,n0[11] ,n2519);
    nor g4763(n2915 ,n0[67] ,n2527);
    nor g4764(n2914 ,n0[35] ,n2525);
    nor g4765(n2913 ,n2367 ,n2480);
    nor g4766(n2912 ,n0[83] ,n2522);
    nor g4767(n2911 ,n2367 ,n2469);
    nor g4768(n2910 ,n1049 ,n2439);
    nor g4769(n2909 ,n2441 ,n2520);
    nor g4770(n2908 ,n1048 ,n2114);
    nor g4771(n2907 ,n0[43] ,n2489);
    nor g4772(n2906 ,n1048 ,n2073);
    nor g4773(n2905 ,n1049 ,n2378);
    nor g4774(n2904 ,n0[75] ,n2492);
    nor g4775(n2903 ,n2367 ,n2476);
    nor g4776(n2902 ,n1048 ,n2127);
    nor g4777(n2901 ,n1048 ,n2479);
    nor g4778(n2900 ,n1048 ,n2126);
    nor g4779(n2899 ,n1051 ,n2104);
    nor g4780(n2898 ,n2367 ,n2094);
    nor g4781(n2897 ,n1048 ,n2474);
    nor g4782(n2896 ,n1[55] ,n1999);
    nor g4783(n2895 ,n1064 ,n2263);
    nor g4784(n2894 ,n1048 ,n2125);
    nor g4785(n2893 ,n1049 ,n2211);
    nor g4786(n2892 ,n1049 ,n2436);
    nor g4787(n2891 ,n1064 ,n2258);
    nor g4788(n2890 ,n1064 ,n2291);
    nor g4789(n2889 ,n2367 ,n2132);
    nor g4790(n2888 ,n1051 ,n2212);
    nor g4791(n2887 ,n1054 ,n2000);
    nor g4792(n2886 ,n1052 ,n2075);
    nor g4793(n2885 ,n0[23] ,n1056);
    nor g4794(n2884 ,n1056 ,n2064);
    nor g4795(n2883 ,n1056 ,n2074);
    nor g4796(n2882 ,n1054 ,n2374);
    nor g4797(n2881 ,n2367 ,n2437);
    nor g4798(n2880 ,n1052 ,n2049);
    nor g4799(n2879 ,n1054 ,n2378);
    nor g4800(n2878 ,n1048 ,n2213);
    nor g4801(n2877 ,n1054 ,n2385);
    nor g4802(n2876 ,n1054 ,n2071);
    nor g4803(n2875 ,n1052 ,n2088);
    nor g4804(n2874 ,n1052 ,n2070);
    nor g4805(n2873 ,n1056 ,n2073);
    nor g4806(n2872 ,n1054 ,n2401);
    nor g4807(n2871 ,n1054 ,n2069);
    nor g4808(n2870 ,n1054 ,n2416);
    nor g4809(n2869 ,n1056 ,n2371);
    nor g4810(n2868 ,n1056 ,n2376);
    nor g4811(n2867 ,n1056 ,n2415);
    nor g4812(n2866 ,n1056 ,n2065);
    nor g4813(n2865 ,n1056 ,n2060);
    nor g4814(n2864 ,n1056 ,n2002);
    nor g4815(n2863 ,n1054 ,n2090);
    nor g4816(n2862 ,n1056 ,n2383);
    nor g4817(n2861 ,n1056 ,n2413);
    nor g4818(n2860 ,n1056 ,n2373);
    nor g4819(n2859 ,n1048 ,n2108);
    nor g4820(n2858 ,n1056 ,n2067);
    nor g4821(n2857 ,n1049 ,n2129);
    nor g4822(n2856 ,n1056 ,n2425);
    nor g4823(n2855 ,n1051 ,n2401);
    nor g4824(n2854 ,n2367 ,n2067);
    nor g4825(n2853 ,n1[85] ,n1051);
    or g4826(n2852 ,n0[85] ,n1051);
    nor g4827(n2851 ,n1051 ,n2477);
    nor g4828(n2850 ,n1054 ,n2085);
    nor g4829(n2849 ,n1[86] ,n1051);
    or g4830(n2848 ,n0[87] ,n1051);
    nor g4831(n2847 ,n1[87] ,n2367);
    nor g4832(n2846 ,n1053 ,n2227);
    nor g4833(n2845 ,n1049 ,n2109);
    nor g4834(n2844 ,n1053 ,n2068);
    nor g4835(n2843 ,n1051 ,n2136);
    nor g4836(n2842 ,n1053 ,n2072);
    nor g4837(n2841 ,n1054 ,n2063);
    or g4838(n2840 ,n1053 ,n2016);
    nor g4839(n2839 ,n1053 ,n2375);
    nor g4840(n3150 ,n0[15] ,n1052);
    nor g4841(n3149 ,n1[36] ,n1052);
    nor g4842(n3147 ,n0[3] ,n1056);
    nor g4843(n3145 ,n0[6] ,n1056);
    nor g4844(n3143 ,n0[30] ,n1054);
    nor g4845(n3141 ,n0[5] ,n1053);
    nor g4846(n3139 ,n0[7] ,n1053);
    nor g4847(n3138 ,n1[56] ,n1053);
    nor g4848(n3136 ,n0[8] ,n1052);
    nor g4849(n3134 ,n0[11] ,n1053);
    nor g4850(n3132 ,n0[17] ,n1056);
    nor g4851(n3130 ,n0[0] ,n1053);
    nor g4852(n3128 ,n0[20] ,n1052);
    nor g4853(n3126 ,n0[9] ,n1052);
    nor g4854(n3125 ,n1[42] ,n1052);
    nor g4855(n3123 ,n0[13] ,n1052);
    nor g4856(n3121 ,n0[22] ,n1052);
    nor g4857(n3119 ,n0[16] ,n1054);
    nor g4858(n3117 ,n0[19] ,n1052);
    nor g4859(n3115 ,n0[21] ,n1056);
    nor g4860(n3113 ,n0[25] ,n1052);
    nor g4861(n3111 ,n0[26] ,n1056);
    nor g4862(n3109 ,n0[27] ,n1052);
    nor g4863(n3107 ,n0[28] ,n1052);
    nor g4864(n3105 ,n0[29] ,n1056);
    nor g4865(n3103 ,n0[2] ,n1052);
    nor g4866(n3101 ,n0[31] ,n1053);
    nor g4867(n3099 ,n0[1] ,n1052);
    nor g4868(n3097 ,n0[12] ,n1054);
    nor g4869(n3095 ,n0[18] ,n1056);
    or g4870(n3094 ,n1020 ,n2248);
    or g4871(n3093 ,n1020 ,n2242);
    or g4872(n3092 ,n1020 ,n2246);
    nor g4873(n2838 ,n2447 ,n2359);
    nor g4874(n3090 ,n1145 ,n1053);
    nor g4875(n3089 ,n0[91] ,n2506);
    nor g4876(n2837 ,n2454 ,n2355);
    nor g4877(n2836 ,n2445 ,n2354);
    nor g4878(n2835 ,n2465 ,n2247);
    nor g4879(n2834 ,n2462 ,n2352);
    nor g4880(n2833 ,n2456 ,n2361);
    nor g4881(n2832 ,n2460 ,n2362);
    nor g4882(n2831 ,n2450 ,n2249);
    nor g4883(n2830 ,n2487 ,n2353);
    nor g4884(n2829 ,n2443 ,n2358);
    nor g4885(n2828 ,n2452 ,n2356);
    nor g4886(n3088 ,n0[59] ,n2499);
    nor g4887(n3087 ,n0[27] ,n2508);
    nor g4888(n2827 ,n2458 ,n2363);
    nor g4889(n2826 ,n2464 ,n2357);
    nor g4890(n2825 ,n2449 ,n2360);
    nor g4891(n3086 ,n1227 ,n1053);
    nor g4892(n3085 ,n1237 ,n1054);
    nor g4893(n3084 ,n1080 ,n1053);
    nor g4894(n3082 ,n1075 ,n1052);
    nor g4895(n3081 ,n1076 ,n1053);
    nor g4896(n3080 ,n1088 ,n1053);
    nor g4897(n3079 ,n1243 ,n1053);
    nor g4898(n3078 ,n1089 ,n1052);
    nor g4899(n3077 ,n1084 ,n1054);
    nor g4900(n3076 ,n1092 ,n1054);
    nor g4901(n3075 ,n1087 ,n1056);
    nor g4902(n3074 ,n1091 ,n1054);
    nor g4903(n3073 ,n1242 ,n1056);
    nor g4904(n3072 ,n1249 ,n1054);
    nor g4905(n3070 ,n1102 ,n1052);
    nor g4906(n3069 ,n1282 ,n1053);
    nor g4907(n3068 ,n1121 ,n1056);
    nor g4908(n3066 ,n1274 ,n1056);
    nor g4909(n3065 ,n1112 ,n1053);
    nor g4910(n3064 ,n1115 ,n1052);
    nor g4911(n3063 ,n1284 ,n1052);
    nor g4912(n3062 ,n1108 ,n1054);
    nor g4913(n3061 ,n1276 ,n1052);
    nor g4914(n3060 ,n1281 ,n1056);
    nor g4915(n3059 ,n1117 ,n1054);
    nor g4916(n3058 ,n1109 ,n1054);
    nor g4917(n3057 ,n1123 ,n1054);
    nor g4918(n3056 ,n1271 ,n1054);
    nor g4919(n3055 ,n1124 ,n1054);
    nor g4920(n3053 ,n1139 ,n1052);
    or g4921(n3052 ,n1356 ,n2368);
    or g4922(n1060 ,n3[0] ,n2229);
    nor g4923(n2824 ,n0[40] ,n1051);
    nor g4924(n2823 ,n1051 ,n2485);
    nor g4925(n2822 ,n0[55] ,n1048);
    nor g4926(n2821 ,n1051 ,n2065);
    nor g4927(n2820 ,n1051 ,n2111);
    nor g4928(n2819 ,n1051 ,n2134);
    nor g4929(n2818 ,n0[53] ,n1049);
    nor g4930(n2817 ,n1049 ,n2000);
    nor g4931(n2816 ,n1048 ,n2106);
    nor g4932(n2815 ,n1051 ,n2468);
    nor g4933(n2814 ,n1048 ,n2096);
    nor g4934(n2813 ,n1048 ,n2483);
    nor g4935(n2812 ,n1051 ,n2471);
    nor g4936(n2811 ,n1051 ,n2484);
    nor g4937(n2810 ,n2367 ,n2063);
    nor g4938(n2809 ,n2367 ,n2072);
    nor g4939(n2808 ,n2367 ,n2375);
    nor g4940(n2807 ,n1048 ,n2120);
    nor g4941(n2806 ,n2367 ,n2098);
    nor g4942(n2805 ,n1049 ,n2222);
    nor g4943(n2804 ,n1049 ,n2075);
    nor g4944(n2803 ,n2367 ,n2115);
    nor g4945(n2802 ,n2367 ,n2064);
    nor g4946(n2801 ,n1051 ,n2074);
    nor g4947(n2800 ,n0[62] ,n1049);
    nor g4948(n2799 ,n1051 ,n2376);
    nor g4949(n2798 ,n1051 ,n2116);
    nor g4950(n2797 ,n1051 ,n2049);
    nor g4951(n2796 ,n1051 ,n2123);
    nor g4952(n2795 ,n1049 ,n2117);
    nor g4953(n2794 ,n1048 ,n2385);
    nor g4954(n2793 ,n2367 ,n2071);
    nor g4955(n2792 ,n1[119] ,n1048);
    or g4956(n2791 ,n0[116] ,n1051);
    nor g4957(n2790 ,n1051 ,n2088);
    nor g4958(n2789 ,n2367 ,n2070);
    nor g4959(n2788 ,n1051 ,n2478);
    nor g4960(n2787 ,n2367 ,n2069);
    nor g4961(n2786 ,n2367 ,n2119);
    nor g4962(n2785 ,n2367 ,n2113);
    nor g4963(n2784 ,n1048 ,n2118);
    nor g4964(n2783 ,n1049 ,n2130);
    nor g4965(n2782 ,n1048 ,n2415);
    nor g4966(n2781 ,n0[61] ,n1048);
    nor g4967(n2780 ,n0[35] ,n1051);
    or g4968(n2779 ,n0[86] ,n1051);
    nor g4969(n2778 ,n1049 ,n2060);
    nor g4970(n2777 ,n2367 ,n2105);
    nor g4971(n2776 ,n1051 ,n2425);
    nor g4972(n2775 ,n2367 ,n2135);
    nor g4973(n2774 ,n2367 ,n2090);
    nor g4974(n2773 ,n2367 ,n2383);
    nor g4975(n2772 ,n1[43] ,n1049);
    nor g4976(n2771 ,n1049 ,n2413);
    nor g4977(n2770 ,n1051 ,n2068);
    nor g4978(n2769 ,n0[43] ,n1051);
    nor g4979(n2768 ,n1048 ,n2438);
    nor g4980(n2767 ,n2367 ,n2085);
    nor g4981(n2766 ,n0[52] ,n1049);
    nor g4982(n2765 ,n1051 ,n2121);
    nor g4983(n2764 ,n0[48] ,n2367);
    nor g4984(n2763 ,n1051 ,n2107);
    nor g4985(n2762 ,n1[116] ,n1051);
    nor g4986(n2761 ,n1044 ,n1929);
    nor g4987(n2760 ,n1044 ,n1966);
    nor g4988(n2759 ,n1042 ,n1945);
    or g4989(n2758 ,n1400 ,n1039);
    nor g4990(n2757 ,n1042 ,n1939);
    or g4991(n2756 ,n1498 ,n1039);
    nor g4992(n2755 ,n1044 ,n1986);
    or g4993(n2754 ,n1360 ,n1039);
    nor g4994(n2753 ,n1040 ,n1886);
    nor g4995(n2752 ,n1040 ,n1924);
    nor g4996(n2751 ,n1040 ,n1917);
    nor g4997(n2750 ,n1042 ,n1887);
    nor g4998(n2749 ,n1044 ,n1923);
    nor g4999(n2748 ,n1044 ,n1880);
    nor g5000(n2747 ,n1044 ,n1998);
    nor g5001(n2746 ,n1041 ,n1889);
    nor g5002(n2745 ,n1041 ,n1905);
    nor g5003(n2744 ,n1044 ,n1884);
    nor g5004(n2743 ,n1044 ,n1888);
    nor g5005(n2742 ,n1041 ,n1927);
    nor g5006(n2741 ,n1042 ,n1890);
    nor g5007(n2740 ,n1041 ,n1891);
    nor g5008(n2739 ,n1044 ,n1883);
    nor g5009(n2738 ,n1042 ,n1892);
    nor g5010(n2737 ,n1039 ,n1978);
    nor g5011(n2736 ,n1040 ,n1976);
    nor g5012(n2735 ,n1042 ,n1882);
    nor g5013(n2734 ,n1040 ,n1935);
    nor g5014(n2733 ,n1040 ,n1946);
    nor g5015(n2732 ,n1044 ,n1961);
    nor g5016(n2731 ,n1039 ,n1906);
    nor g5017(n2730 ,n1041 ,n1902);
    nor g5018(n2729 ,n1041 ,n1926);
    nor g5019(n2728 ,n1044 ,n1893);
    nor g5020(n2727 ,n1044 ,n1931);
    nor g5021(n2726 ,n1041 ,n1894);
    nor g5022(n2725 ,n1039 ,n1933);
    nor g5023(n2724 ,n1040 ,n1895);
    nor g5024(n2723 ,n1042 ,n1934);
    nor g5025(n2722 ,n1039 ,n1911);
    nor g5026(n2721 ,n1042 ,n1896);
    nor g5027(n2720 ,n1041 ,n1936);
    nor g5028(n2719 ,n1041 ,n1897);
    nor g5029(n2718 ,n1044 ,n1899);
    nor g5030(n2717 ,n1044 ,n1983);
    nor g5031(n2716 ,n1044 ,n1908);
    nor g5032(n2715 ,n1044 ,n1940);
    nor g5033(n2714 ,n1042 ,n1901);
    nor g5034(n2713 ,n1040 ,n1977);
    nor g5035(n2712 ,n1042 ,n1941);
    nor g5036(n2711 ,n1044 ,n1963);
    nor g5037(n2710 ,n1042 ,n1942);
    nor g5038(n2709 ,n1044 ,n1993);
    nor g5039(n2708 ,n1040 ,n1992);
    nor g5040(n2707 ,n1041 ,n1947);
    or g5041(n2706 ,n1478 ,n1039);
    nor g5042(n2705 ,n1044 ,n1970);
    nor g5043(n2704 ,n1041 ,n1957);
    nor g5044(n2703 ,n1040 ,n1885);
    nor g5045(n2702 ,n1044 ,n1909);
    nor g5046(n2701 ,n1039 ,n1910);
    nor g5047(n2700 ,n1042 ,n1904);
    nor g5048(n2699 ,n1044 ,n1964);
    nor g5049(n2698 ,n1044 ,n1994);
    nor g5050(n2697 ,n1039 ,n1881);
    or g5051(n2696 ,n1401 ,n1039);
    nor g5052(n2695 ,n1039 ,n1919);
    or g5053(n2694 ,n1434 ,n1039);
    nor g5054(n2693 ,n1039 ,n1953);
    nor g5055(n2692 ,n1040 ,n1954);
    nor g5056(n2691 ,n1040 ,n1900);
    or g5057(n2690 ,n1381 ,n1039);
    nor g5058(n2689 ,n1042 ,n1921);
    nor g5059(n2688 ,n1042 ,n1944);
    nor g5060(n2687 ,n1041 ,n1958);
    nor g5061(n2686 ,n1041 ,n1988);
    nor g5062(n2685 ,n1040 ,n1974);
    nor g5063(n2684 ,n1041 ,n1920);
    nor g5064(n2683 ,n1040 ,n1960);
    nor g5065(n2682 ,n1044 ,n1952);
    nor g5066(n2681 ,n1044 ,n1914);
    nor g5067(n2680 ,n1041 ,n1956);
    nor g5068(n2679 ,n1044 ,n1962);
    nor g5069(n2678 ,n1040 ,n1922);
    or g5070(n2677 ,n1365 ,n1042);
    nor g5071(n2676 ,n1041 ,n1943);
    nor g5072(n2675 ,n1041 ,n1975);
    nor g5073(n2674 ,n1044 ,n1948);
    nor g5074(n2673 ,n1040 ,n1965);
    nor g5075(n2672 ,n1044 ,n1990);
    nor g5076(n2671 ,n1044 ,n1912);
    nor g5077(n2670 ,n1041 ,n1968);
    nor g5078(n2669 ,n1040 ,n1997);
    nor g5079(n2668 ,n1040 ,n1984);
    nor g5080(n2667 ,n1044 ,n1898);
    nor g5081(n2666 ,n1041 ,n1938);
    nor g5082(n2665 ,n1042 ,n1972);
    nor g5083(n2664 ,n1039 ,n1995);
    nor g5084(n2663 ,n1042 ,n1913);
    nor g5085(n2662 ,n1044 ,n1951);
    nor g5086(n2661 ,n1042 ,n1928);
    or g5087(n2660 ,n1383 ,n1039);
    nor g5088(n2659 ,n1040 ,n1903);
    nor g5089(n2658 ,n1040 ,n1981);
    nor g5090(n2657 ,n1040 ,n1987);
    nor g5091(n2656 ,n1040 ,n1955);
    nor g5092(n2655 ,n1044 ,n1973);
    nor g5093(n2654 ,n1041 ,n1959);
    nor g5094(n2653 ,n1040 ,n1930);
    nor g5095(n2652 ,n1040 ,n1918);
    nor g5096(n2651 ,n1040 ,n1915);
    nor g5097(n2650 ,n1040 ,n1967);
    nor g5098(n2649 ,n1041 ,n1985);
    nor g5099(n2648 ,n1042 ,n1950);
    nor g5100(n2647 ,n1040 ,n1937);
    nor g5101(n2646 ,n1041 ,n1949);
    nor g5102(n2645 ,n1040 ,n1969);
    nor g5103(n2644 ,n1041 ,n1982);
    nor g5104(n2643 ,n1042 ,n1980);
    nor g5105(n2642 ,n1041 ,n1925);
    nor g5106(n2641 ,n1041 ,n1971);
    nor g5107(n2640 ,n1040 ,n1996);
    nor g5108(n2639 ,n1042 ,n1907);
    nor g5109(n2638 ,n1042 ,n1979);
    nor g5110(n2637 ,n1041 ,n1991);
    nor g5111(n2636 ,n1042 ,n1932);
    nor g5112(n2635 ,n1044 ,n1989);
    nor g5113(n2634 ,n1042 ,n1916);
    nor g5114(n2633 ,n0[72] ,n2240);
    nor g5115(n2632 ,n1026 ,n2395);
    nor g5116(n2631 ,n1026 ,n2419);
    nor g5117(n2630 ,n1026 ,n2390);
    nor g5118(n2629 ,n1028 ,n2417);
    nor g5119(n2628 ,n1027 ,n2391);
    nor g5120(n2627 ,n1030 ,n2420);
    nor g5121(n2626 ,n1026 ,n2418);
    nor g5122(n2625 ,n1514 ,n2339);
    nor g5123(n2624 ,n0[8] ,n2231);
    nor g5124(n2623 ,n1026 ,n2414);
    or g5125(n2622 ,n1684 ,n2300);
    nor g5126(n2621 ,n1026 ,n2409);
    nor g5127(n2620 ,n0[80] ,n2235);
    nor g5128(n2619 ,n1030 ,n2405);
    or g5129(n2618 ,n1618 ,n2313);
    nor g5130(n2617 ,n1030 ,n2434);
    nor g5131(n2616 ,n1027 ,n2380);
    nor g5132(n2615 ,n1027 ,n2406);
    nor g5133(n2614 ,n1028 ,n2412);
    nor g5134(n2613 ,n1028 ,n2392);
    nor g5135(n2612 ,n1027 ,n2431);
    nor g5136(n2611 ,n1027 ,n2398);
    nor g5137(n2610 ,n1028 ,n2511);
    nor g5138(n2609 ,n1027 ,n2429);
    nor g5139(n2608 ,n1030 ,n2388);
    nor g5140(n2607 ,n1030 ,n2424);
    nor g5141(n2606 ,n1026 ,n2394);
    nor g5142(n2605 ,n1027 ,n2407);
    or g5143(n2604 ,n1623 ,n2301);
    nor g5144(n2603 ,n1028 ,n2393);
    nor g5145(n2602 ,n1028 ,n2421);
    nor g5146(n2601 ,n1030 ,n2509);
    nor g5147(n2600 ,n1026 ,n2423);
    nor g5148(n2599 ,n1030 ,n2426);
    nor g5149(n2598 ,n1030 ,n2430);
    nor g5150(n2597 ,n1027 ,n2427);
    nor g5151(n2596 ,n1026 ,n2433);
    or g5152(n2595 ,n1673 ,n2346);
    nor g5153(n2594 ,n1030 ,n2490);
    nor g5154(n2593 ,n1026 ,n2387);
    nor g5155(n2592 ,n1028 ,n2396);
    or g5156(n2591 ,n1692 ,n2314);
    nor g5157(n2590 ,n1027 ,n2400);
    or g5158(n2589 ,n1627 ,n2302);
    or g5159(n2588 ,n1681 ,n2312);
    or g5160(n2587 ,n1543 ,n2497);
    nor g5161(n2586 ,n1026 ,n2382);
    or g5162(n2585 ,n1713 ,n2321);
    nor g5163(n2584 ,n1027 ,n2428);
    or g5164(n2583 ,n1705 ,n2307);
    nor g5165(n2582 ,n1030 ,n2399);
    or g5166(n2581 ,n1645 ,n2344);
    or g5167(n2580 ,n1668 ,n2308);
    or g5168(n2579 ,n1683 ,n2350);
    nor g5169(n2578 ,n0[123] ,n2497);
    or g5170(n2577 ,n1664 ,n2323);
    nor g5171(n2576 ,n1030 ,n2377);
    nor g5172(n2575 ,n1027 ,n2404);
    nor g5173(n2574 ,n1027 ,n2397);
    or g5174(n2573 ,n1662 ,n2349);
    or g5175(n2572 ,n1659 ,n2348);
    nor g5176(n2571 ,n0[64] ,n2236);
    nor g5177(n2570 ,n1027 ,n2502);
    nor g5178(n2569 ,n1028 ,n2389);
    nor g5179(n2568 ,n1026 ,n2403);
    or g5180(n2567 ,n1676 ,n2310);
    or g5181(n2566 ,n1657 ,n2267);
    nor g5182(n2565 ,n0[112] ,n2239);
    or g5183(n2564 ,n1642 ,n2343);
    nor g5184(n2563 ,n1030 ,n2381);
    nor g5185(n2562 ,n0[104] ,n2232);
    or g5186(n2561 ,n1628 ,n2347);
    or g5187(n2560 ,n1625 ,n2345);
    or g5188(n2559 ,n1712 ,n2264);
    nor g5189(n2558 ,n1028 ,n2496);
    nor g5190(n2557 ,n1026 ,n2379);
    or g5191(n2556 ,n1654 ,n2311);
    or g5192(n2555 ,n1698 ,n2316);
    or g5193(n2554 ,n1634 ,n2351);
    nor g5194(n2553 ,n1028 ,n2384);
    nor g5195(n2552 ,n1026 ,n2408);
    nor g5196(n2551 ,n0[96] ,n2233);
    nor g5197(n2550 ,n0[32] ,n2234);
    nor g5198(n2549 ,n1030 ,n2411);
    nor g5199(n2548 ,n1027 ,n2432);
    nor g5200(n2547 ,n1030 ,n2495);
    or g5201(n2546 ,n1679 ,n2268);
    nor g5202(n2545 ,n0[40] ,n2238);
    or g5203(n2544 ,n1648 ,n2255);
    or g5204(n2543 ,n1646 ,n2309);
    nor g5205(n2542 ,n0[91] ,n2505);
    nor g5206(n2541 ,n0[51] ,n2253);
    nor g5207(n2540 ,n0[3] ,n2252);
    nor g5208(n2539 ,n0[11] ,n2518);
    nor g5209(n2538 ,n0[19] ,n2251);
    nor g5210(n2537 ,n0[27] ,n2507);
    nor g5211(n2536 ,n0[107] ,n2500);
    nor g5212(n2535 ,n0[115] ,n2503);
    nor g5213(n2534 ,n0[99] ,n2493);
    nor g5214(n2533 ,n0[75] ,n2491);
    nor g5215(n2532 ,n0[35] ,n2524);
    nor g5216(n2531 ,n0[43] ,n2488);
    nor g5217(n2530 ,n0[67] ,n2526);
    nor g5218(n2529 ,n0[59] ,n2498);
    nor g5219(n2528 ,n0[83] ,n2521);
    not g5220(n2527 ,n2526);
    not g5221(n2525 ,n2524);
    not g5222(n2522 ,n2521);
    not g5223(n2519 ,n2518);
    not g5224(n2517 ,n2516);
    not g5225(n2515 ,n2514);
    not g5226(n2513 ,n2512);
    not g5227(n2508 ,n2507);
    not g5228(n2506 ,n2505);
    not g5229(n2504 ,n2503);
    not g5230(n2501 ,n2500);
    not g5231(n2499 ,n2498);
    not g5232(n2494 ,n2493);
    not g5233(n2492 ,n2491);
    not g5234(n2489 ,n2488);
    not g5235(n2487 ,n2486);
    not g5236(n2464 ,n2463);
    not g5237(n2462 ,n2461);
    not g5238(n2460 ,n2459);
    not g5239(n2458 ,n2457);
    not g5240(n2456 ,n2455);
    not g5241(n2454 ,n2453);
    not g5242(n2452 ,n2451);
    not g5243(n2449 ,n2448);
    not g5244(n2447 ,n2446);
    not g5245(n2445 ,n2444);
    not g5246(n2443 ,n2442);
    not g5247(n2441 ,n2440);
    not g5248(n2373 ,n2372);
    not g5249(n2371 ,n2370);
    not g5250(n2369 ,n2368);
    not g5251(n1054 ,n1055);
    not g5252(n1053 ,n1055);
    not g5253(n1052 ,n1055);
    not g5254(n1055 ,n1056);
    not g5255(n1049 ,n1050);
    not g5256(n1048 ,n1050);
    not g5257(n2367 ,n1050);
    not g5258(n1050 ,n1051);
    not g5259(n2366 ,n1047);
    not g5260(n2365 ,n1047);
    not g5261(n1045 ,n1047);
    not g5262(n1047 ,n1046);
    not g5263(n1042 ,n1043);
    not g5264(n1039 ,n1043);
    not g5265(n1040 ,n1043);
    not g5266(n1041 ,n1043);
    not g5267(n1043 ,n1044);
    not g5268(n2364 ,n1037);
    not g5269(n1034 ,n1037);
    not g5270(n1035 ,n1037);
    not g5271(n1036 ,n1037);
    not g5272(n1037 ,n1038);
    nor g5273(n2363 ,n1253 ,n1448);
    nor g5274(n2362 ,n1097 ,n1526);
    nor g5275(n2361 ,n1101 ,n1520);
    nor g5276(n2360 ,n1251 ,n1522);
    nor g5277(n2359 ,n1094 ,n1529);
    nor g5278(n2358 ,n1086 ,n1413);
    nor g5279(n2357 ,n1081 ,n1539);
    nor g5280(n2356 ,n1236 ,n1426);
    nor g5281(n2355 ,n1070 ,n1553);
    nor g5282(n2354 ,n1077 ,n1531);
    nor g5283(n2353 ,n1233 ,n1542);
    nor g5284(n2352 ,n1228 ,n1535);
    nor g5285(n2351 ,n1152 ,n1730);
    nor g5286(n2350 ,n1303 ,n1032);
    nor g5287(n2349 ,n1305 ,n1032);
    nor g5288(n2348 ,n1153 ,n1032);
    nor g5289(n2347 ,n1151 ,n1032);
    nor g5290(n2346 ,n1149 ,n1032);
    nor g5291(n2345 ,n1147 ,n1730);
    nor g5292(n2344 ,n1302 ,n1729);
    nor g5293(n2343 ,n1306 ,n1729);
    nor g5294(n2342 ,n1301 ,n1032);
    nor g5295(n2341 ,n1148 ,n1032);
    nor g5296(n2340 ,n1304 ,n1032);
    nor g5297(n2339 ,n1227 ,n1743);
    nor g5298(n2338 ,n1113 ,n1032);
    nor g5299(n2337 ,n1277 ,n1032);
    nor g5300(n2336 ,n1275 ,n1032);
    nor g5301(n2335 ,n1283 ,n1730);
    nor g5302(n2334 ,n1279 ,n1032);
    nor g5303(n2333 ,n1272 ,n1032);
    nor g5304(n2332 ,n1111 ,n1032);
    nor g5305(n2331 ,n1269 ,n1032);
    nor g5306(n2330 ,n1120 ,n1032);
    nor g5307(n2329 ,n1273 ,n1730);
    nor g5308(n2328 ,n1107 ,n1032);
    nor g5309(n2327 ,n1278 ,n1032);
    nor g5310(n2326 ,n1110 ,n1032);
    nor g5311(n2325 ,n1280 ,n1730);
    nor g5312(n2324 ,n1119 ,n1032);
    nor g5313(n2323 ,n1112 ,n11);
    nor g5314(n2322 ,n1116 ,n1032);
    nor g5315(n2321 ,n1266 ,n1032);
    nor g5316(n2320 ,n1118 ,n1730);
    nor g5317(n2319 ,n1114 ,n1730);
    nor g5318(n2318 ,n1268 ,n1730);
    nor g5319(n2317 ,n1256 ,n1032);
    nor g5320(n2316 ,n1255 ,n1032);
    nor g5321(n2315 ,n1105 ,n1032);
    nor g5322(n2314 ,n1104 ,n1730);
    nor g5323(n2313 ,n1260 ,n11);
    nor g5324(n2312 ,n1253 ,n1032);
    nor g5325(n2311 ,n1262 ,n1032);
    nor g5326(n2310 ,n1264 ,n1032);
    nor g5327(n2309 ,n1103 ,n1730);
    nor g5328(n2308 ,n1094 ,n1729);
    nor g5329(n2307 ,n1095 ,n1032);
    nor g5330(n2306 ,n1245 ,n1032);
    nor g5331(n2305 ,n1099 ,n1730);
    nor g5332(n2304 ,n1097 ,n11);
    nor g5333(n2303 ,n1250 ,n1032);
    nor g5334(n2302 ,n1098 ,n1032);
    nor g5335(n2301 ,n1252 ,n1730);
    nor g5336(n2300 ,n1101 ,n1032);
    nor g5337(n2299 ,n1100 ,n1032);
    nor g5338(n2298 ,n1247 ,n11);
    nor g5339(n2297 ,n1248 ,n1730);
    nor g5340(n2296 ,n1251 ,n1730);
    nor g5341(n2295 ,n1097 ,n1549);
    nor g5342(n2294 ,n1101 ,n1536);
    nor g5343(n2293 ,n1251 ,n1524);
    nor g5344(n2292 ,n1094 ,n1550);
    nor g5345(n2291 ,n1098 ,n1615);
    nor g5346(n2290 ,n1093 ,n1032);
    nor g5347(n2289 ,n1240 ,n1032);
    nor g5348(n2288 ,n1083 ,n1730);
    nor g5349(n2287 ,n1086 ,n1730);
    nor g5350(n2286 ,n1244 ,n11);
    nor g5351(n2285 ,n1085 ,n1032);
    nor g5352(n2284 ,n1090 ,n1032);
    nor g5353(n2283 ,n1241 ,n1730);
    nor g5354(n2282 ,n1092 ,n1544);
    nor g5355(n2281 ,n1231 ,n1729);
    nor g5356(n2280 ,n1070 ,n1729);
    nor g5357(n2279 ,n1233 ,n11);
    nor g5358(n2278 ,n1078 ,n1032);
    nor g5359(n2277 ,n1238 ,n1032);
    nor g5360(n2276 ,n1074 ,n11);
    nor g5361(n2275 ,n1232 ,n1730);
    nor g5362(n2274 ,n1234 ,n1032);
    nor g5363(n2273 ,n1235 ,n1730);
    nor g5364(n2272 ,n1079 ,n1032);
    nor g5365(n2271 ,n1230 ,n1730);
    nor g5366(n2270 ,n1073 ,n1729);
    nor g5367(n2269 ,n1071 ,n1032);
    nor g5368(n2268 ,n1236 ,n1032);
    nor g5369(n2267 ,n1072 ,n1032);
    nor g5370(n2266 ,n1081 ,n1032);
    nor g5371(n2265 ,n1077 ,n1032);
    nor g5372(n2264 ,n1239 ,n1032);
    nor g5373(n2263 ,n1071 ,n1609);
    nor g5374(n2262 ,n1231 ,n1363);
    nor g5375(n2261 ,n1233 ,n1540);
    nor g5376(n2260 ,n1077 ,n1532);
    nor g5377(n2259 ,n1070 ,n1551);
    nor g5378(n2258 ,n1076 ,n1608);
    nor g5379(n2257 ,n1081 ,n1537);
    nor g5380(n2256 ,n1229 ,n1730);
    nor g5381(n2255 ,n1228 ,n1729);
    nor g5382(n2254 ,n1228 ,n1533);
    nor g5383(n2253 ,n1064 ,n1516);
    nor g5384(n2252 ,n1064 ,n1527);
    nor g5385(n2251 ,n1020 ,n1523);
    nor g5386(n2250 ,n1226 ,n1729);
    nor g5387(n2249 ,n0[49] ,n1745);
    nor g5388(n2248 ,n0[19] ,n1523);
    nor g5389(n2247 ,n0[1] ,n1742);
    nor g5390(n2246 ,n0[3] ,n1527);
    nor g5391(n2245 ,n0[120] ,n1602);
    nor g5392(n2244 ,n0[0] ,n1738);
    nor g5393(n2243 ,n0[48] ,n1735);
    nor g5394(n2242 ,n0[51] ,n1516);
    nor g5395(n2241 ,n0[16] ,n1743);
    nor g5396(n2240 ,n1064 ,n1403);
    nor g5397(n2239 ,n1064 ,n1394);
    nor g5398(n2238 ,n1064 ,n1422);
    nor g5399(n2237 ,n1064 ,n1543);
    nor g5400(n2236 ,n1064 ,n1430);
    nor g5401(n2235 ,n1064 ,n1377);
    nor g5402(n2234 ,n1064 ,n1396);
    nor g5403(n2233 ,n1064 ,n1428);
    nor g5404(n2232 ,n1064 ,n1399);
    nor g5405(n2231 ,n1064 ,n1376);
    nor g5406(n2230 ,n1603 ,n1537);
    or g5407(n2229 ,n1351 ,n1513);
    nor g5408(n2228 ,n1601 ,n1532);
    xnor g5409(n2227 ,n0[14] ,n1[46]);
    or g5410(n2226 ,n1736 ,n1466);
    xnor g5411(n2225 ,n0[50] ,n1[50]);
    nor g5412(n2224 ,n1613 ,n1549);
    nor g5413(n2223 ,n1605 ,n1551);
    xnor g5414(n2222 ,n0[97] ,n1[97]);
    nor g5415(n2221 ,n1614 ,n1524);
    xnor g5416(n2220 ,n0[56] ,n1[56]);
    nor g5417(n2219 ,n1611 ,n1536);
    nor g5418(n2218 ,n1600 ,n1533);
    nor g5419(n2217 ,n1606 ,n1550);
    or g5420(n2216 ,n1736 ,n1514);
    nor g5421(n2215 ,n1604 ,n1540);
    xnor g5422(n2214 ,n0[120] ,n1[120]);
    xnor g5423(n2213 ,n0[83] ,n1[83]);
    xnor g5424(n2212 ,n0[82] ,n1[82]);
    xnor g5425(n2211 ,n0[80] ,n1[80]);
    xnor g5426(n2210 ,n0[20] ,n4[28]);
    xnor g5427(n2209 ,n0[28] ,n4[4]);
    xnor g5428(n2208 ,n0[29] ,n4[5]);
    xnor g5429(n2207 ,n0[30] ,n4[6]);
    xnor g5430(n2206 ,n0[31] ,n4[7]);
    xnor g5431(n2205 ,n0[108] ,n4[4]);
    nor g5432(n2526 ,n1064 ,n1367);
    xnor g5433(n2204 ,n0[116] ,n4[4]);
    nor g5434(n2524 ,n1064 ,n1436);
    nor g5435(n2523 ,n1095 ,n1734);
    nor g5436(n2521 ,n1064 ,n1366);
    nor g5437(n2520 ,n1226 ,n1402);
    xnor g5438(n2203 ,n0[68] ,n4[28]);
    nor g5439(n2518 ,n1064 ,n1357);
    xnor g5440(n2202 ,n0[70] ,n1[86]);
    xnor g5441(n2201 ,n0[18] ,n4[26]);
    xnor g5442(n2200 ,n0[71] ,n1[87]);
    nor g5443(n2516 ,n1260 ,n1375);
    xnor g5444(n2199 ,n0[110] ,n4[6]);
    nor g5445(n2514 ,n1084 ,n1397);
    xnor g5446(n2198 ,n0[122] ,n4[10]);
    xnor g5447(n2197 ,n0[123] ,n4[11]);
    xnor g5448(n2196 ,n0[0] ,n4[16]);
    nor g5449(n2512 ,n1244 ,n1384);
    xnor g5450(n2195 ,n0[89] ,n4[17]);
    xnor g5451(n2194 ,n0[11] ,n4[27]);
    xnor g5452(n2193 ,n0[121] ,n4[9]);
    xnor g5453(n2192 ,n0[88] ,n4[16]);
    xnor g5454(n2191 ,n0[76] ,n4[4]);
    xnor g5455(n2190 ,n0[118] ,n4[6]);
    xnor g5456(n2189 ,n0[78] ,n4[6]);
    xnor g5457(n2188 ,n0[77] ,n4[5]);
    xnor g5458(n2187 ,n0[117] ,n4[5]);
    nor g5459(n2186 ,n1518 ,n1515);
    xnor g5460(n2185 ,n0[33] ,n1[49]);
    xnor g5461(n2184 ,n0[97] ,n4[9]);
    xnor g5462(n2183 ,n0[41] ,n1[57]);
    xnor g5463(n2182 ,n0[58] ,n4[18]);
    xnor g5464(n2181 ,n0[65] ,n4[25]);
    xnor g5465(n2180 ,n0[79] ,n4[7]);
    xnor g5466(n2179 ,n0[16] ,n4[24]);
    xnor g5467(n2178 ,n0[120] ,n4[8]);
    nor g5468(n2511 ,n1447 ,n1546);
    nor g5469(n2177 ,n1740 ,n1517);
    xnor g5470(n2176 ,n0[119] ,n4[7]);
    nor g5471(n2510 ,n1237 ,n1737);
    xnor g5472(n2175 ,n0[32] ,n1[48]);
    xnor g5473(n2174 ,n0[42] ,n4[18]);
    xnor g5474(n2173 ,n0[64] ,n1[80]);
    xnor g5475(n2172 ,n0[66] ,n1[82]);
    nor g5476(n2509 ,n1445 ,n1517);
    xnor g5477(n2171 ,n0[67] ,n1[83]);
    xnor g5478(n2170 ,n0[39] ,n1[55]);
    nor g5479(n2507 ,n0[26] ,n1547);
    xnor g5480(n2169 ,n0[105] ,n4[1]);
    nor g5481(n2505 ,n0[90] ,n1545);
    xnor g5482(n2168 ,n0[113] ,n4[1]);
    xnor g5483(n2167 ,n0[109] ,n4[5]);
    xnor g5484(n2166 ,n0[9] ,n4[25]);
    xnor g5485(n2165 ,n0[17] ,n4[25]);
    xnor g5486(n2164 ,n0[43] ,n1[59]);
    xnor g5487(n2163 ,n0[73] ,n4[1]);
    xnor g5488(n2162 ,n0[26] ,n4[2]);
    nor g5489(n2503 ,n1064 ,n1369);
    xnor g5490(n2161 ,n0[90] ,n4[18]);
    nor g5491(n2502 ,n1739 ,n1439);
    nor g5492(n2500 ,n1064 ,n1359);
    xnor g5493(n2160 ,n0[119] ,n0[103]);
    nor g5494(n2498 ,n0[58] ,n1548);
    nor g5495(n2497 ,n0[121] ,n1364);
    nor g5496(n2496 ,n1740 ,n1432);
    nor g5497(n2495 ,n1518 ,n1494);
    xnor g5498(n2159 ,n0[75] ,n4[3]);
    nor g5499(n2493 ,n1064 ,n1358);
    xnor g5500(n2158 ,n0[111] ,n4[7]);
    nor g5501(n2491 ,n1064 ,n1362);
    xnor g5502(n2157 ,n0[115] ,n4[3]);
    xnor g5503(n2156 ,n0[25] ,n4[1]);
    nor g5504(n2155 ,n1739 ,n1546);
    xnor g5505(n2154 ,n0[112] ,n4[0]);
    xnor g5506(n2153 ,n0[107] ,n4[3]);
    xnor g5507(n2152 ,n0[114] ,n4[2]);
    xnor g5508(n2151 ,n0[35] ,n1[51]);
    xnor g5509(n2150 ,n0[106] ,n4[2]);
    nor g5510(n2490 ,n1559 ,n1515);
    xnor g5511(n2149 ,n0[74] ,n4[2]);
    nor g5512(n2488 ,n1064 ,n1472);
    xnor g5513(n2148 ,n0[106] ,n0[74]);
    xnor g5514(n2147 ,n0[40] ,n0[24]);
    xnor g5515(n2146 ,n0[35] ,n0[19]);
    xnor g5516(n2145 ,n0[43] ,n0[27]);
    xnor g5517(n2144 ,n0[97] ,n0[81]);
    xnor g5518(n2143 ,n0[40] ,n1[56]);
    xnor g5519(n2142 ,n0[69] ,n1[85]);
    xnor g5520(n2141 ,n0[34] ,n1[50]);
    xnor g5521(n2140 ,n0[72] ,n4[0]);
    xnor g5522(n2139 ,n1[43] ,n4[3]);
    xnor g5523(n2138 ,n0[84] ,n4[28]);
    xnor g5524(n2137 ,n0[12] ,n4[28]);
    nor g5525(n2486 ,n1064 ,n1405);
    xnor g5526(n2485 ,n0[34] ,n1[34]);
    xnor g5527(n2484 ,n0[32] ,n1[32]);
    xnor g5528(n2483 ,n0[33] ,n1[33]);
    xnor g5529(n2482 ,n0[58] ,n1[58]);
    xnor g5530(n2481 ,n0[41] ,n1[41]);
    xnor g5531(n2480 ,n0[121] ,n1[121]);
    xnor g5532(n2479 ,n0[115] ,n1[115]);
    xnor g5533(n2478 ,n0[122] ,n1[122]);
    xnor g5534(n2477 ,n0[114] ,n1[114]);
    xnor g5535(n2476 ,n0[75] ,n1[75]);
    xnor g5536(n2475 ,n0[105] ,n1[105]);
    xnor g5537(n2474 ,n0[112] ,n1[112]);
    xnor g5538(n2473 ,n0[106] ,n1[106]);
    xnor g5539(n2472 ,n0[123] ,n1[123]);
    xnor g5540(n2471 ,n0[74] ,n1[74]);
    xnor g5541(n2470 ,n0[89] ,n1[89]);
    xnor g5542(n2469 ,n0[72] ,n1[72]);
    xnor g5543(n2468 ,n0[104] ,n1[104]);
    xnor g5544(n2467 ,n0[107] ,n1[107]);
    xnor g5545(n2466 ,n0[42] ,n1[42]);
    or g5546(n2465 ,n1020 ,n1418);
    nor g5547(n2463 ,n1064 ,n1425);
    nor g5548(n2461 ,n1064 ,n1414);
    nor g5549(n2459 ,n1064 ,n1463);
    nor g5550(n2457 ,n1064 ,n1437);
    nor g5551(n2455 ,n1020 ,n1449);
    nor g5552(n2453 ,n1020 ,n1412);
    nor g5553(n2451 ,n1064 ,n1395);
    or g5554(n2450 ,n1020 ,n1454);
    nor g5555(n2448 ,n1064 ,n1423);
    nor g5556(n2446 ,n1064 ,n1453);
    nor g5557(n2444 ,n1064 ,n1409);
    nor g5558(n2442 ,n1064 ,n1398);
    nor g5559(n2440 ,n1064 ,n1374);
    xnor g5560(n2439 ,n0[73] ,n1[73]);
    xnor g5561(n2438 ,n0[90] ,n1[90]);
    xnor g5562(n2437 ,n0[113] ,n1[113]);
    xnor g5563(n2436 ,n0[81] ,n1[81]);
    xnor g5564(n2435 ,n0[88] ,n1[88]);
    nor g5565(n2434 ,n1599 ,n1497);
    nor g5566(n2433 ,n1587 ,n1475);
    nor g5567(n2432 ,n1506 ,n1491);
    nor g5568(n2431 ,n1558 ,n1582);
    nor g5569(n2430 ,n1715 ,n1485);
    nor g5570(n2429 ,n1446 ,n1573);
    nor g5571(n2428 ,n1596 ,n1487);
    nor g5572(n2427 ,n1507 ,n1492);
    nor g5573(n2426 ,n1588 ,n1469);
    xnor g5574(n2425 ,n0[3] ,n1[3]);
    nor g5575(n2424 ,n1595 ,n1480);
    nor g5576(n2423 ,n1557 ,n1575);
    xnor g5577(n2422 ,n0[80] ,n4[24]);
    nor g5578(n2421 ,n1597 ,n1468);
    nor g5579(n2420 ,n1563 ,n1489);
    nor g5580(n2419 ,n1612 ,n1568);
    nor g5581(n2418 ,n1594 ,n1474);
    nor g5582(n2417 ,n1512 ,n1583);
    xnor g5583(n2416 ,n0[11] ,n1[11]);
    xnor g5584(n2415 ,n0[8] ,n1[8]);
    nor g5585(n2414 ,n1727 ,n1490);
    xnor g5586(n2413 ,n0[0] ,n1[0]);
    nor g5587(n2412 ,n1502 ,n1500);
    nor g5588(n2411 ,n1511 ,n1499);
    xnor g5589(n2410 ,n0[83] ,n4[27]);
    nor g5590(n2409 ,n1610 ,n1471);
    nor g5591(n2408 ,n1617 ,n1493);
    nor g5592(n2407 ,n1590 ,n1488);
    nor g5593(n2406 ,n1725 ,n1574);
    nor g5594(n2405 ,n1607 ,n1496);
    nor g5595(n2404 ,n1504 ,n1473);
    nor g5596(n2403 ,n1505 ,n1577);
    xnor g5597(n2402 ,n0[82] ,n4[26]);
    xnor g5598(n2401 ,n0[25] ,n1[25]);
    nor g5599(n2400 ,n1571 ,n1495);
    nor g5600(n2399 ,n1570 ,n1481);
    nor g5601(n2398 ,n1591 ,n1482);
    nor g5602(n2397 ,n1503 ,n1457);
    nor g5603(n2396 ,n1589 ,n1483);
    nor g5604(n2395 ,n1510 ,n1584);
    nor g5605(n2394 ,n1562 ,n1476);
    nor g5606(n2393 ,n1508 ,n1501);
    nor g5607(n2392 ,n1572 ,n1484);
    nor g5608(n2391 ,n1554 ,n1567);
    nor g5609(n2390 ,n1561 ,n1564);
    nor g5610(n2389 ,n1593 ,n1470);
    nor g5611(n2388 ,n1616 ,n1477);
    nor g5612(n2387 ,n1556 ,n1580);
    xnor g5613(n2386 ,n0[116] ,n0[100]);
    xnor g5614(n2385 ,n0[16] ,n1[16]);
    nor g5615(n2384 ,n1635 ,n1581);
    xnor g5616(n2383 ,n0[1] ,n1[1]);
    nor g5617(n2382 ,n1592 ,n1467);
    nor g5618(n2381 ,n1586 ,n1440);
    nor g5619(n2380 ,n1555 ,n1579);
    nor g5620(n2379 ,n1509 ,n1576);
    xnor g5621(n2378 ,n0[17] ,n1[17]);
    nor g5622(n2377 ,n1560 ,n1578);
    xnor g5623(n2376 ,n0[9] ,n1[9]);
    xnor g5624(n2375 ,n0[27] ,n1[27]);
    xnor g5625(n2374 ,n0[19] ,n1[19]);
    xnor g5626(n2372 ,n1[24] ,n1236);
    xnor g5627(n2370 ,n1[10] ,n1228);
    nor g5628(n2368 ,n7663 ,n1732);
    or g5629(n1056 ,n7664 ,n1733);
    or g5630(n1051 ,n7665 ,n1638);
    or g5631(n1046 ,n1733 ,n1513);
    or g5632(n1044 ,n7665 ,n1732);
    or g5633(n1038 ,n1726 ,n1513);
    not g5634(n2093 ,n2092);
    not g5635(n2082 ,n2081);
    not g5636(n2080 ,n2079);
    not g5637(n2077 ,n2076);
    not g5638(n2062 ,n2061);
    not g5639(n2059 ,n2058);
    not g5640(n2057 ,n2056);
    not g5641(n2055 ,n2054);
    not g5642(n2053 ,n2052);
    not g5643(n2051 ,n2050);
    not g5644(n2048 ,n2047);
    not g5645(n2045 ,n2044);
    not g5646(n2042 ,n2041);
    not g5647(n2039 ,n2038);
    not g5648(n2037 ,n2036);
    not g5649(n2029 ,n2028);
    not g5650(n2027 ,n2026);
    not g5651(n2025 ,n2024);
    not g5652(n2023 ,n2022);
    not g5653(n2021 ,n2020);
    not g5654(n2019 ,n2018);
    not g5655(n2017 ,n2016);
    not g5656(n2015 ,n2014);
    not g5657(n2013 ,n2012);
    not g5658(n2011 ,n2010);
    not g5659(n2009 ,n2008);
    not g5660(n2007 ,n2006);
    not g5661(n2005 ,n2004);
    not g5662(n2002 ,n2001);
    not g5663(n2000 ,n1999);
    xnor g5664(n1998 ,n1[49] ,n2[49]);
    xnor g5665(n1997 ,n1[122] ,n2[58]);
    xnor g5666(n1996 ,n1[101] ,n2[37]);
    xnor g5667(n1995 ,n1[117] ,n2[53]);
    xnor g5668(n1994 ,n1[84] ,n2[20]);
    xnor g5669(n1993 ,n1[30] ,n2[30]);
    xnor g5670(n1992 ,n1[93] ,n2[29]);
    xnor g5671(n1991 ,n1[89] ,n2[25]);
    xnor g5672(n1990 ,n1[98] ,n2[34]);
    xnor g5673(n1989 ,n1[102] ,n2[38]);
    xnor g5674(n1988 ,n1[75] ,n2[11]);
    xnor g5675(n1987 ,n1[0] ,n2[0]);
    xnor g5676(n1986 ,n1[18] ,n2[18]);
    xnor g5677(n1985 ,n1[105] ,n2[41]);
    xnor g5678(n1984 ,n1[107] ,n2[43]);
    xnor g5679(n1983 ,n1[109] ,n2[45]);
    xnor g5680(n1982 ,n1[31] ,n2[31]);
    xnor g5681(n1981 ,n1[111] ,n2[47]);
    xnor g5682(n1980 ,n1[100] ,n2[36]);
    xnor g5683(n1979 ,n1[114] ,n2[50]);
    xnor g5684(n1978 ,n1[15] ,n2[15]);
    xnor g5685(n1977 ,n1[27] ,n2[27]);
    xnor g5686(n1976 ,n1[103] ,n2[39]);
    xnor g5687(n1975 ,n1[3] ,n2[3]);
    xnor g5688(n1974 ,n1[11] ,n2[11]);
    xnor g5689(n1973 ,n1[110] ,n2[46]);
    xnor g5690(n1972 ,n1[118] ,n2[54]);
    xnor g5691(n1971 ,n1[99] ,n2[35]);
    xnor g5692(n1970 ,n1[10] ,n2[10]);
    xnor g5693(n1969 ,n1[1] ,n2[1]);
    xnor g5694(n1968 ,n1[2] ,n2[2]);
    xnor g5695(n1967 ,n1[106] ,n2[42]);
    xnor g5696(n1966 ,n1[19] ,n2[19]);
    xnor g5697(n1965 ,n1[125] ,n2[61]);
    xnor g5698(n1964 ,n1[70] ,n2[6]);
    xnor g5699(n1963 ,n1[73] ,n2[9]);
    xnor g5700(n1962 ,n1[68] ,n2[4]);
    xnor g5701(n1961 ,n1[29] ,n2[29]);
    xnor g5702(n1960 ,n1[72] ,n2[8]);
    xnor g5703(n1959 ,n1[79] ,n2[15]);
    xnor g5704(n1958 ,n1[76] ,n2[12]);
    xnor g5705(n1957 ,n1[88] ,n2[24]);
    xnor g5706(n1956 ,n1[5] ,n2[5]);
    xnor g5707(n1955 ,n1[22] ,n2[22]);
    xnor g5708(n1954 ,n1[24] ,n2[24]);
    xnor g5709(n1953 ,n1[81] ,n2[17]);
    xnor g5710(n1952 ,n1[71] ,n2[7]);
    xnor g5711(n1951 ,n1[115] ,n2[51]);
    xnor g5712(n1950 ,n1[28] ,n2[28]);
    xnor g5713(n1949 ,n1[124] ,n2[60]);
    xnor g5714(n1948 ,n1[6] ,n2[6]);
    xnor g5715(n1947 ,n1[91] ,n2[27]);
    xnor g5716(n1946 ,n1[126] ,n2[62]);
    xnor g5717(n1945 ,n1[92] ,n2[28]);
    xnor g5718(n1944 ,n1[77] ,n2[13]);
    xnor g5719(n1943 ,n1[64] ,n2[0]);
    xnor g5720(n1942 ,n1[94] ,n2[30]);
    xnor g5721(n1941 ,n1[95] ,n2[31]);
    xnor g5722(n1940 ,n1[12] ,n2[12]);
    xnor g5723(n1939 ,n1[23] ,n2[23]);
    xnor g5724(n1938 ,n1[9] ,n2[9]);
    xnor g5725(n1937 ,n1[104] ,n2[40]);
    xnor g5726(n1936 ,n1[13] ,n2[13]);
    xnor g5727(n1935 ,n1[96] ,n2[32]);
    xnor g5728(n1934 ,n1[4] ,n2[4]);
    xnor g5729(n1933 ,n1[14] ,n2[14]);
    xnor g5730(n1932 ,n1[20] ,n2[20]);
    xnor g5731(n1931 ,n1[25] ,n2[25]);
    xnor g5732(n1930 ,n1[108] ,n2[44]);
    xnor g5733(n1929 ,n1[26] ,n2[26]);
    xnor g5734(n1928 ,n1[113] ,n2[49]);
    xnor g5735(n1927 ,n1[16] ,n2[16]);
    xnor g5736(n1926 ,n1[21] ,n2[21]);
    xnor g5737(n1925 ,n1[69] ,n2[5]);
    xnor g5738(n1924 ,n1[121] ,n2[57]);
    xnor g5739(n1923 ,n1[17] ,n2[17]);
    xnor g5740(n1922 ,n1[67] ,n2[3]);
    xnor g5741(n1921 ,n1[7] ,n2[7]);
    xnor g5742(n1920 ,n1[74] ,n2[10]);
    xnor g5743(n1919 ,n1[8] ,n2[8]);
    xnor g5744(n1918 ,n1[127] ,n2[63]);
    xnor g5745(n1917 ,n1[66] ,n2[2]);
    xnor g5746(n1916 ,n1[63] ,n2[63]);
    xnor g5747(n1915 ,n1[62] ,n2[62]);
    xnor g5748(n1914 ,n1[120] ,n2[56]);
    xnor g5749(n1913 ,n1[116] ,n2[52]);
    xnor g5750(n1912 ,n1[97] ,n2[33]);
    xnor g5751(n1911 ,n1[38] ,n2[38]);
    xnor g5752(n1910 ,n1[86] ,n2[22]);
    xnor g5753(n1909 ,n1[83] ,n2[19]);
    xnor g5754(n1908 ,n1[34] ,n2[34]);
    xnor g5755(n1907 ,n1[59] ,n2[59]);
    xnor g5756(n1906 ,n1[42] ,n2[42]);
    xnor g5757(n1905 ,n1[58] ,n2[58]);
    xnor g5758(n1904 ,n1[85] ,n2[21]);
    xnor g5759(n1903 ,n1[61] ,n2[61]);
    xnor g5760(n1902 ,n1[60] ,n2[60]);
    xnor g5761(n1901 ,n1[32] ,n2[32]);
    xnor g5762(n1900 ,n1[80] ,n2[16]);
    xnor g5763(n1899 ,n1[35] ,n2[35]);
    xnor g5764(n1898 ,n1[119] ,n2[55]);
    xnor g5765(n1897 ,n1[36] ,n2[36]);
    xnor g5766(n1896 ,n1[37] ,n2[37]);
    xnor g5767(n1895 ,n1[39] ,n2[39]);
    xnor g5768(n1894 ,n1[40] ,n2[40]);
    xnor g5769(n1893 ,n1[41] ,n2[41]);
    xnor g5770(n1892 ,n1[44] ,n2[44]);
    xnor g5771(n1891 ,n1[45] ,n2[45]);
    xnor g5772(n1890 ,n1[46] ,n2[46]);
    xnor g5773(n1889 ,n1[48] ,n2[48]);
    xnor g5774(n1888 ,n1[57] ,n2[57]);
    xnor g5775(n1887 ,n1[51] ,n2[51]);
    xnor g5776(n1886 ,n1[52] ,n2[52]);
    xnor g5777(n1885 ,n1[87] ,n2[23]);
    xnor g5778(n1884 ,n1[47] ,n2[47]);
    xnor g5779(n1883 ,n1[33] ,n2[33]);
    xnor g5780(n1882 ,n1[43] ,n2[43]);
    xnor g5781(n1881 ,n1[56] ,n2[56]);
    xnor g5782(n1880 ,n1[50] ,n2[50]);
    xnor g5783(n1879 ,n7435 ,n7434);
    xnor g5784(n1878 ,n7495 ,n7494);
    xnor g5785(n1877 ,n7416 ,n7417);
    xnor g5786(n1876 ,n1[35] ,n4[27]);
    xnor g5787(n1875 ,n7456 ,n7457);
    xnor g5788(n1874 ,n7504 ,n7503);
    xnor g5789(n1873 ,n7423 ,n7422);
    xnor g5790(n1872 ,n7669 ,n7627);
    xnor g5791(n1871 ,n7412 ,n7413);
    xnor g5792(n1870 ,n7524 ,n7525);
    xnor g5793(n1869 ,n1[119] ,n4[15]);
    xnor g5794(n1868 ,n7449 ,n7447);
    xnor g5795(n1867 ,n7523 ,n7522);
    xnor g5796(n1866 ,n7444 ,n7445);
    xnor g5797(n1865 ,n7451 ,n7450);
    xnor g5798(n1864 ,n7468 ,n7469);
    xnor g5799(n1863 ,n7667 ,n7625);
    xnor g5800(n1862 ,n7480 ,n7481);
    xnor g5801(n1861 ,n1[36] ,n1[4]);
    xnor g5802(n1860 ,n7559 ,n7526);
    xnor g5803(n1859 ,n1[42] ,n1[10]);
    xnor g5804(n1858 ,n7452 ,n7453);
    xnor g5805(n1857 ,n7520 ,n7521);
    xnor g5806(n1856 ,n7479 ,n7478);
    xnor g5807(n1855 ,n7436 ,n7437);
    xnor g5808(n1854 ,n7428 ,n7429);
    xnor g5809(n1853 ,n0[80] ,n7682);
    xnor g5810(n1852 ,n0[82] ,n7684);
    xnor g5811(n1851 ,n0[104] ,n7674);
    xnor g5812(n1850 ,n0[89] ,n7691);
    xnor g5813(n1849 ,n0[83] ,n7685);
    xnor g5814(n1848 ,n0[122] ,n7692);
    xnor g5815(n1847 ,n0[107] ,n7677);
    xnor g5816(n1846 ,n0[88] ,n7690);
    xnor g5817(n1845 ,n0[91] ,n7693);
    xnor g5818(n1844 ,n0[73] ,n7675);
    xnor g5819(n1843 ,n0[113] ,n7683);
    xnor g5820(n1842 ,n0[102] ,n7672);
    xnor g5821(n1841 ,n0[79] ,n7681);
    xnor g5822(n1840 ,n0[78] ,n7680);
    xnor g5823(n1839 ,n7666 ,n7624);
    xnor g5824(n1838 ,n0[77] ,n7679);
    xnor g5825(n1837 ,n0[76] ,n7678);
    xnor g5826(n1836 ,n7419 ,n7418);
    xnor g5827(n1835 ,n0[95] ,n7697);
    xnor g5828(n1834 ,n0[92] ,n7694);
    xnor g5829(n1833 ,n0[94] ,n7696);
    xnor g5830(n1832 ,n7420 ,n7421);
    xnor g5831(n1831 ,n0[68] ,n7670);
    xnor g5832(n1830 ,n0[69] ,n7671);
    xnor g5833(n1829 ,n0[71] ,n7673);
    xnor g5834(n1828 ,n0[93] ,n7695);
    xnor g5835(n1827 ,n0[84] ,n7686);
    xnor g5836(n1826 ,n7628 ,n7629);
    xnor g5837(n1825 ,n7668 ,n7626);
    xnor g5838(n1824 ,n0[86] ,n7688);
    xnor g5839(n1823 ,n7511 ,n7510);
    xnor g5840(n1822 ,n7475 ,n7474);
    xnor g5841(n1821 ,n7427 ,n7426);
    xnor g5842(n1820 ,n7440 ,n7441);
    xnor g5843(n1819 ,n1[116] ,n4[12]);
    xnor g5844(n1818 ,n7519 ,n7518);
    xnor g5845(n1817 ,n7431 ,n7430);
    xnor g5846(n1816 ,n7432 ,n7433);
    xnor g5847(n1815 ,n7439 ,n7438);
    xnor g5848(n1814 ,n7424 ,n7425);
    xnor g5849(n1813 ,n0[22] ,n4[30]);
    xnor g5850(n1812 ,n0[3] ,n4[19]);
    xnor g5851(n1811 ,n7411 ,n7410);
    xnor g5852(n1810 ,n0[85] ,n7687);
    xnor g5853(n1809 ,n0[125] ,n4[13]);
    xnor g5854(n1808 ,n0[126] ,n4[14]);
    xnor g5855(n1807 ,n7472 ,n7471);
    xnor g5856(n1806 ,n7443 ,n7442);
    xnor g5857(n1805 ,n0[6] ,n4[22]);
    xnor g5858(n1804 ,n0[23] ,n4[31]);
    xnor g5859(n1803 ,n0[21] ,n4[29]);
    xnor g5860(n1802 ,n7493 ,n7491);
    xnor g5861(n1801 ,n0[92] ,n4[20]);
    xnor g5862(n1800 ,n0[127] ,n4[15]);
    xnor g5863(n1799 ,n0[95] ,n4[23]);
    xnor g5864(n1798 ,n0[87] ,n7689);
    xnor g5865(n1797 ,n7448 ,n7446);
    xnor g5866(n1796 ,n0[93] ,n4[21]);
    xnor g5867(n1795 ,n7512 ,n7513);
    xnor g5868(n1794 ,n7508 ,n7509);
    xnor g5869(n1793 ,n0[94] ,n4[22]);
    xnor g5870(n1792 ,n7500 ,n7501);
    xnor g5871(n1791 ,n7455 ,n7454);
    xnor g5872(n1790 ,n7460 ,n7461);
    xnor g5873(n1789 ,n7415 ,n7414);
    xnor g5874(n1788 ,n7459 ,n7458);
    xnor g5875(n1787 ,n0[15] ,n4[31]);
    xnor g5876(n1786 ,n7404 ,n7402);
    xnor g5877(n1785 ,n7487 ,n7486);
    xnor g5878(n1784 ,n7505 ,n7502);
    xnor g5879(n1783 ,n7464 ,n7462);
    xnor g5880(n1782 ,n0[124] ,n4[12]);
    xnor g5881(n1781 ,n0[36] ,n1[52]);
    xnor g5882(n1780 ,n7465 ,n7463);
    xnor g5883(n1779 ,n0[37] ,n1[53]);
    xnor g5884(n1778 ,n0[44] ,n1[60]);
    xnor g5885(n1777 ,n0[45] ,n1[61]);
    xnor g5886(n1776 ,n0[46] ,n1[62]);
    xnor g5887(n1775 ,n0[47] ,n1[63]);
    xnor g5888(n1774 ,n1[56] ,n1[24]);
    xnor g5889(n1773 ,n7467 ,n7466);
    xnor g5890(n1772 ,n0[4] ,n4[20]);
    xnor g5891(n1771 ,n7405 ,n7403);
    xnor g5892(n1770 ,n7473 ,n7470);
    xnor g5893(n1769 ,n7492 ,n7490);
    xnor g5894(n1768 ,n7407 ,n7406);
    xnor g5895(n1767 ,n7515 ,n7514);
    xnor g5896(n1766 ,n1[55] ,n1[23]);
    xnor g5897(n1765 ,n0[38] ,n1[54]);
    xnor g5898(n1764 ,n7476 ,n7477);
    xnor g5899(n1763 ,n7516 ,n7517);
    xnor g5900(n1762 ,n0[14] ,n4[30]);
    xnor g5901(n1761 ,n0[102] ,n4[14]);
    xnor g5902(n1760 ,n7499 ,n7498);
    xnor g5903(n1759 ,n0[101] ,n4[13]);
    xnor g5904(n1758 ,n0[98] ,n4[10]);
    xnor g5905(n1757 ,n7507 ,n7506);
    xnor g5906(n1756 ,n0[96] ,n4[8]);
    xnor g5907(n1755 ,n0[99] ,n4[11]);
    xnor g5908(n1754 ,n1[97] ,n4[25]);
    xnor g5909(n1753 ,n1[40] ,n4[0]);
    xnor g5910(n1752 ,n1[120] ,n4[0]);
    xnor g5911(n1751 ,n7484 ,n7485);
    xnor g5912(n1750 ,n0[91] ,n4[19]);
    xnor g5913(n1749 ,n7483 ,n7482);
    xnor g5914(n1748 ,n7488 ,n7489);
    xnor g5915(n1747 ,n7496 ,n7497);
    xnor g5916(n1746 ,n7408 ,n7409);
    xnor g5917(n2136 ,n0[95] ,n1[95]);
    xnor g5918(n2135 ,n0[117] ,n1[117]);
    xnor g5919(n2134 ,n0[37] ,n1[37]);
    xnor g5920(n2133 ,n0[108] ,n1[108]);
    xnor g5921(n2132 ,n0[65] ,n1[65]);
    xnor g5922(n2131 ,n0[111] ,n1[111]);
    xnor g5923(n2130 ,n0[93] ,n1[93]);
    xnor g5924(n2129 ,n0[84] ,n1[84]);
    xnor g5925(n2128 ,n0[125] ,n1[125]);
    xnor g5926(n2127 ,n0[76] ,n1[76]);
    xnor g5927(n2126 ,n0[77] ,n1[77]);
    xnor g5928(n2125 ,n0[79] ,n1[79]);
    xnor g5929(n2124 ,n0[68] ,n1[68]);
    xnor g5930(n2123 ,n0[118] ,n1[118]);
    xnor g5931(n2122 ,n0[69] ,n1[69]);
    xnor g5932(n2121 ,n0[67] ,n1[67]);
    xnor g5933(n2120 ,n0[98] ,n1[98]);
    xnor g5934(n2119 ,n0[99] ,n1[99]);
    xnor g5935(n2118 ,n0[102] ,n1[102]);
    xnor g5936(n2117 ,n0[101] ,n1[101]);
    xnor g5937(n2116 ,n0[96] ,n1[96]);
    xnor g5938(n2115 ,n0[109] ,n1[109]);
    xnor g5939(n2114 ,n0[127] ,n1[127]);
    xnor g5940(n2113 ,n0[94] ,n1[94]);
    xnor g5941(n2112 ,n0[39] ,n1[39]);
    xnor g5942(n2111 ,n0[38] ,n1[38]);
    xnor g5943(n2110 ,n0[66] ,n1[66]);
    xnor g5944(n2109 ,n0[103] ,n1[103]);
    xnor g5945(n2108 ,n0[124] ,n1[124]);
    xnor g5946(n2107 ,n0[46] ,n1[46]);
    xnor g5947(n2106 ,n0[36] ,n1[36]);
    xnor g5948(n2105 ,n0[44] ,n1[44]);
    xnor g5949(n2104 ,n0[64] ,n1[64]);
    xnor g5950(n2103 ,n0[45] ,n1[45]);
    xnor g5951(n2102 ,n0[47] ,n1[47]);
    xnor g5952(n2101 ,n0[70] ,n1[70]);
    xnor g5953(n2100 ,n0[92] ,n1[92]);
    xnor g5954(n2099 ,n0[71] ,n1[71]);
    xnor g5955(n2098 ,n0[91] ,n1[91]);
    xnor g5956(n2097 ,n0[110] ,n1[110]);
    xnor g5957(n2096 ,n0[100] ,n1[100]);
    xnor g5958(n2095 ,n0[126] ,n1[126]);
    xnor g5959(n2094 ,n0[78] ,n1[78]);
    xnor g5960(n2092 ,n1[12] ,n1285);
    xnor g5961(n2091 ,n0[57] ,n4[17]);
    xnor g5962(n2090 ,n0[2] ,n1[2]);
    xnor g5963(n2089 ,n0[48] ,n4[8]);
    xnor g5964(n2088 ,n0[14] ,n1[14]);
    xnor g5965(n2087 ,n0[59] ,n4[19]);
    xnor g5966(n2086 ,n0[56] ,n4[16]);
    xnor g5967(n2085 ,n0[26] ,n1[26]);
    xnor g5968(n2084 ,n0[51] ,n4[11]);
    xnor g5969(n2083 ,n0[49] ,n4[9]);
    xnor g5970(n2081 ,n1[18] ,n1258);
    xnor g5971(n2079 ,n1[3] ,n1146);
    xnor g5972(n2078 ,n0[53] ,n4[13]);
    xnor g5973(n2076 ,n1[11] ,n1267);
    xnor g5974(n2075 ,n0[22] ,n1[22]);
    xnor g5975(n2074 ,n0[20] ,n1[20]);
    xnor g5976(n2073 ,n0[28] ,n1[28]);
    xnor g5977(n2072 ,n0[29] ,n1[29]);
    xnor g5978(n2071 ,n0[15] ,n1[15]);
    xnor g5979(n2070 ,n0[13] ,n1[13]);
    xnor g5980(n2069 ,n0[12] ,n1[12]);
    xnor g5981(n2068 ,n0[31] ,n1[31]);
    xnor g5982(n2067 ,n0[5] ,n1[5]);
    xnor g5983(n2066 ,n0[50] ,n4[10]);
    xnor g5984(n2065 ,n0[7] ,n1[7]);
    xnor g5985(n2064 ,n0[21] ,n1[21]);
    xnor g5986(n2063 ,n0[30] ,n1[30]);
    xnor g5987(n2061 ,n1[22] ,n1122);
    xnor g5988(n2060 ,n0[6] ,n1[6]);
    xnor g5989(n2058 ,n1[29] ,n1300);
    xnor g5990(n2056 ,n1[6] ,n1287);
    xnor g5991(n2054 ,n1[1] ,n1296);
    xnor g5992(n2052 ,n1[27] ,n1136);
    xnor g5993(n2050 ,n1[25] ,n1135);
    xnor g5994(n2049 ,n0[18] ,n1[18]);
    xnor g5995(n2047 ,n1[2] ,n1141);
    xnor g5996(n2046 ,n0[55] ,n4[15]);
    xnor g5997(n2044 ,n1[28] ,n1140);
    xnor g5998(n2043 ,n0[52] ,n4[12]);
    xnor g5999(n2041 ,n1[26] ,n1132);
    xnor g6000(n2040 ,n0[87] ,n4[31]);
    xnor g6001(n2038 ,n1[16] ,n1130);
    xnor g6002(n2036 ,n1[0] ,n1142);
    xnor g6003(n2035 ,n0[54] ,n4[14]);
    xnor g6004(n2034 ,n0[61] ,n4[21]);
    xnor g6005(n2033 ,n0[60] ,n4[20]);
    xnor g6006(n2032 ,n0[62] ,n4[22]);
    xnor g6007(n2031 ,n0[63] ,n4[23]);
    xnor g6008(n2030 ,n0[86] ,n4[30]);
    xnor g6009(n2028 ,n1[5] ,n1134);
    xnor g6010(n2026 ,n1[8] ,n1133);
    xnor g6011(n2024 ,n1[7] ,n1143);
    xnor g6012(n2022 ,n1[13] ,n1286);
    xnor g6013(n2020 ,n1[15] ,n1129);
    xnor g6014(n2018 ,n1[30] ,n1290);
    xnor g6015(n2016 ,n1[46] ,n1[14]);
    xnor g6016(n2014 ,n1[17] ,n1125);
    xnor g6017(n2012 ,n1[19] ,n1297);
    xnor g6018(n2010 ,n1[20] ,n1295);
    xnor g6019(n2008 ,n1[21] ,n1294);
    xnor g6020(n2006 ,n1[9] ,n1292);
    xnor g6021(n2004 ,n1[31] ,n1293);
    xnor g6022(n2003 ,n0[85] ,n4[29]);
    xnor g6023(n2001 ,n1[4] ,n1105);
    xnor g6024(n1999 ,n1[23] ,n1112);
    not g6025(n1745 ,n1744);
    not g6026(n1742 ,n1741);
    not g6027(n1738 ,n1737);
    not g6028(n1735 ,n1734);
    not g6029(n1033 ,n1731);
    not g6030(n11 ,n1031);
    not g6031(n1730 ,n1031);
    not g6032(n1729 ,n1031);
    not g6033(n1031 ,n1032);
    nor g6034(n1728 ,n1177 ,n1017);
    nor g6035(n1727 ,n1279 ,n1025);
    nor g6036(n1726 ,n1224 ,n1182);
    nor g6037(n1725 ,n1272 ,n1025);
    nor g6038(n1724 ,n1310 ,n1314);
    nor g6039(n1723 ,n1309 ,n1161);
    nor g6040(n1722 ,n1308 ,n1311);
    nor g6041(n1721 ,n1157 ,n1159);
    nor g6042(n1720 ,n1154 ,n1312);
    nor g6043(n1719 ,n1127 ,n1315);
    nor g6044(n1718 ,n1294 ,n1313);
    nor g6045(n1717 ,n1122 ,n1163);
    nor g6046(n1716 ,n1265 ,n1160);
    nor g6047(n1715 ,n1278 ,n1025);
    nor g6048(n1714 ,n1196 ,n1019);
    nor g6049(n1713 ,n1340 ,n1019);
    nor g6050(n1712 ,n1201 ,n1019);
    nor g6051(n1711 ,n1178 ,n1017);
    nor g6052(n1710 ,n1181 ,n1018);
    nor g6053(n1709 ,n1316 ,n1018);
    nor g6054(n1708 ,n1195 ,n1018);
    nor g6055(n1707 ,n1217 ,n1017);
    nor g6056(n1706 ,n1174 ,n1019);
    nor g6057(n1705 ,n1339 ,n1018);
    nor g6058(n1704 ,n1168 ,n1019);
    nor g6059(n1703 ,n1330 ,n1017);
    nor g6060(n1702 ,n1348 ,n1019);
    nor g6061(n1701 ,n1165 ,n1019);
    nor g6062(n1700 ,n1345 ,n1018);
    nor g6063(n1699 ,n1337 ,n1017);
    nor g6064(n1698 ,n1214 ,n1018);
    nor g6065(n1697 ,n1200 ,n1017);
    nor g6066(n1696 ,n1347 ,n1017);
    nor g6067(n1695 ,n1344 ,n1018);
    nor g6068(n1694 ,n1328 ,n1019);
    nor g6069(n1693 ,n1215 ,n1017);
    nor g6070(n1692 ,n1197 ,n1017);
    nor g6071(n1691 ,n1334 ,n1017);
    nor g6072(n1690 ,n1198 ,n1018);
    nor g6073(n1689 ,n1342 ,n1017);
    nor g6074(n1688 ,n1205 ,n1019);
    nor g6075(n1687 ,n1212 ,n1019);
    nor g6076(n1686 ,n1166 ,n1018);
    nor g6077(n1685 ,n1327 ,n1019);
    nor g6078(n1684 ,n1209 ,n1018);
    nor g6079(n1683 ,n1176 ,n1018);
    nor g6080(n1682 ,n1173 ,n1019);
    nor g6081(n1681 ,n1343 ,n1017);
    nor g6082(n1680 ,n1320 ,n1017);
    nor g6083(n1679 ,n1352 ,n1018);
    nor g6084(n1678 ,n1341 ,n1017);
    nor g6085(n1677 ,n1323 ,n1018);
    nor g6086(n1676 ,n1187 ,n1018);
    nor g6087(n1675 ,n1336 ,n1018);
    nor g6088(n1674 ,n1188 ,n1019);
    nor g6089(n1673 ,n1333 ,n1017);
    nor g6090(n1672 ,n1189 ,n1019);
    nor g6091(n1671 ,n1355 ,n1019);
    nor g6092(n1670 ,n1213 ,n1018);
    nor g6093(n1669 ,n1338 ,n1018);
    nor g6094(n1668 ,n1321 ,n1017);
    nor g6095(n1667 ,n1190 ,n1018);
    nor g6096(n1666 ,n1346 ,n1019);
    nor g6097(n1665 ,n1192 ,n1018);
    nor g6098(n1664 ,n1319 ,n1018);
    nor g6099(n1663 ,n1186 ,n1018);
    nor g6100(n1662 ,n1354 ,n1018);
    nor g6101(n1661 ,n1218 ,n1018);
    nor g6102(n1660 ,n1183 ,n1019);
    nor g6103(n1659 ,n1194 ,n1018);
    nor g6104(n1658 ,n1350 ,n1017);
    nor g6105(n1657 ,n1317 ,n1017);
    nor g6106(n1656 ,n1171 ,n1017);
    nor g6107(n1655 ,n1185 ,n1018);
    nor g6108(n1654 ,n1322 ,n1018);
    nor g6109(n1653 ,n1204 ,n1017);
    nor g6110(n1652 ,n1220 ,n1017);
    nor g6111(n1651 ,n1169 ,n1018);
    nor g6112(n1650 ,n1199 ,n1018);
    nor g6113(n1649 ,n1324 ,n1018);
    nor g6114(n1648 ,n1193 ,n1019);
    nor g6115(n1647 ,n1325 ,n1017);
    nor g6116(n1646 ,n1329 ,n1017);
    nor g6117(n1645 ,n1191 ,n1017);
    nor g6118(n1644 ,n1349 ,n1018);
    nor g6119(n1643 ,n1222 ,n1017);
    nor g6120(n1642 ,n1179 ,n1018);
    nor g6121(n1641 ,n1216 ,n1019);
    nor g6122(n1640 ,n1206 ,n1019);
    nor g6123(n1639 ,n1167 ,n1018);
    or g6124(n1638 ,n1162 ,n3[1]);
    nor g6125(n1637 ,n1208 ,n1019);
    nor g6126(n1636 ,n1331 ,n1017);
    nor g6127(n1635 ,n1110 ,n1023);
    nor g6128(n1634 ,n1210 ,n1019);
    nor g6129(n1633 ,n1202 ,n1017);
    nor g6130(n1632 ,n1221 ,n1019);
    nor g6131(n1631 ,n1211 ,n1017);
    nor g6132(n1630 ,n1184 ,n1019);
    nor g6133(n1629 ,n1326 ,n1017);
    nor g6134(n1628 ,n1219 ,n1019);
    nor g6135(n1627 ,n1175 ,n1019);
    nor g6136(n1626 ,n1332 ,n1017);
    nor g6137(n1625 ,n1318 ,n1019);
    nor g6138(n1624 ,n1207 ,n1017);
    nor g6139(n1623 ,n1353 ,n1019);
    nor g6140(n1622 ,n1335 ,n1019);
    nor g6141(n1621 ,n1180 ,n1019);
    nor g6142(n1620 ,n1164 ,n1019);
    nor g6143(n1619 ,n1172 ,n1017);
    nor g6144(n1618 ,n1203 ,n1019);
    nor g6145(n1617 ,n1276 ,n1023);
    nor g6146(n1616 ,n1283 ,n1025);
    nor g6147(n1615 ,n1104 ,n1260);
    nor g6148(n1614 ,n1247 ,n1245);
    nor g6149(n1613 ,n1248 ,n1250);
    nor g6150(n1612 ,n1112 ,n1023);
    nor g6151(n1611 ,n1239 ,n1252);
    nor g6152(n1610 ,n1124 ,n1025);
    nor g6153(n1609 ,n1241 ,n1244);
    nor g6154(n1608 ,n1089 ,n1084);
    nor g6155(n1607 ,n1269 ,n1023);
    nor g6156(n1606 ,n1082 ,n1072);
    nor g6157(n1605 ,n1078 ,n1238);
    nor g6158(n1604 ,n1230 ,n1074);
    nor g6159(n1603 ,n1234 ,n1235);
    or g6160(n1602 ,n1079 ,n1231);
    nor g6161(n1601 ,n1073 ,n1232);
    nor g6162(n1600 ,n1075 ,n1080);
    nor g6163(n1599 ,n1114 ,n1023);
    nor g6164(n1598 ,n1242 ,n1227);
    nor g6165(n1597 ,n1147 ,n1023);
    nor g6166(n1596 ,n1304 ,n1023);
    nor g6167(n1595 ,n1152 ,n1025);
    nor g6168(n1594 ,n1149 ,n1025);
    nor g6169(n1593 ,n1148 ,n1025);
    nor g6170(n1592 ,n1301 ,n1025);
    nor g6171(n1591 ,n1302 ,n1023);
    nor g6172(n1590 ,n1151 ,n1025);
    nor g6173(n1589 ,n1153 ,n1025);
    nor g6174(n1588 ,n1305 ,n1025);
    nor g6175(n1587 ,n1306 ,n1023);
    nor g6176(n1586 ,n1303 ,n1023);
    nor g6177(n1585 ,n1150 ,n1028);
    nor g6178(n1584 ,n1149 ,n1024);
    nor g6179(n1583 ,n1148 ,n1022);
    nor g6180(n1582 ,n1302 ,n1022);
    nor g6181(n1581 ,n1147 ,n1022);
    nor g6182(n1580 ,n1153 ,n1022);
    nor g6183(n1579 ,n1301 ,n1024);
    nor g6184(n1578 ,n1306 ,n1024);
    nor g6185(n1577 ,n1152 ,n1024);
    nor g6186(n1576 ,n1151 ,n1024);
    nor g6187(n1575 ,n1305 ,n1024);
    nor g6188(n1574 ,n1304 ,n1024);
    nor g6189(n1573 ,n1303 ,n1022);
    nor g6190(n1572 ,n1126 ,n1023);
    nor g6191(n1571 ,n1299 ,n1023);
    nor g6192(n1570 ,n1131 ,n1023);
    nor g6193(n1569 ,n1289 ,n1028);
    nor g6194(n1568 ,n1131 ,n1024);
    nor g6195(n1567 ,n1299 ,n1022);
    nor g6196(n1566 ,n1138 ,n1030);
    nor g6197(n1565 ,n1291 ,n1027);
    nor g6198(n1564 ,n1126 ,n1024);
    nor g6199(n1563 ,n1271 ,n1023);
    nor g6200(n1562 ,n1118 ,n1023);
    nor g6201(n1561 ,n1274 ,n1023);
    nor g6202(n1560 ,n1111 ,n1023);
    nor g6203(n1559 ,n1119 ,n1025);
    nor g6204(n1558 ,n1123 ,n1023);
    nor g6205(n1557 ,n1117 ,n1023);
    nor g6206(n1556 ,n1281 ,n1023);
    nor g6207(n1555 ,n1120 ,n1023);
    nor g6208(n1554 ,n1121 ,n1023);
    nor g6209(n1744 ,n1266 ,n1095);
    or g6210(n1743 ,n1092 ,n1242);
    nor g6211(n1741 ,n1249 ,n1237);
    nor g6212(n1740 ,n1282 ,n1023);
    nor g6213(n1739 ,n1284 ,n1025);
    nor g6214(n1737 ,n1087 ,n1249);
    nor g6215(n1736 ,n1091 ,n1227);
    nor g6216(n1734 ,n1262 ,n1266);
    or g6217(n1733 ,n1351 ,n1223);
    or g6218(n1732 ,n1162 ,n1170);
    or g6219(n1731 ,n1225 ,n1356);
    or g6220(n1032 ,n1351 ,n1162);
    not g6221(n1553 ,n1552);
    not g6222(n1542 ,n1541);
    not g6223(n1539 ,n1538);
    not g6224(n1535 ,n1534);
    not g6225(n1531 ,n1530);
    not g6226(n1529 ,n1528);
    not g6227(n1526 ,n1525);
    not g6228(n1522 ,n1521);
    not g6229(n1520 ,n1519);
    nor g6230(n1512 ,n1277 ,n1025);
    nor g6231(n1511 ,n1108 ,n1023);
    nor g6232(n1510 ,n1268 ,n1023);
    nor g6233(n1509 ,n1107 ,n1025);
    nor g6234(n1508 ,n1116 ,n1025);
    nor g6235(n1507 ,n1115 ,n1025);
    nor g6236(n1506 ,n1109 ,n1025);
    nor g6237(n1505 ,n1273 ,n1025);
    nor g6238(n1504 ,n1113 ,n1023);
    nor g6239(n1503 ,n1275 ,n1023);
    nor g6240(n1502 ,n1280 ,n1023);
    nor g6241(n1501 ,n1108 ,n1022);
    nor g6242(n1500 ,n1113 ,n1022);
    nor g6243(n1499 ,n1116 ,n1022);
    nor g6244(n1498 ,n1[54] ,n2[54]);
    nor g6245(n1497 ,n1115 ,n1024);
    nor g6246(n1496 ,n1284 ,n1022);
    nor g6247(n1495 ,n1121 ,n1024);
    nor g6248(n1494 ,n1119 ,n1022);
    nor g6249(n1493 ,n1280 ,n1022);
    nor g6250(n1492 ,n1114 ,n1022);
    nor g6251(n1491 ,n1118 ,n1024);
    nor g6252(n1490 ,n1271 ,n1022);
    nor g6253(n1489 ,n1279 ,n1024);
    nor g6254(n1488 ,n1107 ,n1022);
    nor g6255(n1487 ,n1272 ,n1024);
    nor g6256(n1486 ,n1270 ,n1030);
    nor g6257(n1485 ,n1282 ,n1024);
    nor g6258(n1484 ,n1274 ,n1024);
    nor g6259(n1483 ,n1281 ,n1024);
    nor g6260(n1482 ,n1123 ,n1024);
    nor g6261(n1481 ,n1112 ,n1024);
    nor g6262(n1480 ,n1273 ,n1022);
    nor g6263(n1479 ,n1266 ,n1067);
    nor g6264(n1478 ,n1[90] ,n2[26]);
    nor g6265(n1477 ,n1124 ,n1024);
    nor g6266(n1476 ,n1109 ,n1024);
    nor g6267(n1475 ,n1111 ,n1022);
    nor g6268(n1474 ,n1268 ,n1024);
    nor g6269(n1473 ,n1276 ,n1022);
    or g6270(n1472 ,n0[42] ,n0[40]);
    nor g6271(n1471 ,n1283 ,n1024);
    nor g6272(n1470 ,n1277 ,n1024);
    nor g6273(n1469 ,n1117 ,n1024);
    nor g6274(n1468 ,n1110 ,n1022);
    nor g6275(n1467 ,n1120 ,n1024);
    nor g6276(n1466 ,n0[19] ,n0[17]);
    nor g6277(n1465 ,n1261 ,n1030);
    nor g6278(n1464 ,n1260 ,n1066);
    nor g6279(n1463 ,n1256 ,n0[64]);
    nor g6280(n1462 ,n1262 ,n0[49]);
    nor g6281(n1461 ,n1256 ,n1067);
    nor g6282(n1460 ,n1264 ,n1066);
    nor g6283(n1459 ,n1259 ,n1028);
    nor g6284(n1458 ,n1263 ,n1028);
    nor g6285(n1457 ,n1105 ,n1022);
    nor g6286(n1456 ,n1254 ,n1030);
    nor g6287(n1455 ,n1106 ,n1028);
    nor g6288(n1454 ,n1103 ,n0[48]);
    nor g6289(n1453 ,n1264 ,n0[40]);
    nor g6290(n1452 ,n1255 ,n1066);
    nor g6291(n1451 ,n1257 ,n1030);
    nor g6292(n1450 ,n1104 ,n0[57]);
    nor g6293(n1449 ,n1255 ,n0[32]);
    or g6294(n1448 ,n1260 ,n0[57]);
    nor g6295(n1447 ,n1100 ,n1023);
    nor g6296(n1446 ,n1246 ,n1023);
    nor g6297(n1445 ,n1099 ,n1023);
    nor g6298(n1444 ,n1101 ,n1069);
    nor g6299(n1443 ,n1248 ,n0[65]);
    nor g6300(n1442 ,n0[48] ,n1069);
    nor g6301(n1441 ,n1247 ,n0[97]);
    nor g6302(n1440 ,n1246 ,n1024);
    nor g6303(n1439 ,n1100 ,n1024);
    nor g6304(n1438 ,n1094 ,n1067);
    nor g6305(n1437 ,n1098 ,n0[56]);
    or g6306(n1436 ,n0[34] ,n0[32]);
    nor g6307(n1435 ,n1251 ,n1067);
    nor g6308(n1434 ,n1[123] ,n2[59]);
    nor g6309(n1433 ,n1096 ,n1030);
    nor g6310(n1432 ,n1099 ,n1024);
    nor g6311(n1431 ,n1098 ,n1066);
    nor g6312(n1430 ,n1248 ,n0[66]);
    nor g6313(n1429 ,n1097 ,n1069);
    nor g6314(n1428 ,n1247 ,n0[98]);
    nor g6315(n1427 ,n1249 ,n1069);
    or g6316(n1426 ,n1084 ,n0[25]);
    nor g6317(n1425 ,n1083 ,n0[72]);
    nor g6318(n1424 ,n1090 ,n1067);
    nor g6319(n1423 ,n1085 ,n0[96]);
    nor g6320(n1422 ,n1082 ,n0[42]);
    nor g6321(n1421 ,n1087 ,n0[1]);
    nor g6322(n1420 ,n1082 ,n0[41]);
    nor g6323(n1419 ,n1240 ,n1068);
    nor g6324(n1418 ,n1088 ,n0[0]);
    nor g6325(n1417 ,n1084 ,n1069);
    nor g6326(n1416 ,n1093 ,n1068);
    nor g6327(n1415 ,n1083 ,n1066);
    nor g6328(n1414 ,n1243 ,n0[8]);
    or g6329(n1413 ,n1244 ,n0[89]);
    nor g6330(n1412 ,n1240 ,n0[80]);
    nor g6331(n1411 ,n1243 ,n1067);
    nor g6332(n1410 ,n1089 ,n0[25]);
    nor g6333(n1409 ,n1090 ,n0[104]);
    nor g6334(n1408 ,n1241 ,n0[89]);
    nor g6335(n1407 ,n1244 ,n1067);
    nor g6336(n1406 ,n1085 ,n1069);
    nor g6337(n1405 ,n1093 ,n0[112]);
    nor g6338(n1404 ,n1239 ,n0[33]);
    nor g6339(n1403 ,n1234 ,n0[74]);
    or g6340(n1402 ,n1231 ,n0[121]);
    nor g6341(n1401 ,n1[82] ,n2[18]);
    nor g6342(n1400 ,n1[55] ,n2[55]);
    nor g6343(n1399 ,n1073 ,n0[106]);
    nor g6344(n1398 ,n1071 ,n0[88]);
    nor g6345(n1397 ,n0[27] ,n0[25]);
    nor g6346(n1396 ,n1239 ,n0[34]);
    nor g6347(n1395 ,n1076 ,n0[24]);
    nor g6348(n1394 ,n1230 ,n0[114]);
    nor g6349(n1393 ,n1075 ,n0[9]);
    nor g6350(n1392 ,n1233 ,n1068);
    nor g6351(n1391 ,n1231 ,n1067);
    nor g6352(n1390 ,n1073 ,n0[105]);
    nor g6353(n1389 ,n1070 ,n1068);
    nor g6354(n1388 ,n1077 ,n1069);
    nor g6355(n1387 ,n1076 ,n1066);
    nor g6356(n1386 ,n1078 ,n0[81]);
    nor g6357(n1385 ,n1079 ,n0[121]);
    nor g6358(n1384 ,n0[91] ,n0[89]);
    nor g6359(n1383 ,n1[112] ,n2[48]);
    nor g6360(n1382 ,n1234 ,n0[73]);
    nor g6361(n1381 ,n1[78] ,n2[14]);
    nor g6362(n1380 ,n1230 ,n0[113]);
    nor g6363(n1379 ,n1071 ,n1069);
    nor g6364(n1378 ,n1081 ,n1068);
    nor g6365(n1377 ,n1078 ,n0[82]);
    nor g6366(n1376 ,n1075 ,n0[10]);
    nor g6367(n1375 ,n0[59] ,n0[57]);
    nor g6368(n1374 ,n1229 ,n0[120]);
    nor g6369(n1373 ,n1229 ,n1068);
    nor g6370(n1372 ,n1228 ,n1066);
    nor g6371(n1371 ,n0[0] ,n1068);
    nor g6372(n1370 ,n0[16] ,n1066);
    or g6373(n1369 ,n0[114] ,n0[112]);
    or g6374(n1368 ,n1020 ,n0[123]);
    or g6375(n1367 ,n0[66] ,n0[64]);
    or g6376(n1366 ,n0[82] ,n0[80]);
    nor g6377(n1365 ,n1[65] ,n2[1]);
    nor g6378(n1364 ,n0[122] ,n0[120]);
    nor g6379(n1363 ,n0[123] ,n0[121]);
    or g6380(n1362 ,n0[74] ,n0[72]);
    nor g6381(n1361 ,n0[18] ,n1068);
    nor g6382(n1360 ,n1[53] ,n2[53]);
    or g6383(n1359 ,n0[106] ,n0[104]);
    or g6384(n1358 ,n0[98] ,n0[96]);
    or g6385(n1357 ,n0[10] ,n0[8]);
    nor g6386(n1552 ,n1238 ,n0[81]);
    nor g6387(n1551 ,n0[83] ,n0[81]);
    nor g6388(n1550 ,n0[43] ,n0[41]);
    nor g6389(n1549 ,n0[67] ,n0[65]);
    or g6390(n1548 ,n1020 ,n0[56]);
    or g6391(n1547 ,n1020 ,n0[24]);
    nor g6392(n1546 ,n1269 ,n1024);
    or g6393(n1545 ,n1020 ,n0[88]);
    nor g6394(n1544 ,n1227 ,n0[18]);
    nor g6395(n1543 ,n1229 ,n0[122]);
    nor g6396(n1541 ,n1074 ,n0[113]);
    nor g6397(n1540 ,n0[115] ,n0[113]);
    nor g6398(n1538 ,n1235 ,n0[73]);
    nor g6399(n1537 ,n0[75] ,n0[73]);
    nor g6400(n1536 ,n0[35] ,n0[33]);
    nor g6401(n1534 ,n1080 ,n0[9]);
    nor g6402(n1533 ,n0[11] ,n0[9]);
    nor g6403(n1532 ,n0[107] ,n0[105]);
    nor g6404(n1530 ,n1232 ,n0[105]);
    nor g6405(n1528 ,n1072 ,n0[41]);
    or g6406(n1527 ,n0[2] ,n0[0]);
    nor g6407(n1525 ,n1250 ,n0[65]);
    nor g6408(n1524 ,n0[99] ,n0[97]);
    or g6409(n1523 ,n0[18] ,n0[16]);
    nor g6410(n1521 ,n1245 ,n0[97]);
    nor g6411(n1519 ,n1252 ,n0[33]);
    nor g6412(n1518 ,n1105 ,n1023);
    nor g6413(n1517 ,n1278 ,n1024);
    or g6414(n1516 ,n0[50] ,n0[48]);
    nor g6415(n1515 ,n1275 ,n1024);
    nor g6416(n1514 ,n0[17] ,n0[16]);
    or g6417(n1513 ,n3[2] ,n3[1]);
    not g6418(n1356 ,n7397);
    not g6419(n1355 ,n7454);
    not g6420(n1354 ,n7457);
    not g6421(n1353 ,n7405);
    not g6422(n1352 ,n7498);
    not g6423(n1351 ,n3[3]);
    not g6424(n1350 ,n7515);
    not g6425(n1349 ,n7518);
    not g6426(n1348 ,n7459);
    not g6427(n1347 ,n7422);
    not g6428(n1346 ,n7497);
    not g6429(n1345 ,n7514);
    not g6430(n1344 ,n7491);
    not g6431(n1343 ,n7501);
    not g6432(n1342 ,n7507);
    not g6433(n1341 ,n7450);
    not g6434(n1340 ,n7477);
    not g6435(n1339 ,n7469);
    not g6436(n1338 ,n7439);
    not g6437(n1337 ,n7475);
    not g6438(n1336 ,n7430);
    not g6439(n1335 ,n7499);
    not g6440(n1334 ,n7479);
    not g6441(n1333 ,n7629);
    not g6442(n1332 ,n7423);
    not g6443(n1331 ,n7474);
    not g6444(n1330 ,n7411);
    not g6445(n1329 ,n7473);
    not g6446(n1328 ,n7402);
    not g6447(n1327 ,n7447);
    not g6448(n1326 ,n7427);
    not g6449(n1325 ,n7485);
    not g6450(n1324 ,n7446);
    not g6451(n1323 ,n7522);
    not g6452(n1322 ,n7481);
    not g6453(n1321 ,n7445);
    not g6454(n1320 ,n7419);
    not g6455(n1319 ,n7494);
    not g6456(n1318 ,n7421);
    not g6457(n1317 ,n7437);
    not g6458(n1316 ,n7511);
    not g6459(n1315 ,n2[18]);
    not g6460(n1314 ,n2[26]);
    not g6461(n1313 ,n2[53]);
    not g6462(n1312 ,n2[1]);
    not g6463(n1311 ,n2[14]);
    not g6464(n1310 ,n1[90]);
    not g6465(n1309 ,n1[112]);
    not g6466(n1308 ,n1[78]);
    not g6467(n1307 ,n1[95]);
    not g6468(n1306 ,n0[39]);
    not g6469(n1305 ,n0[45]);
    not g6470(n1304 ,n0[61]);
    not g6471(n1303 ,n0[46]);
    not g6472(n1302 ,n0[47]);
    not g6473(n1301 ,n0[60]);
    not g6474(n1300 ,n1[61]);
    not g6475(n1299 ,n0[85]);
    not g6476(n1298 ,n1[85]);
    not g6477(n1297 ,n1[51]);
    not g6478(n1296 ,n1[33]);
    not g6479(n1295 ,n1[52]);
    not g6480(n1294 ,n1[53]);
    not g6481(n1293 ,n1[63]);
    not g6482(n1292 ,n1[41]);
    not g6483(n1291 ,n0[52]);
    not g6484(n1290 ,n1[62]);
    not g6485(n1289 ,n0[55]);
    not g6486(n1288 ,n1[116]);
    not g6487(n1287 ,n1[38]);
    not g6488(n1286 ,n1[45]);
    not g6489(n1285 ,n1[44]);
    not g6490(n1284 ,n0[6]);
    not g6491(n1283 ,n0[124]);
    not g6492(n1282 ,n0[5]);
    not g6493(n1281 ,n0[12]);
    not g6494(n1280 ,n0[103]);
    not g6495(n1279 ,n0[84]);
    not g6496(n1278 ,n0[109]);
    not g6497(n1277 ,n0[94]);
    not g6498(n1276 ,n0[7]);
    not g6499(n1275 ,n0[108]);
    not g6500(n1274 ,n0[22]);
    not g6501(n1273 ,n0[70]);
    not g6502(n1272 ,n0[93]);
    not g6503(n1271 ,n0[20]);
    not g6504(n1270 ,n0[116]);
    not g6505(n1269 ,n0[110]);
    not g6506(n1268 ,n0[95]);
    not g6507(n1267 ,n1[43]);
    not g6508(n1266 ,n0[50]);
    not g6509(n1265 ,n1[55]);
    not g6510(n1264 ,n0[41]);
    not g6511(n1263 ,n0[77]);
    not g6512(n1262 ,n0[51]);
    not g6513(n1261 ,n0[76]);
    not g6514(n1260 ,n0[58]);
    not g6515(n1259 ,n0[78]);
    not g6516(n1258 ,n1[50]);
    not g6517(n1257 ,n0[118]);
    not g6518(n1256 ,n0[65]);
    not g6519(n1255 ,n0[33]);
    not g6520(n1254 ,n0[79]);
    not g6521(n1253 ,n0[56]);
    not g6522(n1252 ,n0[32]);
    not g6523(n1251 ,n0[98]);
    not g6524(n1250 ,n0[64]);
    not g6525(n1249 ,n0[2]);
    not g6526(n1248 ,n0[67]);
    not g6527(n1247 ,n0[99]);
    not g6528(n1246 ,n0[14]);
    not g6529(n1245 ,n0[96]);
    not g6530(n1244 ,n0[90]);
    not g6531(n1243 ,n0[9]);
    not g6532(n1242 ,n0[18]);
    not g6533(n1241 ,n0[91]);
    not g6534(n1240 ,n0[81]);
    not g6535(n1239 ,n0[35]);
    not g6536(n1238 ,n0[80]);
    not g6537(n1237 ,n0[0]);
    not g6538(n1236 ,n0[24]);
    not g6539(n1235 ,n0[72]);
    not g6540(n1234 ,n0[75]);
    not g6541(n1233 ,n0[114]);
    not g6542(n1232 ,n0[104]);
    not g6543(n1231 ,n0[122]);
    not g6544(n1230 ,n0[115]);
    not g6545(n1229 ,n0[121]);
    not g6546(n1228 ,n0[10]);
    not g6547(n1227 ,n0[16]);
    not g6548(n1226 ,n0[120]);
    not g6549(n1225 ,n7399);
    not g6550(n1029 ,n1030);
    not g6551(n1027 ,n1029);
    not g6552(n1028 ,n1029);
    not g6553(n1026 ,n1029);
    not g6554(n1030 ,n7312);
    not g6555(n1025 ,n1024);
    buf g6556(n1024 ,n8);
    not g6557(n1023 ,n1022);
    not g6558(n1021 ,n1022);
    buf g6559(n1022 ,n8);
    not g6560(n1224 ,n7663);
    not g6561(n1223 ,n3[0]);
    not g6562(n1222 ,n7495);
    not g6563(n1221 ,n7490);
    not g6564(n1220 ,n7526);
    not g6565(n1219 ,n7425);
    not g6566(n1218 ,n7449);
    not g6567(n1217 ,n7470);
    not g6568(n1216 ,n7482);
    not g6569(n1215 ,n7431);
    not g6570(n1214 ,n7409);
    not g6571(n1213 ,n7525);
    not g6572(n1212 ,n7471);
    not g6573(n1211 ,n7493);
    not g6574(n1210 ,n7429);
    not g6575(n1209 ,n7413);
    not g6576(n1208 ,n7489);
    not g6577(n1207 ,n7523);
    not g6578(n1206 ,n7438);
    not g6579(n1205 ,n7414);
    not g6580(n1204 ,n7451);
    not g6581(n1203 ,n7509);
    not g6582(n1202 ,n7434);
    not g6583(n1201 ,n7417);
    not g6584(n1200 ,n7487);
    not g6585(n1199 ,n7502);
    not g6586(n1198 ,n7418);
    not g6587(n1197 ,n7513);
    not g6588(n1196 ,n7483);
    not g6589(n1195 ,n7462);
    not g6590(n1194 ,n7453);
    not g6591(n1193 ,n7442);
    not g6592(n1192 ,n7559);
    not g6593(n1191 ,n7465);
    not g6594(n1190 ,n7503);
    not g6595(n1189 ,n7486);
    not g6596(n1188 ,n7478);
    not g6597(n1187 ,n7441);
    not g6598(n1186 ,n7410);
    not g6599(n1185 ,n7517);
    not g6600(n1184 ,n7426);
    not g6601(n1183 ,n7406);
    not g6602(n1182 ,n7665);
    not g6603(n1181 ,n7467);
    not g6604(n1180 ,n7403);
    not g6605(n1179 ,n7433);
    not g6606(n1178 ,n7466);
    not g6607(n1177 ,n7458);
    not g6608(n1176 ,n7461);
    not g6609(n1175 ,n7505);
    not g6610(n1174 ,n7407);
    not g6611(n1173 ,n7463);
    not g6612(n1172 ,n7506);
    not g6613(n1171 ,n7435);
    not g6614(n1170 ,n3[1]);
    not g6615(n1169 ,n7510);
    not g6616(n1168 ,n7443);
    not g6617(n1167 ,n7455);
    not g6618(n1166 ,n7519);
    not g6619(n1165 ,n7415);
    not g6620(n1164 ,n7521);
    not g6621(n1163 ,n2[54]);
    not g6622(n1162 ,n3[2]);
    not g6623(n1161 ,n2[48]);
    not g6624(n1160 ,n2[55]);
    not g6625(n1159 ,n2[59]);
    not g6626(n1158 ,n1[64]);
    not g6627(n1157 ,n1[123]);
    not g6628(n1156 ,n1[94]);
    not g6629(n1155 ,n1[93]);
    not g6630(n1154 ,n1[65]);
    not g6631(n1153 ,n0[44]);
    not g6632(n1152 ,n0[38]);
    not g6633(n1151 ,n0[37]);
    not g6634(n1150 ,n0[54]);
    not g6635(n1149 ,n0[63]);
    not g6636(n1148 ,n0[62]);
    not g6637(n1147 ,n0[36]);
    not g6638(n1146 ,n1[35]);
    not g6639(n1145 ,n1[42]);
    not g6640(n1144 ,n1[119]);
    not g6641(n1143 ,n1[39]);
    not g6642(n1142 ,n1[32]);
    not g6643(n1141 ,n1[34]);
    not g6644(n1140 ,n1[60]);
    not g6645(n1139 ,n1[36]);
    not g6646(n1138 ,n0[53]);
    not g6647(n1137 ,n1[87]);
    not g6648(n1136 ,n1[59]);
    not g6649(n1135 ,n1[57]);
    not g6650(n1134 ,n1[37]);
    not g6651(n1133 ,n1[40]);
    not g6652(n1132 ,n1[58]);
    not g6653(n1131 ,n0[87]);
    not g6654(n1130 ,n1[48]);
    not g6655(n1129 ,n1[47]);
    not g6656(n1128 ,n1[86]);
    not g6657(n1127 ,n1[82]);
    not g6658(n1126 ,n0[86]);
    not g6659(n1125 ,n1[49]);
    not g6660(n1124 ,n0[28]);
    not g6661(n1123 ,n0[15]);
    not g6662(n1122 ,n1[54]);
    not g6663(n1121 ,n0[21]);
    not g6664(n1120 ,n0[92]);
    not g6665(n1119 ,n0[100]);
    not g6666(n1118 ,n0[127]);
    not g6667(n1117 ,n0[13]);
    not g6668(n1116 ,n0[125]);
    not g6669(n1115 ,n0[30]);
    not g6670(n1114 ,n0[126]);
    not g6671(n1113 ,n0[111]);
    not g6672(n1112 ,n0[23]);
    not g6673(n1111 ,n0[71]);
    not g6674(n1110 ,n0[68]);
    not g6675(n1109 ,n0[31]);
    not g6676(n1108 ,n0[29]);
    not g6677(n1107 ,n0[69]);
    not g6678(n1106 ,n0[117]);
    not g6679(n1105 ,n0[4]);
    not g6680(n1104 ,n0[59]);
    not g6681(n1103 ,n0[49]);
    not g6682(n1102 ,n1[56]);
    not g6683(n1101 ,n0[34]);
    not g6684(n1100 ,n0[102]);
    not g6685(n1099 ,n0[101]);
    not g6686(n1098 ,n0[57]);
    not g6687(n1097 ,n0[66]);
    not g6688(n1096 ,n0[119]);
    not g6689(n1095 ,n0[48]);
    not g6690(n1094 ,n0[42]);
    not g6691(n1093 ,n0[113]);
    not g6692(n1092 ,n0[19]);
    not g6693(n1091 ,n0[17]);
    not g6694(n1090 ,n0[105]);
    not g6695(n1089 ,n0[27]);
    not g6696(n1088 ,n0[1]);
    not g6697(n1087 ,n0[3]);
    not g6698(n1086 ,n0[88]);
    not g6699(n1085 ,n0[97]);
    not g6700(n1084 ,n0[26]);
    not g6701(n1083 ,n0[73]);
    not g6702(n1082 ,n0[43]);
    not g6703(n1081 ,n0[74]);
    not g6704(n1080 ,n0[8]);
    not g6705(n1079 ,n0[123]);
    not g6706(n1078 ,n0[83]);
    not g6707(n1077 ,n0[106]);
    not g6708(n1076 ,n0[25]);
    not g6709(n1075 ,n0[11]);
    not g6710(n1074 ,n0[112]);
    not g6711(n1073 ,n0[107]);
    not g6712(n1072 ,n0[40]);
    not g6713(n1071 ,n0[89]);
    not g6714(n1070 ,n0[82]);
    not g6715(n1069 ,n7311);
    not g6716(n1068 ,n7311);
    not g6717(n1067 ,n7311);
    not g6718(n1066 ,n7311);
    not g6719(n1020 ,n1065);
    not g6720(n1065 ,n7311);
    not g6721(n1064 ,n1063);
    not g6722(n1063 ,n7311);
    not g6723(n1018 ,n1062);
    not g6724(n1019 ,n1062);
    not g6725(n1017 ,n1062);
    not g6726(n1062 ,n7400);
    or g6727(n1016 ,n3998 ,n5087);
    xor g6728(n1015 ,n2436 ,n6499);
    xor g6729(n1014 ,n2439 ,n6496);
    xor g6730(n1013 ,n2484 ,n6495);
    xor g6731(n1012 ,n3197 ,n6293);
    xor g6732(n1011 ,n6081 ,n6567);
    xor g6733(n1010 ,n2438 ,n5977);
    xor g6734(n1009 ,n5578 ,n5977);
    xor g6735(n1008 ,n4318 ,n3408);
    xor g6736(n1007 ,n4309 ,n3406);
    xor g6737(n1006 ,n4308 ,n3401);
    xor g6738(n1005 ,n4307 ,n3398);
    or g6739(n7657 ,n983 ,n949);
    or g6740(n7660 ,n997 ,n954);
    or g6741(n7658 ,n993 ,n958);
    or g6742(n7655 ,n999 ,n965);
    or g6743(n7636 ,n1002 ,n971);
    or g6744(n7635 ,n1001 ,n969);
    or g6745(n7648 ,n998 ,n967);
    or g6746(n7634 ,n977 ,n968);
    or g6747(n7633 ,n996 ,n962);
    or g6748(n7654 ,n989 ,n959);
    or g6749(n7647 ,n995 ,n963);
    or g6750(n7632 ,n994 ,n964);
    or g6751(n7646 ,n988 ,n961);
    or g6752(n7631 ,n992 ,n966);
    or g6753(n7630 ,n1000 ,n960);
    or g6754(n7661 ,n1004 ,n972);
    or g6755(n7637 ,n973 ,n941);
    or g6756(n7645 ,n987 ,n957);
    or g6757(n7644 ,n985 ,n955);
    or g6758(n7643 ,n984 ,n952);
    or g6759(n7659 ,n974 ,n956);
    or g6760(n7652 ,n982 ,n950);
    or g6761(n7642 ,n981 ,n951);
    or g6762(n7641 ,n980 ,n948);
    or g6763(n7651 ,n979 ,n946);
    or g6764(n7640 ,n978 ,n947);
    or g6765(n7656 ,n975 ,n942);
    or g6766(n7650 ,n990 ,n943);
    or g6767(n7639 ,n976 ,n945);
    or g6768(n7638 ,n991 ,n944);
    or g6769(n7649 ,n1003 ,n970);
    or g6770(n7653 ,n986 ,n953);
    nor g6771(n1004 ,n891 ,n909);
    nor g6772(n1003 ,n877 ,n909);
    nor g6773(n1002 ,n924 ,n909);
    nor g6774(n1001 ,n935 ,n909);
    nor g6775(n1000 ,n881 ,n909);
    nor g6776(n999 ,n921 ,n909);
    nor g6777(n998 ,n925 ,n909);
    nor g6778(n997 ,n896 ,n909);
    nor g6779(n996 ,n939 ,n909);
    nor g6780(n995 ,n937 ,n909);
    nor g6781(n994 ,n886 ,n909);
    nor g6782(n993 ,n885 ,n909);
    nor g6783(n992 ,n887 ,n909);
    nor g6784(n991 ,n913 ,n909);
    nor g6785(n990 ,n911 ,n909);
    nor g6786(n989 ,n876 ,n909);
    nor g6787(n988 ,n917 ,n909);
    nor g6788(n987 ,n919 ,n909);
    nor g6789(n986 ,n914 ,n909);
    nor g6790(n985 ,n894 ,n909);
    nor g6791(n984 ,n908 ,n909);
    nor g6792(n983 ,n934 ,n909);
    nor g6793(n982 ,n899 ,n909);
    nor g6794(n981 ,n889 ,n909);
    nor g6795(n980 ,n931 ,n909);
    nor g6796(n979 ,n898 ,n909);
    nor g6797(n978 ,n927 ,n909);
    nor g6798(n977 ,n922 ,n909);
    nor g6799(n976 ,n883 ,n909);
    nor g6800(n975 ,n900 ,n909);
    nor g6801(n974 ,n888 ,n909);
    nor g6802(n973 ,n936 ,n909);
    nor g6803(n972 ,n932 ,n7400);
    nor g6804(n971 ,n938 ,n7400);
    nor g6805(n970 ,n929 ,n7400);
    nor g6806(n969 ,n930 ,n7400);
    nor g6807(n968 ,n928 ,n7400);
    nor g6808(n967 ,n923 ,n7400);
    nor g6809(n966 ,n915 ,n7400);
    nor g6810(n965 ,n920 ,n7400);
    nor g6811(n964 ,n905 ,n7400);
    nor g6812(n963 ,n901 ,n7400);
    nor g6813(n962 ,n916 ,n7400);
    nor g6814(n961 ,n879 ,n7400);
    nor g6815(n960 ,n892 ,n7400);
    nor g6816(n959 ,n897 ,n7400);
    nor g6817(n958 ,n895 ,n7400);
    nor g6818(n957 ,n884 ,n7400);
    nor g6819(n956 ,n933 ,n7400);
    nor g6820(n955 ,n878 ,n7400);
    nor g6821(n954 ,n910 ,n7400);
    nor g6822(n953 ,n893 ,n7400);
    nor g6823(n952 ,n882 ,n7400);
    nor g6824(n951 ,n903 ,n7400);
    nor g6825(n950 ,n902 ,n7400);
    nor g6826(n949 ,n926 ,n7400);
    nor g6827(n948 ,n940 ,n7400);
    nor g6828(n947 ,n890 ,n7400);
    nor g6829(n946 ,n918 ,n7400);
    nor g6830(n945 ,n907 ,n7400);
    nor g6831(n944 ,n912 ,n7400);
    nor g6832(n943 ,n880 ,n7400);
    nor g6833(n942 ,n906 ,n7400);
    nor g6834(n941 ,n904 ,n7400);
    not g6835(n940 ,n0[75]);
    not g6836(n939 ,n1[3]);
    not g6837(n938 ,n0[70]);
    not g6838(n937 ,n1[17]);
    not g6839(n936 ,n1[7]);
    not g6840(n935 ,n1[5]);
    not g6841(n934 ,n1[27]);
    not g6842(n933 ,n0[93]);
    not g6843(n932 ,n0[95]);
    not g6844(n931 ,n1[11]);
    not g6845(n930 ,n0[69]);
    not g6846(n929 ,n0[83]);
    not g6847(n928 ,n0[68]);
    not g6848(n927 ,n1[10]);
    not g6849(n926 ,n0[91]);
    not g6850(n925 ,n1[18]);
    not g6851(n924 ,n1[6]);
    not g6852(n923 ,n0[82]);
    not g6853(n922 ,n1[4]);
    not g6854(n921 ,n1[25]);
    not g6855(n920 ,n0[89]);
    not g6856(n919 ,n1[15]);
    not g6857(n918 ,n0[85]);
    not g6858(n917 ,n1[16]);
    not g6859(n916 ,n0[67]);
    not g6860(n915 ,n0[65]);
    not g6861(n914 ,n1[23]);
    not g6862(n913 ,n1[8]);
    not g6863(n912 ,n0[72]);
    not g6864(n911 ,n1[20]);
    not g6865(n910 ,n0[94]);
    not g6866(n909 ,n7662);
    not g6867(n908 ,n1[13]);
    not g6868(n907 ,n0[73]);
    not g6869(n906 ,n0[90]);
    not g6870(n905 ,n0[66]);
    not g6871(n904 ,n0[71]);
    not g6872(n903 ,n0[76]);
    not g6873(n902 ,n0[86]);
    not g6874(n901 ,n0[81]);
    not g6875(n900 ,n1[26]);
    not g6876(n899 ,n1[22]);
    not g6877(n898 ,n1[21]);
    not g6878(n897 ,n0[88]);
    not g6879(n896 ,n1[30]);
    not g6880(n895 ,n0[92]);
    not g6881(n894 ,n1[14]);
    not g6882(n893 ,n0[87]);
    not g6883(n892 ,n0[64]);
    not g6884(n891 ,n1[31]);
    not g6885(n890 ,n0[74]);
    not g6886(n889 ,n1[12]);
    not g6887(n888 ,n1[29]);
    not g6888(n887 ,n1[1]);
    not g6889(n886 ,n1[2]);
    not g6890(n885 ,n1[28]);
    not g6891(n884 ,n0[79]);
    not g6892(n883 ,n1[9]);
    not g6893(n882 ,n0[77]);
    not g6894(n881 ,n1[0]);
    not g6895(n880 ,n0[84]);
    not g6896(n879 ,n0[80]);
    not g6897(n878 ,n0[78]);
    not g6898(n877 ,n1[19]);
    not g6899(n876 ,n1[24]);
    xor g6900(n7629 ,n148 ,n227);
    nor g6901(n227 ,n125 ,n226);
    xor g6902(n7525 ,n147 ,n225);
    nor g6903(n226 ,n78 ,n225);
    nor g6904(n225 ,n106 ,n224);
    xor g6905(n7521 ,n146 ,n223);
    nor g6906(n224 ,n88 ,n223);
    nor g6907(n223 ,n109 ,n222);
    xor g6908(n7517 ,n145 ,n221);
    nor g6909(n222 ,n80 ,n221);
    nor g6910(n221 ,n112 ,n220);
    xor g6911(n7513 ,n144 ,n219);
    nor g6912(n220 ,n79 ,n219);
    nor g6913(n219 ,n131 ,n218);
    xor g6914(n7509 ,n143 ,n217);
    nor g6915(n218 ,n103 ,n217);
    nor g6916(n217 ,n130 ,n216);
    xor g6917(n7505 ,n142 ,n215);
    nor g6918(n216 ,n86 ,n215);
    nor g6919(n215 ,n113 ,n214);
    xor g6920(n7501 ,n141 ,n213);
    nor g6921(n214 ,n81 ,n213);
    nor g6922(n213 ,n116 ,n212);
    xor g6923(n7497 ,n140 ,n211);
    nor g6924(n212 ,n104 ,n211);
    nor g6925(n211 ,n110 ,n210);
    xor g6926(n7493 ,n139 ,n209);
    nor g6927(n210 ,n90 ,n209);
    nor g6928(n209 ,n118 ,n208);
    xor g6929(n7489 ,n138 ,n207);
    nor g6930(n208 ,n99 ,n207);
    nor g6931(n207 ,n107 ,n206);
    xor g6932(n7485 ,n137 ,n205);
    nor g6933(n206 ,n94 ,n205);
    nor g6934(n205 ,n127 ,n204);
    xor g6935(n7481 ,n167 ,n203);
    nor g6936(n204 ,n102 ,n203);
    nor g6937(n203 ,n122 ,n202);
    xor g6938(n7477 ,n166 ,n201);
    nor g6939(n202 ,n95 ,n201);
    nor g6940(n201 ,n128 ,n200);
    xor g6941(n7473 ,n165 ,n199);
    nor g6942(n200 ,n83 ,n199);
    nor g6943(n199 ,n119 ,n198);
    xor g6944(n7469 ,n164 ,n197);
    nor g6945(n198 ,n82 ,n197);
    nor g6946(n197 ,n117 ,n196);
    xor g6947(n7465 ,n163 ,n195);
    nor g6948(n196 ,n85 ,n195);
    nor g6949(n195 ,n114 ,n194);
    xor g6950(n7461 ,n162 ,n193);
    nor g6951(n194 ,n100 ,n193);
    nor g6952(n193 ,n111 ,n192);
    xor g6953(n7457 ,n161 ,n191);
    nor g6954(n192 ,n87 ,n191);
    nor g6955(n191 ,n108 ,n190);
    xor g6956(n7453 ,n160 ,n189);
    nor g6957(n190 ,n89 ,n189);
    nor g6958(n189 ,n105 ,n188);
    xor g6959(n7449 ,n159 ,n187);
    nor g6960(n188 ,n97 ,n187);
    nor g6961(n187 ,n133 ,n186);
    xor g6962(n7445 ,n158 ,n185);
    nor g6963(n186 ,n93 ,n185);
    nor g6964(n185 ,n129 ,n184);
    xor g6965(n7441 ,n157 ,n183);
    nor g6966(n184 ,n75 ,n183);
    nor g6967(n183 ,n126 ,n182);
    xor g6968(n7437 ,n156 ,n181);
    nor g6969(n182 ,n98 ,n181);
    nor g6970(n181 ,n124 ,n180);
    xor g6971(n7433 ,n155 ,n179);
    nor g6972(n180 ,n74 ,n179);
    nor g6973(n179 ,n123 ,n178);
    xor g6974(n7429 ,n154 ,n177);
    nor g6975(n178 ,n96 ,n177);
    nor g6976(n177 ,n134 ,n176);
    xor g6977(n7425 ,n153 ,n175);
    nor g6978(n176 ,n91 ,n175);
    nor g6979(n175 ,n121 ,n174);
    xor g6980(n7421 ,n152 ,n173);
    nor g6981(n174 ,n77 ,n173);
    nor g6982(n173 ,n132 ,n172);
    xor g6983(n7417 ,n151 ,n171);
    nor g6984(n172 ,n76 ,n171);
    nor g6985(n171 ,n120 ,n170);
    xor g6986(n7413 ,n150 ,n169);
    nor g6987(n170 ,n92 ,n169);
    xnor g6988(n7409 ,n149 ,n135);
    nor g6989(n169 ,n115 ,n168);
    nor g6990(n7405 ,n135 ,n101);
    nor g6991(n168 ,n136 ,n84);
    xnor g6992(n167 ,n0[19] ,n7649);
    xnor g6993(n166 ,n0[18] ,n7648);
    xnor g6994(n165 ,n0[17] ,n7647);
    xnor g6995(n164 ,n0[16] ,n7646);
    xnor g6996(n163 ,n0[15] ,n7645);
    xnor g6997(n162 ,n0[14] ,n7644);
    xnor g6998(n161 ,n0[13] ,n7643);
    xnor g6999(n160 ,n0[12] ,n7642);
    xnor g7000(n159 ,n0[11] ,n7641);
    xnor g7001(n158 ,n0[10] ,n7640);
    xnor g7002(n157 ,n0[9] ,n7639);
    xnor g7003(n156 ,n0[8] ,n7638);
    xnor g7004(n155 ,n0[7] ,n7637);
    xnor g7005(n154 ,n0[6] ,n7636);
    xnor g7006(n153 ,n0[5] ,n7635);
    xnor g7007(n152 ,n0[4] ,n7634);
    xnor g7008(n151 ,n0[3] ,n7633);
    xnor g7009(n150 ,n0[2] ,n7632);
    xnor g7010(n149 ,n0[1] ,n7631);
    xnor g7011(n148 ,n7661 ,n0[31]);
    xnor g7012(n147 ,n0[30] ,n7660);
    xnor g7013(n146 ,n0[29] ,n7659);
    xnor g7014(n145 ,n0[28] ,n7658);
    xnor g7015(n144 ,n0[27] ,n7657);
    xnor g7016(n143 ,n0[26] ,n7656);
    xnor g7017(n142 ,n0[25] ,n7655);
    xnor g7018(n141 ,n0[24] ,n7654);
    xnor g7019(n140 ,n0[23] ,n7653);
    xnor g7020(n139 ,n0[22] ,n7652);
    xnor g7021(n138 ,n0[21] ,n7651);
    xnor g7022(n137 ,n0[20] ,n7650);
    not g7023(n136 ,n135);
    nor g7024(n134 ,n42 ,n22);
    nor g7025(n133 ,n64 ,n68);
    nor g7026(n132 ,n35 ,n33);
    nor g7027(n131 ,n15 ,n45);
    nor g7028(n130 ,n38 ,n26);
    nor g7029(n129 ,n13 ,n52);
    nor g7030(n128 ,n56 ,n23);
    nor g7031(n127 ,n30 ,n70);
    nor g7032(n126 ,n46 ,n16);
    nor g7033(n125 ,n53 ,n69);
    nor g7034(n124 ,n34 ,n28);
    nor g7035(n123 ,n27 ,n55);
    nor g7036(n122 ,n39 ,n57);
    nor g7037(n121 ,n37 ,n44);
    nor g7038(n120 ,n24 ,n60);
    nor g7039(n119 ,n19 ,n51);
    nor g7040(n118 ,n58 ,n67);
    nor g7041(n117 ,n66 ,n72);
    nor g7042(n116 ,n54 ,n31);
    nor g7043(n115 ,n32 ,n71);
    nor g7044(n114 ,n65 ,n36);
    nor g7045(n113 ,n62 ,n40);
    nor g7046(n112 ,n50 ,n25);
    nor g7047(n111 ,n29 ,n47);
    nor g7048(n110 ,n63 ,n61);
    nor g7049(n109 ,n12 ,n20);
    nor g7050(n108 ,n21 ,n18);
    nor g7051(n107 ,n17 ,n48);
    nor g7052(n106 ,n49 ,n59);
    nor g7053(n105 ,n14 ,n41);
    nor g7054(n135 ,n73 ,n43);
    nor g7055(n104 ,n7653 ,n0[23]);
    nor g7056(n103 ,n7656 ,n0[26]);
    nor g7057(n102 ,n7649 ,n0[19]);
    nor g7058(n101 ,n7630 ,n0[0]);
    nor g7059(n100 ,n7644 ,n0[14]);
    nor g7060(n99 ,n7651 ,n0[21]);
    nor g7061(n98 ,n7638 ,n0[8]);
    nor g7062(n97 ,n7641 ,n0[11]);
    nor g7063(n96 ,n7636 ,n0[6]);
    nor g7064(n95 ,n7648 ,n0[18]);
    nor g7065(n94 ,n7650 ,n0[20]);
    nor g7066(n93 ,n7640 ,n0[10]);
    nor g7067(n92 ,n7632 ,n0[2]);
    nor g7068(n91 ,n7635 ,n0[5]);
    nor g7069(n90 ,n7652 ,n0[22]);
    nor g7070(n89 ,n7642 ,n0[12]);
    nor g7071(n88 ,n7659 ,n0[29]);
    nor g7072(n87 ,n7643 ,n0[13]);
    nor g7073(n86 ,n7655 ,n0[25]);
    nor g7074(n85 ,n7645 ,n0[15]);
    nor g7075(n84 ,n7631 ,n0[1]);
    nor g7076(n83 ,n7647 ,n0[17]);
    nor g7077(n82 ,n7646 ,n0[16]);
    nor g7078(n81 ,n7654 ,n0[24]);
    nor g7079(n80 ,n7658 ,n0[28]);
    nor g7080(n79 ,n7657 ,n0[27]);
    nor g7081(n78 ,n7660 ,n0[30]);
    nor g7082(n77 ,n7634 ,n0[4]);
    nor g7083(n76 ,n7633 ,n0[3]);
    nor g7084(n75 ,n7639 ,n0[9]);
    nor g7085(n74 ,n7637 ,n0[7]);
    not g7086(n73 ,n7630);
    not g7087(n72 ,n0[15]);
    not g7088(n71 ,n0[1]);
    not g7089(n70 ,n0[19]);
    not g7090(n69 ,n0[30]);
    not g7091(n68 ,n0[10]);
    not g7092(n67 ,n0[21]);
    not g7093(n66 ,n7645);
    not g7094(n65 ,n7644);
    not g7095(n64 ,n7640);
    not g7096(n63 ,n7652);
    not g7097(n62 ,n7654);
    not g7098(n61 ,n0[22]);
    not g7099(n60 ,n0[2]);
    not g7100(n59 ,n0[29]);
    not g7101(n58 ,n7651);
    not g7102(n57 ,n0[18]);
    not g7103(n56 ,n7647);
    not g7104(n55 ,n0[6]);
    not g7105(n54 ,n7653);
    not g7106(n53 ,n7660);
    not g7107(n52 ,n0[9]);
    not g7108(n51 ,n0[16]);
    not g7109(n50 ,n7657);
    not g7110(n49 ,n7659);
    not g7111(n48 ,n0[20]);
    not g7112(n47 ,n0[13]);
    not g7113(n46 ,n7638);
    not g7114(n45 ,n0[26]);
    not g7115(n44 ,n0[4]);
    not g7116(n43 ,n0[0]);
    not g7117(n42 ,n7635);
    not g7118(n41 ,n0[11]);
    not g7119(n40 ,n0[24]);
    not g7120(n39 ,n7648);
    not g7121(n38 ,n7655);
    not g7122(n37 ,n7634);
    not g7123(n36 ,n0[14]);
    not g7124(n35 ,n7633);
    not g7125(n34 ,n7637);
    not g7126(n33 ,n0[3]);
    not g7127(n32 ,n7631);
    not g7128(n31 ,n0[23]);
    not g7129(n30 ,n7649);
    not g7130(n29 ,n7643);
    not g7131(n28 ,n0[7]);
    not g7132(n27 ,n7636);
    not g7133(n26 ,n0[25]);
    not g7134(n25 ,n0[27]);
    not g7135(n24 ,n7632);
    not g7136(n23 ,n0[17]);
    not g7137(n22 ,n0[5]);
    not g7138(n21 ,n7642);
    not g7139(n20 ,n0[28]);
    not g7140(n19 ,n7646);
    not g7141(n18 ,n0[12]);
    not g7142(n17 ,n7650);
    not g7143(n16 ,n0[8]);
    not g7144(n15 ,n7656);
    not g7145(n14 ,n7641);
    not g7146(n13 ,n7639);
    not g7147(n12 ,n7658);
    xor g7148(n7628 ,n364 ,n443);
    nor g7149(n443 ,n341 ,n442);
    xor g7150(n7524 ,n363 ,n441);
    nor g7151(n442 ,n294 ,n441);
    nor g7152(n441 ,n322 ,n440);
    xor g7153(n7520 ,n362 ,n439);
    nor g7154(n440 ,n304 ,n439);
    nor g7155(n439 ,n325 ,n438);
    xor g7156(n7516 ,n361 ,n437);
    nor g7157(n438 ,n296 ,n437);
    nor g7158(n437 ,n328 ,n436);
    xor g7159(n7512 ,n360 ,n435);
    nor g7160(n436 ,n295 ,n435);
    nor g7161(n435 ,n347 ,n434);
    xor g7162(n7508 ,n359 ,n433);
    nor g7163(n434 ,n319 ,n433);
    nor g7164(n433 ,n346 ,n432);
    xor g7165(n7504 ,n358 ,n431);
    nor g7166(n432 ,n302 ,n431);
    nor g7167(n431 ,n329 ,n430);
    xor g7168(n7500 ,n357 ,n429);
    nor g7169(n430 ,n297 ,n429);
    nor g7170(n429 ,n332 ,n428);
    xor g7171(n7496 ,n356 ,n427);
    nor g7172(n428 ,n320 ,n427);
    nor g7173(n427 ,n326 ,n426);
    xor g7174(n7492 ,n355 ,n425);
    nor g7175(n426 ,n306 ,n425);
    nor g7176(n425 ,n334 ,n424);
    xor g7177(n7488 ,n354 ,n423);
    nor g7178(n424 ,n315 ,n423);
    nor g7179(n423 ,n323 ,n422);
    xor g7180(n7484 ,n353 ,n421);
    nor g7181(n422 ,n310 ,n421);
    nor g7182(n421 ,n343 ,n420);
    xor g7183(n7480 ,n383 ,n419);
    nor g7184(n420 ,n318 ,n419);
    nor g7185(n419 ,n338 ,n418);
    xor g7186(n7476 ,n382 ,n417);
    nor g7187(n418 ,n311 ,n417);
    nor g7188(n417 ,n344 ,n416);
    xor g7189(n7472 ,n381 ,n415);
    nor g7190(n416 ,n299 ,n415);
    nor g7191(n415 ,n335 ,n414);
    xor g7192(n7468 ,n380 ,n413);
    nor g7193(n414 ,n298 ,n413);
    nor g7194(n413 ,n333 ,n412);
    xor g7195(n7464 ,n379 ,n411);
    nor g7196(n412 ,n301 ,n411);
    nor g7197(n411 ,n330 ,n410);
    xor g7198(n7460 ,n378 ,n409);
    nor g7199(n410 ,n316 ,n409);
    nor g7200(n409 ,n327 ,n408);
    xor g7201(n7456 ,n377 ,n407);
    nor g7202(n408 ,n303 ,n407);
    nor g7203(n407 ,n324 ,n406);
    xor g7204(n7452 ,n376 ,n405);
    nor g7205(n406 ,n305 ,n405);
    nor g7206(n405 ,n321 ,n404);
    xor g7207(n7448 ,n375 ,n403);
    nor g7208(n404 ,n313 ,n403);
    nor g7209(n403 ,n349 ,n402);
    xor g7210(n7444 ,n374 ,n401);
    nor g7211(n402 ,n309 ,n401);
    nor g7212(n401 ,n345 ,n400);
    xor g7213(n7440 ,n373 ,n399);
    nor g7214(n400 ,n291 ,n399);
    nor g7215(n399 ,n342 ,n398);
    xor g7216(n7436 ,n372 ,n397);
    nor g7217(n398 ,n314 ,n397);
    nor g7218(n397 ,n340 ,n396);
    xor g7219(n7432 ,n371 ,n395);
    nor g7220(n396 ,n290 ,n395);
    nor g7221(n395 ,n339 ,n394);
    xor g7222(n7428 ,n370 ,n393);
    nor g7223(n394 ,n312 ,n393);
    nor g7224(n393 ,n350 ,n392);
    xor g7225(n7424 ,n369 ,n391);
    nor g7226(n392 ,n307 ,n391);
    nor g7227(n391 ,n337 ,n390);
    xor g7228(n7420 ,n368 ,n389);
    nor g7229(n390 ,n293 ,n389);
    nor g7230(n389 ,n348 ,n388);
    xor g7231(n7416 ,n367 ,n387);
    nor g7232(n388 ,n292 ,n387);
    nor g7233(n387 ,n336 ,n386);
    xor g7234(n7412 ,n366 ,n385);
    nor g7235(n386 ,n308 ,n385);
    xnor g7236(n7408 ,n365 ,n351);
    nor g7237(n385 ,n331 ,n384);
    nor g7238(n7404 ,n351 ,n317);
    nor g7239(n384 ,n352 ,n300);
    xnor g7240(n383 ,n1[51] ,n0[51]);
    xnor g7241(n382 ,n1[50] ,n0[50]);
    xnor g7242(n381 ,n1[49] ,n0[49]);
    xnor g7243(n380 ,n1[48] ,n0[48]);
    xnor g7244(n379 ,n1[47] ,n0[47]);
    xnor g7245(n378 ,n1[46] ,n0[46]);
    xnor g7246(n377 ,n1[45] ,n0[45]);
    xnor g7247(n376 ,n1[44] ,n0[44]);
    xnor g7248(n375 ,n1[43] ,n0[43]);
    xnor g7249(n374 ,n1[42] ,n0[42]);
    xnor g7250(n373 ,n1[41] ,n0[41]);
    xnor g7251(n372 ,n1[40] ,n0[40]);
    xnor g7252(n371 ,n1[39] ,n0[39]);
    xnor g7253(n370 ,n1[38] ,n0[38]);
    xnor g7254(n369 ,n1[37] ,n0[37]);
    xnor g7255(n368 ,n1[36] ,n0[36]);
    xnor g7256(n367 ,n1[35] ,n0[35]);
    xnor g7257(n366 ,n1[34] ,n0[34]);
    xnor g7258(n365 ,n1[33] ,n0[33]);
    xnor g7259(n364 ,n0[63] ,n1[63]);
    xnor g7260(n363 ,n1[62] ,n0[62]);
    xnor g7261(n362 ,n1[61] ,n0[61]);
    xnor g7262(n361 ,n1[60] ,n0[60]);
    xnor g7263(n360 ,n1[59] ,n0[59]);
    xnor g7264(n359 ,n1[58] ,n0[58]);
    xnor g7265(n358 ,n1[57] ,n0[57]);
    xnor g7266(n357 ,n1[56] ,n0[56]);
    xnor g7267(n356 ,n1[55] ,n0[55]);
    xnor g7268(n355 ,n1[54] ,n0[54]);
    xnor g7269(n354 ,n1[53] ,n0[53]);
    xnor g7270(n353 ,n1[52] ,n0[52]);
    not g7271(n352 ,n351);
    nor g7272(n350 ,n258 ,n238);
    nor g7273(n349 ,n280 ,n284);
    nor g7274(n348 ,n251 ,n249);
    nor g7275(n347 ,n231 ,n261);
    nor g7276(n346 ,n254 ,n242);
    nor g7277(n345 ,n229 ,n268);
    nor g7278(n344 ,n272 ,n239);
    nor g7279(n343 ,n246 ,n286);
    nor g7280(n342 ,n262 ,n232);
    nor g7281(n341 ,n269 ,n285);
    nor g7282(n340 ,n250 ,n244);
    nor g7283(n339 ,n243 ,n271);
    nor g7284(n338 ,n255 ,n273);
    nor g7285(n337 ,n253 ,n260);
    nor g7286(n336 ,n240 ,n276);
    nor g7287(n335 ,n235 ,n267);
    nor g7288(n334 ,n274 ,n283);
    nor g7289(n333 ,n282 ,n288);
    nor g7290(n332 ,n270 ,n247);
    nor g7291(n331 ,n248 ,n287);
    nor g7292(n330 ,n281 ,n252);
    nor g7293(n329 ,n278 ,n256);
    nor g7294(n328 ,n266 ,n241);
    nor g7295(n327 ,n245 ,n263);
    nor g7296(n326 ,n279 ,n277);
    nor g7297(n325 ,n228 ,n236);
    nor g7298(n324 ,n237 ,n234);
    nor g7299(n323 ,n233 ,n264);
    nor g7300(n322 ,n265 ,n275);
    nor g7301(n321 ,n230 ,n257);
    nor g7302(n351 ,n289 ,n259);
    nor g7303(n320 ,n0[55] ,n1[55]);
    nor g7304(n319 ,n0[58] ,n1[58]);
    nor g7305(n318 ,n0[51] ,n1[51]);
    nor g7306(n317 ,n0[32] ,n1[32]);
    nor g7307(n316 ,n0[46] ,n1[46]);
    nor g7308(n315 ,n0[53] ,n1[53]);
    nor g7309(n314 ,n0[40] ,n1[40]);
    nor g7310(n313 ,n0[43] ,n1[43]);
    nor g7311(n312 ,n0[38] ,n1[38]);
    nor g7312(n311 ,n0[50] ,n1[50]);
    nor g7313(n310 ,n0[52] ,n1[52]);
    nor g7314(n309 ,n0[42] ,n1[42]);
    nor g7315(n308 ,n0[34] ,n1[34]);
    nor g7316(n307 ,n0[37] ,n1[37]);
    nor g7317(n306 ,n0[54] ,n1[54]);
    nor g7318(n305 ,n0[44] ,n1[44]);
    nor g7319(n304 ,n0[61] ,n1[61]);
    nor g7320(n303 ,n0[45] ,n1[45]);
    nor g7321(n302 ,n0[57] ,n1[57]);
    nor g7322(n301 ,n0[47] ,n1[47]);
    nor g7323(n300 ,n0[33] ,n1[33]);
    nor g7324(n299 ,n0[49] ,n1[49]);
    nor g7325(n298 ,n0[48] ,n1[48]);
    nor g7326(n297 ,n0[56] ,n1[56]);
    nor g7327(n296 ,n0[60] ,n1[60]);
    nor g7328(n295 ,n0[59] ,n1[59]);
    nor g7329(n294 ,n0[62] ,n1[62]);
    nor g7330(n293 ,n0[36] ,n1[36]);
    nor g7331(n292 ,n0[35] ,n1[35]);
    nor g7332(n291 ,n0[41] ,n1[41]);
    nor g7333(n290 ,n0[39] ,n1[39]);
    not g7334(n289 ,n0[32]);
    not g7335(n288 ,n1[47]);
    not g7336(n287 ,n1[33]);
    not g7337(n286 ,n1[51]);
    not g7338(n285 ,n1[62]);
    not g7339(n284 ,n1[42]);
    not g7340(n283 ,n1[53]);
    not g7341(n282 ,n0[47]);
    not g7342(n281 ,n0[46]);
    not g7343(n280 ,n0[42]);
    not g7344(n279 ,n0[54]);
    not g7345(n278 ,n0[56]);
    not g7346(n277 ,n1[54]);
    not g7347(n276 ,n1[34]);
    not g7348(n275 ,n1[61]);
    not g7349(n274 ,n0[53]);
    not g7350(n273 ,n1[50]);
    not g7351(n272 ,n0[49]);
    not g7352(n271 ,n1[38]);
    not g7353(n270 ,n0[55]);
    not g7354(n269 ,n0[62]);
    not g7355(n268 ,n1[41]);
    not g7356(n267 ,n1[48]);
    not g7357(n266 ,n0[59]);
    not g7358(n265 ,n0[61]);
    not g7359(n264 ,n1[52]);
    not g7360(n263 ,n1[45]);
    not g7361(n262 ,n0[40]);
    not g7362(n261 ,n1[58]);
    not g7363(n260 ,n1[36]);
    not g7364(n259 ,n1[32]);
    not g7365(n258 ,n0[37]);
    not g7366(n257 ,n1[43]);
    not g7367(n256 ,n1[56]);
    not g7368(n255 ,n0[50]);
    not g7369(n254 ,n0[57]);
    not g7370(n253 ,n0[36]);
    not g7371(n252 ,n1[46]);
    not g7372(n251 ,n0[35]);
    not g7373(n250 ,n0[39]);
    not g7374(n249 ,n1[35]);
    not g7375(n248 ,n0[33]);
    not g7376(n247 ,n1[55]);
    not g7377(n246 ,n0[51]);
    not g7378(n245 ,n0[45]);
    not g7379(n244 ,n1[39]);
    not g7380(n243 ,n0[38]);
    not g7381(n242 ,n1[57]);
    not g7382(n241 ,n1[59]);
    not g7383(n240 ,n0[34]);
    not g7384(n239 ,n1[49]);
    not g7385(n238 ,n1[37]);
    not g7386(n237 ,n0[44]);
    not g7387(n236 ,n1[60]);
    not g7388(n235 ,n0[48]);
    not g7389(n234 ,n1[44]);
    not g7390(n233 ,n0[52]);
    not g7391(n232 ,n1[40]);
    not g7392(n231 ,n0[58]);
    not g7393(n230 ,n0[43]);
    not g7394(n229 ,n0[41]);
    not g7395(n228 ,n0[60]);
    xor g7396(n7559 ,n580 ,n659);
    nor g7397(n659 ,n557 ,n658);
    xor g7398(n7523 ,n579 ,n657);
    nor g7399(n658 ,n510 ,n657);
    nor g7400(n657 ,n538 ,n656);
    xor g7401(n7519 ,n578 ,n655);
    nor g7402(n656 ,n520 ,n655);
    nor g7403(n655 ,n541 ,n654);
    xor g7404(n7515 ,n577 ,n653);
    nor g7405(n654 ,n512 ,n653);
    nor g7406(n653 ,n544 ,n652);
    xor g7407(n7511 ,n576 ,n651);
    nor g7408(n652 ,n511 ,n651);
    nor g7409(n651 ,n563 ,n650);
    xor g7410(n7507 ,n575 ,n649);
    nor g7411(n650 ,n535 ,n649);
    nor g7412(n649 ,n562 ,n648);
    xor g7413(n7503 ,n574 ,n647);
    nor g7414(n648 ,n518 ,n647);
    nor g7415(n647 ,n545 ,n646);
    xor g7416(n7499 ,n573 ,n645);
    nor g7417(n646 ,n513 ,n645);
    nor g7418(n645 ,n548 ,n644);
    xor g7419(n7495 ,n572 ,n643);
    nor g7420(n644 ,n536 ,n643);
    nor g7421(n643 ,n542 ,n642);
    xor g7422(n7491 ,n571 ,n641);
    nor g7423(n642 ,n522 ,n641);
    nor g7424(n641 ,n550 ,n640);
    xor g7425(n7487 ,n570 ,n639);
    nor g7426(n640 ,n531 ,n639);
    nor g7427(n639 ,n539 ,n638);
    xor g7428(n7483 ,n569 ,n637);
    nor g7429(n638 ,n526 ,n637);
    nor g7430(n637 ,n559 ,n636);
    xor g7431(n7479 ,n599 ,n635);
    nor g7432(n636 ,n534 ,n635);
    nor g7433(n635 ,n554 ,n634);
    xor g7434(n7475 ,n598 ,n633);
    nor g7435(n634 ,n527 ,n633);
    nor g7436(n633 ,n560 ,n632);
    xor g7437(n7471 ,n597 ,n631);
    nor g7438(n632 ,n515 ,n631);
    nor g7439(n631 ,n551 ,n630);
    xor g7440(n7467 ,n596 ,n629);
    nor g7441(n630 ,n514 ,n629);
    nor g7442(n629 ,n549 ,n628);
    xor g7443(n7463 ,n595 ,n627);
    nor g7444(n628 ,n517 ,n627);
    nor g7445(n627 ,n546 ,n626);
    xor g7446(n7459 ,n594 ,n625);
    nor g7447(n626 ,n532 ,n625);
    nor g7448(n625 ,n543 ,n624);
    xor g7449(n7455 ,n593 ,n623);
    nor g7450(n624 ,n519 ,n623);
    nor g7451(n623 ,n540 ,n622);
    xor g7452(n7451 ,n592 ,n621);
    nor g7453(n622 ,n521 ,n621);
    nor g7454(n621 ,n537 ,n620);
    xor g7455(n7447 ,n591 ,n619);
    nor g7456(n620 ,n529 ,n619);
    nor g7457(n619 ,n565 ,n618);
    xor g7458(n7443 ,n590 ,n617);
    nor g7459(n618 ,n525 ,n617);
    nor g7460(n617 ,n561 ,n616);
    xor g7461(n7439 ,n589 ,n615);
    nor g7462(n616 ,n507 ,n615);
    nor g7463(n615 ,n558 ,n614);
    xor g7464(n7435 ,n588 ,n613);
    nor g7465(n614 ,n530 ,n613);
    nor g7466(n613 ,n556 ,n612);
    xor g7467(n7431 ,n587 ,n611);
    nor g7468(n612 ,n506 ,n611);
    nor g7469(n611 ,n555 ,n610);
    xor g7470(n7427 ,n586 ,n609);
    nor g7471(n610 ,n528 ,n609);
    nor g7472(n609 ,n566 ,n608);
    xor g7473(n7423 ,n585 ,n607);
    nor g7474(n608 ,n523 ,n607);
    nor g7475(n607 ,n553 ,n606);
    xor g7476(n7419 ,n584 ,n605);
    nor g7477(n606 ,n509 ,n605);
    nor g7478(n605 ,n564 ,n604);
    xor g7479(n7415 ,n583 ,n603);
    nor g7480(n604 ,n508 ,n603);
    nor g7481(n603 ,n552 ,n602);
    xor g7482(n7411 ,n582 ,n601);
    nor g7483(n602 ,n524 ,n601);
    xnor g7484(n7407 ,n581 ,n567);
    nor g7485(n601 ,n547 ,n600);
    nor g7486(n7403 ,n567 ,n533);
    nor g7487(n600 ,n568 ,n516);
    xnor g7488(n599 ,n7579 ,n7611);
    xnor g7489(n598 ,n7578 ,n7610);
    xnor g7490(n597 ,n7577 ,n7609);
    xnor g7491(n596 ,n7576 ,n7608);
    xnor g7492(n595 ,n7575 ,n7607);
    xnor g7493(n594 ,n7574 ,n7606);
    xnor g7494(n593 ,n7573 ,n7605);
    xnor g7495(n592 ,n7572 ,n7604);
    xnor g7496(n591 ,n7571 ,n7603);
    xnor g7497(n590 ,n7570 ,n7602);
    xnor g7498(n589 ,n7569 ,n7601);
    xnor g7499(n588 ,n7568 ,n7600);
    xnor g7500(n587 ,n7567 ,n7599);
    xnor g7501(n586 ,n7566 ,n7598);
    xnor g7502(n585 ,n7565 ,n7597);
    xnor g7503(n584 ,n7564 ,n7596);
    xnor g7504(n583 ,n7563 ,n7595);
    xnor g7505(n582 ,n7562 ,n7594);
    xnor g7506(n581 ,n7561 ,n7593);
    xnor g7507(n580 ,n7623 ,n7591);
    xnor g7508(n579 ,n7590 ,n7622);
    xnor g7509(n578 ,n7589 ,n7621);
    xnor g7510(n577 ,n7588 ,n7620);
    xnor g7511(n576 ,n7587 ,n7619);
    xnor g7512(n575 ,n7586 ,n7618);
    xnor g7513(n574 ,n7585 ,n7617);
    xnor g7514(n573 ,n7584 ,n7616);
    xnor g7515(n572 ,n7583 ,n7615);
    xnor g7516(n571 ,n7582 ,n7614);
    xnor g7517(n570 ,n7581 ,n7613);
    xnor g7518(n569 ,n7580 ,n7612);
    not g7519(n568 ,n567);
    nor g7520(n566 ,n474 ,n454);
    nor g7521(n565 ,n496 ,n500);
    nor g7522(n564 ,n467 ,n465);
    nor g7523(n563 ,n447 ,n477);
    nor g7524(n562 ,n470 ,n458);
    nor g7525(n561 ,n445 ,n484);
    nor g7526(n560 ,n488 ,n455);
    nor g7527(n559 ,n462 ,n502);
    nor g7528(n558 ,n478 ,n448);
    nor g7529(n557 ,n485 ,n501);
    nor g7530(n556 ,n466 ,n460);
    nor g7531(n555 ,n459 ,n487);
    nor g7532(n554 ,n471 ,n489);
    nor g7533(n553 ,n469 ,n476);
    nor g7534(n552 ,n456 ,n492);
    nor g7535(n551 ,n451 ,n483);
    nor g7536(n550 ,n490 ,n499);
    nor g7537(n549 ,n498 ,n504);
    nor g7538(n548 ,n486 ,n463);
    nor g7539(n547 ,n464 ,n503);
    nor g7540(n546 ,n497 ,n468);
    nor g7541(n545 ,n494 ,n472);
    nor g7542(n544 ,n482 ,n457);
    nor g7543(n543 ,n461 ,n479);
    nor g7544(n542 ,n495 ,n493);
    nor g7545(n541 ,n444 ,n452);
    nor g7546(n540 ,n453 ,n450);
    nor g7547(n539 ,n449 ,n480);
    nor g7548(n538 ,n481 ,n491);
    nor g7549(n537 ,n446 ,n473);
    nor g7550(n567 ,n505 ,n475);
    nor g7551(n536 ,n7615 ,n7583);
    nor g7552(n535 ,n7618 ,n7586);
    nor g7553(n534 ,n7611 ,n7579);
    nor g7554(n533 ,n7592 ,n7560);
    nor g7555(n532 ,n7606 ,n7574);
    nor g7556(n531 ,n7613 ,n7581);
    nor g7557(n530 ,n7600 ,n7568);
    nor g7558(n529 ,n7603 ,n7571);
    nor g7559(n528 ,n7598 ,n7566);
    nor g7560(n527 ,n7610 ,n7578);
    nor g7561(n526 ,n7612 ,n7580);
    nor g7562(n525 ,n7602 ,n7570);
    nor g7563(n524 ,n7594 ,n7562);
    nor g7564(n523 ,n7597 ,n7565);
    nor g7565(n522 ,n7614 ,n7582);
    nor g7566(n521 ,n7604 ,n7572);
    nor g7567(n520 ,n7621 ,n7589);
    nor g7568(n519 ,n7605 ,n7573);
    nor g7569(n518 ,n7617 ,n7585);
    nor g7570(n517 ,n7607 ,n7575);
    nor g7571(n516 ,n7593 ,n7561);
    nor g7572(n515 ,n7609 ,n7577);
    nor g7573(n514 ,n7608 ,n7576);
    nor g7574(n513 ,n7616 ,n7584);
    nor g7575(n512 ,n7620 ,n7588);
    nor g7576(n511 ,n7619 ,n7587);
    nor g7577(n510 ,n7622 ,n7590);
    nor g7578(n509 ,n7596 ,n7564);
    nor g7579(n508 ,n7595 ,n7563);
    nor g7580(n507 ,n7601 ,n7569);
    nor g7581(n506 ,n7599 ,n7567);
    not g7582(n505 ,n7592);
    not g7583(n504 ,n7575);
    not g7584(n503 ,n7561);
    not g7585(n502 ,n7579);
    not g7586(n501 ,n7590);
    not g7587(n500 ,n7570);
    not g7588(n499 ,n7581);
    not g7589(n498 ,n7607);
    not g7590(n497 ,n7606);
    not g7591(n496 ,n7602);
    not g7592(n495 ,n7614);
    not g7593(n494 ,n7616);
    not g7594(n493 ,n7582);
    not g7595(n492 ,n7562);
    not g7596(n491 ,n7589);
    not g7597(n490 ,n7613);
    not g7598(n489 ,n7578);
    not g7599(n488 ,n7609);
    not g7600(n487 ,n7566);
    not g7601(n486 ,n7615);
    not g7602(n485 ,n7622);
    not g7603(n484 ,n7569);
    not g7604(n483 ,n7576);
    not g7605(n482 ,n7619);
    not g7606(n481 ,n7621);
    not g7607(n480 ,n7580);
    not g7608(n479 ,n7573);
    not g7609(n478 ,n7600);
    not g7610(n477 ,n7586);
    not g7611(n476 ,n7564);
    not g7612(n475 ,n7560);
    not g7613(n474 ,n7597);
    not g7614(n473 ,n7571);
    not g7615(n472 ,n7584);
    not g7616(n471 ,n7610);
    not g7617(n470 ,n7617);
    not g7618(n469 ,n7596);
    not g7619(n468 ,n7574);
    not g7620(n467 ,n7595);
    not g7621(n466 ,n7599);
    not g7622(n465 ,n7563);
    not g7623(n464 ,n7593);
    not g7624(n463 ,n7583);
    not g7625(n462 ,n7611);
    not g7626(n461 ,n7605);
    not g7627(n460 ,n7567);
    not g7628(n459 ,n7598);
    not g7629(n458 ,n7585);
    not g7630(n457 ,n7587);
    not g7631(n456 ,n7594);
    not g7632(n455 ,n7577);
    not g7633(n454 ,n7565);
    not g7634(n453 ,n7604);
    not g7635(n452 ,n7588);
    not g7636(n451 ,n7608);
    not g7637(n450 ,n7572);
    not g7638(n449 ,n7612);
    not g7639(n448 ,n7568);
    not g7640(n447 ,n7618);
    not g7641(n446 ,n7603);
    not g7642(n445 ,n7601);
    not g7643(n444 ,n7620);
    xor g7644(n7526 ,n796 ,n875);
    nor g7645(n875 ,n773 ,n874);
    xor g7646(n7522 ,n795 ,n873);
    nor g7647(n874 ,n726 ,n873);
    nor g7648(n873 ,n754 ,n872);
    xor g7649(n7518 ,n794 ,n871);
    nor g7650(n872 ,n736 ,n871);
    nor g7651(n871 ,n757 ,n870);
    xor g7652(n7514 ,n793 ,n869);
    nor g7653(n870 ,n728 ,n869);
    nor g7654(n869 ,n760 ,n868);
    xor g7655(n7510 ,n792 ,n867);
    nor g7656(n868 ,n727 ,n867);
    nor g7657(n867 ,n779 ,n866);
    xor g7658(n7506 ,n791 ,n865);
    nor g7659(n866 ,n751 ,n865);
    nor g7660(n865 ,n778 ,n864);
    xor g7661(n7502 ,n790 ,n863);
    nor g7662(n864 ,n734 ,n863);
    nor g7663(n863 ,n761 ,n862);
    xor g7664(n7498 ,n789 ,n861);
    nor g7665(n862 ,n729 ,n861);
    nor g7666(n861 ,n764 ,n860);
    xor g7667(n7494 ,n788 ,n859);
    nor g7668(n860 ,n752 ,n859);
    nor g7669(n859 ,n758 ,n858);
    xor g7670(n7490 ,n787 ,n857);
    nor g7671(n858 ,n738 ,n857);
    nor g7672(n857 ,n766 ,n856);
    xor g7673(n7486 ,n786 ,n855);
    nor g7674(n856 ,n747 ,n855);
    nor g7675(n855 ,n755 ,n854);
    xor g7676(n7482 ,n785 ,n853);
    nor g7677(n854 ,n742 ,n853);
    nor g7678(n853 ,n775 ,n852);
    xor g7679(n7478 ,n815 ,n851);
    nor g7680(n852 ,n750 ,n851);
    nor g7681(n851 ,n770 ,n850);
    xor g7682(n7474 ,n814 ,n849);
    nor g7683(n850 ,n743 ,n849);
    nor g7684(n849 ,n776 ,n848);
    xor g7685(n7470 ,n813 ,n847);
    nor g7686(n848 ,n731 ,n847);
    nor g7687(n847 ,n767 ,n846);
    xor g7688(n7466 ,n812 ,n845);
    nor g7689(n846 ,n730 ,n845);
    nor g7690(n845 ,n765 ,n844);
    xor g7691(n7462 ,n811 ,n843);
    nor g7692(n844 ,n733 ,n843);
    nor g7693(n843 ,n762 ,n842);
    xor g7694(n7458 ,n810 ,n841);
    nor g7695(n842 ,n748 ,n841);
    nor g7696(n841 ,n759 ,n840);
    xor g7697(n7454 ,n809 ,n839);
    nor g7698(n840 ,n735 ,n839);
    nor g7699(n839 ,n756 ,n838);
    xor g7700(n7450 ,n808 ,n837);
    nor g7701(n838 ,n737 ,n837);
    nor g7702(n837 ,n753 ,n836);
    xor g7703(n7446 ,n807 ,n835);
    nor g7704(n836 ,n745 ,n835);
    nor g7705(n835 ,n781 ,n834);
    xor g7706(n7442 ,n806 ,n833);
    nor g7707(n834 ,n741 ,n833);
    nor g7708(n833 ,n777 ,n832);
    xor g7709(n7438 ,n805 ,n831);
    nor g7710(n832 ,n723 ,n831);
    nor g7711(n831 ,n774 ,n830);
    xor g7712(n7434 ,n804 ,n829);
    nor g7713(n830 ,n746 ,n829);
    nor g7714(n829 ,n772 ,n828);
    xor g7715(n7430 ,n803 ,n827);
    nor g7716(n828 ,n722 ,n827);
    nor g7717(n827 ,n771 ,n826);
    xor g7718(n7426 ,n802 ,n825);
    nor g7719(n826 ,n744 ,n825);
    nor g7720(n825 ,n782 ,n824);
    xor g7721(n7422 ,n801 ,n823);
    nor g7722(n824 ,n739 ,n823);
    nor g7723(n823 ,n769 ,n822);
    xor g7724(n7418 ,n800 ,n821);
    nor g7725(n822 ,n725 ,n821);
    nor g7726(n821 ,n780 ,n820);
    xor g7727(n7414 ,n799 ,n819);
    nor g7728(n820 ,n724 ,n819);
    nor g7729(n819 ,n768 ,n818);
    xor g7730(n7410 ,n798 ,n817);
    nor g7731(n818 ,n740 ,n817);
    xnor g7732(n7406 ,n797 ,n783);
    nor g7733(n817 ,n763 ,n816);
    nor g7734(n7402 ,n783 ,n749);
    nor g7735(n816 ,n784 ,n732);
    xnor g7736(n815 ,n7546 ,n0[115]);
    xnor g7737(n814 ,n7545 ,n0[114]);
    xnor g7738(n813 ,n7544 ,n0[113]);
    xnor g7739(n812 ,n7543 ,n0[112]);
    xnor g7740(n811 ,n7542 ,n0[111]);
    xnor g7741(n810 ,n7541 ,n0[110]);
    xnor g7742(n809 ,n7540 ,n0[109]);
    xnor g7743(n808 ,n7539 ,n0[108]);
    xnor g7744(n807 ,n7538 ,n0[107]);
    xnor g7745(n806 ,n7537 ,n0[106]);
    xnor g7746(n805 ,n7536 ,n0[105]);
    xnor g7747(n804 ,n7535 ,n0[104]);
    xnor g7748(n803 ,n7534 ,n0[103]);
    xnor g7749(n802 ,n7533 ,n0[102]);
    xnor g7750(n801 ,n7532 ,n0[101]);
    xnor g7751(n800 ,n7531 ,n0[100]);
    xnor g7752(n799 ,n7530 ,n0[99]);
    xnor g7753(n798 ,n7529 ,n0[98]);
    xnor g7754(n797 ,n7528 ,n0[97]);
    xnor g7755(n796 ,n0[127] ,n7558);
    xnor g7756(n795 ,n7557 ,n0[126]);
    xnor g7757(n794 ,n7556 ,n0[125]);
    xnor g7758(n793 ,n7555 ,n0[124]);
    xnor g7759(n792 ,n7554 ,n0[123]);
    xnor g7760(n791 ,n7553 ,n0[122]);
    xnor g7761(n790 ,n7552 ,n0[121]);
    xnor g7762(n789 ,n7551 ,n0[120]);
    xnor g7763(n788 ,n7550 ,n0[119]);
    xnor g7764(n787 ,n7549 ,n0[118]);
    xnor g7765(n786 ,n7548 ,n0[117]);
    xnor g7766(n785 ,n7547 ,n0[116]);
    not g7767(n784 ,n783);
    nor g7768(n782 ,n690 ,n670);
    nor g7769(n781 ,n712 ,n716);
    nor g7770(n780 ,n683 ,n681);
    nor g7771(n779 ,n663 ,n693);
    nor g7772(n778 ,n686 ,n674);
    nor g7773(n777 ,n661 ,n700);
    nor g7774(n776 ,n704 ,n671);
    nor g7775(n775 ,n678 ,n718);
    nor g7776(n774 ,n694 ,n664);
    nor g7777(n773 ,n701 ,n717);
    nor g7778(n772 ,n682 ,n676);
    nor g7779(n771 ,n675 ,n703);
    nor g7780(n770 ,n687 ,n705);
    nor g7781(n769 ,n685 ,n692);
    nor g7782(n768 ,n672 ,n708);
    nor g7783(n767 ,n667 ,n699);
    nor g7784(n766 ,n706 ,n715);
    nor g7785(n765 ,n714 ,n720);
    nor g7786(n764 ,n702 ,n679);
    nor g7787(n763 ,n680 ,n719);
    nor g7788(n762 ,n713 ,n684);
    nor g7789(n761 ,n710 ,n688);
    nor g7790(n760 ,n698 ,n673);
    nor g7791(n759 ,n677 ,n695);
    nor g7792(n758 ,n711 ,n709);
    nor g7793(n757 ,n660 ,n668);
    nor g7794(n756 ,n669 ,n666);
    nor g7795(n755 ,n665 ,n696);
    nor g7796(n754 ,n697 ,n707);
    nor g7797(n753 ,n662 ,n689);
    nor g7798(n783 ,n721 ,n691);
    nor g7799(n752 ,n0[119] ,n7550);
    nor g7800(n751 ,n0[122] ,n7553);
    nor g7801(n750 ,n0[115] ,n7546);
    nor g7802(n749 ,n0[96] ,n7527);
    nor g7803(n748 ,n0[110] ,n7541);
    nor g7804(n747 ,n0[117] ,n7548);
    nor g7805(n746 ,n0[104] ,n7535);
    nor g7806(n745 ,n0[107] ,n7538);
    nor g7807(n744 ,n0[102] ,n7533);
    nor g7808(n743 ,n0[114] ,n7545);
    nor g7809(n742 ,n0[116] ,n7547);
    nor g7810(n741 ,n0[106] ,n7537);
    nor g7811(n740 ,n0[98] ,n7529);
    nor g7812(n739 ,n0[101] ,n7532);
    nor g7813(n738 ,n0[118] ,n7549);
    nor g7814(n737 ,n0[108] ,n7539);
    nor g7815(n736 ,n0[125] ,n7556);
    nor g7816(n735 ,n0[109] ,n7540);
    nor g7817(n734 ,n0[121] ,n7552);
    nor g7818(n733 ,n0[111] ,n7542);
    nor g7819(n732 ,n0[97] ,n7528);
    nor g7820(n731 ,n0[113] ,n7544);
    nor g7821(n730 ,n0[112] ,n7543);
    nor g7822(n729 ,n0[120] ,n7551);
    nor g7823(n728 ,n0[124] ,n7555);
    nor g7824(n727 ,n0[123] ,n7554);
    nor g7825(n726 ,n0[126] ,n7557);
    nor g7826(n725 ,n0[100] ,n7531);
    nor g7827(n724 ,n0[99] ,n7530);
    nor g7828(n723 ,n0[105] ,n7536);
    nor g7829(n722 ,n0[103] ,n7534);
    not g7830(n721 ,n0[96]);
    not g7831(n720 ,n7542);
    not g7832(n719 ,n7528);
    not g7833(n718 ,n7546);
    not g7834(n717 ,n7557);
    not g7835(n716 ,n7537);
    not g7836(n715 ,n7548);
    not g7837(n714 ,n0[111]);
    not g7838(n713 ,n0[110]);
    not g7839(n712 ,n0[106]);
    not g7840(n711 ,n0[118]);
    not g7841(n710 ,n0[120]);
    not g7842(n709 ,n7549);
    not g7843(n708 ,n7529);
    not g7844(n707 ,n7556);
    not g7845(n706 ,n0[117]);
    not g7846(n705 ,n7545);
    not g7847(n704 ,n0[113]);
    not g7848(n703 ,n7533);
    not g7849(n702 ,n0[119]);
    not g7850(n701 ,n0[126]);
    not g7851(n700 ,n7536);
    not g7852(n699 ,n7543);
    not g7853(n698 ,n0[123]);
    not g7854(n697 ,n0[125]);
    not g7855(n696 ,n7547);
    not g7856(n695 ,n7540);
    not g7857(n694 ,n0[104]);
    not g7858(n693 ,n7553);
    not g7859(n692 ,n7531);
    not g7860(n691 ,n7527);
    not g7861(n690 ,n0[101]);
    not g7862(n689 ,n7538);
    not g7863(n688 ,n7551);
    not g7864(n687 ,n0[114]);
    not g7865(n686 ,n0[121]);
    not g7866(n685 ,n0[100]);
    not g7867(n684 ,n7541);
    not g7868(n683 ,n0[99]);
    not g7869(n682 ,n0[103]);
    not g7870(n681 ,n7530);
    not g7871(n680 ,n0[97]);
    not g7872(n679 ,n7550);
    not g7873(n678 ,n0[115]);
    not g7874(n677 ,n0[109]);
    not g7875(n676 ,n7534);
    not g7876(n675 ,n0[102]);
    not g7877(n674 ,n7552);
    not g7878(n673 ,n7554);
    not g7879(n672 ,n0[98]);
    not g7880(n671 ,n7544);
    not g7881(n670 ,n7532);
    not g7882(n669 ,n0[108]);
    not g7883(n668 ,n7555);
    not g7884(n667 ,n0[112]);
    not g7885(n666 ,n7539);
    not g7886(n665 ,n0[116]);
    not g7887(n664 ,n7535);
    not g7888(n663 ,n0[122]);
    not g7889(n662 ,n0[107]);
    not g7890(n661 ,n0[105]);
    not g7891(n660 ,n0[124]);
endmodule
