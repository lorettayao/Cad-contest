module top(n0, n1, n4, n6, n5, n2, n11, n12, n13, n14, n17, n15, n16, n3, n7, n8, n9, n10);
    input n0, n1, n2, n3;
    input [7:0] n4;
    input [3:0] n5;
    output [7:0] n6, n7, n8, n9, n10;
    output n11, n12, n13, n14, n15, n16;
    output [3:0] n17;
    wire n0, n1, n2, n3;
    wire [7:0] n4;
    wire [3:0] n5;
    wire [7:0] n6, n7, n8, n9, n10;
    wire n11, n12, n13, n14, n15, n16;
    wire [3:0] n17;
    wire [3:0] n18;
    wire [3:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [4:0] n22;
    wire [3:0] n23;
    wire [3:0] n24;
    wire [7:0] n25;
    wire [2:0] n26;
    wire [7:0] n27;
    wire [7:0] n28;
    wire [7:0] n29;
    wire [7:0] n30;
    wire [7:0] n31;
    wire [7:0] n32;
    wire [7:0] n33;
    wire [7:0] n34;
    wire [7:0] n35;
    wire [7:0] n36;
    wire [7:0] n37;
    wire [7:0] n38;
    wire [7:0] n39;
    wire [7:0] n40;
    wire [7:0] n41;
    wire [7:0] n42;
    wire [4:0] n43;
    wire [3:0] n44;
    wire [3:0] n45;
    wire [7:0] n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    buf g0(n45[3], 1'b0);
    buf g1(n45[2], 1'b0);
    buf g2(n45[1], 1'b0);
    buf g3(n45[0], 1'b0);
    buf g4(n23[3], 1'b0);
    buf g5(n23[2], 1'b0);
    buf g6(n23[1], 1'b0);
    buf g7(n23[0], 1'b0);
    buf g8(n10[0], 1'b0);
    buf g9(n10[1], 1'b0);
    buf g10(n10[2], 1'b0);
    buf g11(n10[3], 1'b0);
    buf g12(n10[4], n7[7]);
    buf g13(n10[5], n7[7]);
    buf g14(n9[0], 1'b0);
    buf g15(n9[1], 1'b0);
    buf g16(n9[2], 1'b0);
    buf g17(n9[3], 1'b0);
    buf g18(n9[4], 1'b0);
    buf g19(n9[5], 1'b0);
    buf g20(n9[6], 1'b0);
    buf g21(n9[7], 1'b0);
    buf g22(n8[0], 1'b0);
    buf g23(n8[1], 1'b0);
    buf g24(n8[2], 1'b0);
    buf g25(n8[3], 1'b0);
    buf g26(n8[4], 1'b0);
    buf g27(n8[5], 1'b0);
    buf g28(n8[6], 1'b0);
    buf g29(n8[7], 1'b0);
    buf g30(n7[0], 1'b0);
    buf g31(n7[1], 1'b0);
    buf g32(n7[6], n7[7]);
    buf g33(n14, n13);
    not g34(n1518 ,n1537);
    not g35(n1517 ,n1533);
    not g36(n1516 ,n3);
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1157), .Q(n18[0]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1145), .Q(n18[1]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1119), .Q(n18[2]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1115), .Q(n18[3]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n513), .Q(n19[0]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n606), .Q(n19[1]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n740), .Q(n17[0]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n737), .Q(n17[1]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n748), .Q(n17[2]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n742), .Q(n17[3]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n422), .Q(n7[7]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n402), .Q(n10[6]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n405), .Q(n10[7]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n732), .Q(n16));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n580), .Q(n13));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n627), .Q(n6[0]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n633), .Q(n6[1]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n626), .Q(n6[2]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n635), .Q(n6[3]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n629), .Q(n6[4]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n632), .Q(n6[5]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n630), .Q(n6[6]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n631), .Q(n6[7]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n12));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1480), .Q(n20[0]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1477), .Q(n20[1]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1479), .Q(n20[2]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1478), .Q(n20[3]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1476), .Q(n20[4]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1473), .Q(n20[5]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1475), .Q(n20[6]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1474), .Q(n20[7]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n21[0]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1413), .Q(n21[1]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n21[2]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n21[3]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1410), .Q(n21[4]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n21[5]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n21[6]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n21[7]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1369), .Q(n22[0]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n507), .Q(n22[0]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1368), .Q(n22[1]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n511), .Q(n22[1]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n22[2]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n510), .Q(n22[2]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n22[3]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n506), .Q(n22[3]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n22[4]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n505), .Q(n22[4]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n647), .Q(n23[0]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n648), .Q(n23[1]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n649), .Q(n23[2]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n650), .Q(n23[3]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n24[0]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n24[1]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n24[2]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n24[3]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n25[0]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1312), .Q(n25[1]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n25[2]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n25[3]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1315), .Q(n25[4]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1044), .Q(n25[5]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n25[6]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1184), .Q(n25[7]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n751), .Q(n15));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n739), .Q(n26[0]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n638), .Q(n26[1]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n616), .Q(n7[2]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n578), .Q(n7[3]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n617), .Q(n7[4]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n618), .Q(n7[5]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n11));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1171), .Q(n27[0]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1167), .Q(n27[1]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1162), .Q(n27[2]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1160), .Q(n27[3]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1156), .Q(n27[4]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1153), .Q(n27[5]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1147), .Q(n27[6]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1144), .Q(n27[7]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1141), .Q(n28[0]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1137), .Q(n28[1]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1134), .Q(n28[2]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1131), .Q(n28[3]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1129), .Q(n28[4]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1128), .Q(n28[5]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1127), .Q(n28[6]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1126), .Q(n28[7]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1124), .Q(n29[0]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1122), .Q(n29[1]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1121), .Q(n29[2]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1120), .Q(n29[3]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1118), .Q(n29[4]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1117), .Q(n29[5]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1116), .Q(n29[6]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1113), .Q(n29[7]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1112), .Q(n30[0]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1111), .Q(n30[1]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1110), .Q(n30[2]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1108), .Q(n30[3]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1107), .Q(n30[4]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1106), .Q(n30[5]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1104), .Q(n30[6]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1123), .Q(n30[7]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1130), .Q(n31[0]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1149), .Q(n31[1]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1154), .Q(n31[2]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1183), .Q(n31[3]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1103), .Q(n31[4]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1102), .Q(n31[5]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1101), .Q(n31[6]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1098), .Q(n31[7]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1105), .Q(n32[0]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1066), .Q(n32[1]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1095), .Q(n32[2]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1094), .Q(n32[3]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1093), .Q(n32[4]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1092), .Q(n32[5]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1091), .Q(n32[6]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1088), .Q(n32[7]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1114), .Q(n33[0]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1089), .Q(n33[1]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1125), .Q(n33[2]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1086), .Q(n33[3]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1085), .Q(n33[4]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1084), .Q(n33[5]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1082), .Q(n33[6]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1081), .Q(n33[7]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1079), .Q(n34[0]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1080), .Q(n34[1]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1078), .Q(n34[2]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1077), .Q(n34[3]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1076), .Q(n34[4]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1075), .Q(n34[5]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1074), .Q(n34[6]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1073), .Q(n34[7]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1072), .Q(n35[0]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1071), .Q(n35[1]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1070), .Q(n35[2]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1069), .Q(n35[3]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1068), .Q(n35[4]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1067), .Q(n35[5]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1065), .Q(n35[6]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1064), .Q(n35[7]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1063), .Q(n36[0]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1062), .Q(n36[1]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1061), .Q(n36[2]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1060), .Q(n36[3]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1059), .Q(n36[4]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1058), .Q(n36[5]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1057), .Q(n36[6]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1056), .Q(n36[7]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1055), .Q(n37[0]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1054), .Q(n37[1]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1053), .Q(n37[2]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1052), .Q(n37[3]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1051), .Q(n37[4]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1050), .Q(n37[5]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1049), .Q(n37[6]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1048), .Q(n37[7]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1047), .Q(n38[0]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1046), .Q(n38[1]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1045), .Q(n38[2]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1185), .Q(n38[3]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1180), .Q(n38[4]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1182), .Q(n38[5]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1181), .Q(n38[6]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1179), .Q(n38[7]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1178), .Q(n39[0]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1177), .Q(n39[1]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1176), .Q(n39[2]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1175), .Q(n39[3]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1174), .Q(n39[4]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1173), .Q(n39[5]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1172), .Q(n39[6]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1170), .Q(n39[7]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1169), .Q(n40[0]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1168), .Q(n40[1]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1166), .Q(n40[2]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1165), .Q(n40[3]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1164), .Q(n40[4]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1163), .Q(n40[5]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1161), .Q(n40[6]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1159), .Q(n40[7]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1158), .Q(n41[0]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1155), .Q(n41[1]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1152), .Q(n41[2]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1151), .Q(n41[3]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1150), .Q(n41[4]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1148), .Q(n41[5]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1146), .Q(n41[6]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1143), .Q(n41[7]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1142), .Q(n42[0]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1140), .Q(n42[1]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1139), .Q(n42[2]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1138), .Q(n42[3]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1136), .Q(n42[4]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1135), .Q(n42[5]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1133), .Q(n42[6]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1132), .Q(n42[7]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n640), .Q(n43[0]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n581), .Q(n43[0]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n641), .Q(n43[1]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n584), .Q(n43[1]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n642), .Q(n43[2]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n583), .Q(n43[2]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n643), .Q(n43[3]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n582), .Q(n43[3]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n644), .Q(n43[4]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n579), .Q(n43[4]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n645), .Q(n44[0]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n44[1]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n44[2]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1415), .Q(n44[3]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n45[0]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1362), .Q(n45[1]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n45[2]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1360), .Q(n45[3]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1513), .Q(n46[0]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1514), .Q(n46[1]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1515), .Q(n46[2]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1507), .Q(n46[3]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1510), .Q(n46[4]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1511), .Q(n46[5]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1509), .Q(n46[6]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1512), .Q(n46[7]));
    or g265(n1515 ,n1503 ,n1489);
    or g266(n1514 ,n1491 ,n1502);
    or g267(n1513 ,n1434 ,n1506);
    or g268(n1512 ,n1483 ,n1501);
    or g269(n1511 ,n1437 ,n1505);
    or g270(n1510 ,n1436 ,n1508);
    or g271(n1509 ,n1485 ,n1504);
    or g272(n1508 ,n1424 ,n1500);
    or g273(n1507 ,n1430 ,n1499);
    or g274(n1506 ,n1357 ,n1498);
    or g275(n1505 ,n1422 ,n1495);
    or g276(n1504 ,n1275 ,n1494);
    or g277(n1503 ,n1247 ,n1496);
    or g278(n1502 ,n1256 ,n1497);
    or g279(n1501 ,n1284 ,n1493);
    or g280(n1500 ,n1202 ,n1487);
    or g281(n1499 ,n1425 ,n1488);
    or g282(n1498 ,n1272 ,n1492);
    or g283(n1497 ,n1255 ,n1490);
    or g284(n1496 ,n741 ,n1481);
    or g285(n1495 ,n1208 ,n1486);
    or g286(n1494 ,n1201 ,n1484);
    or g287(n1493 ,n1193 ,n1482);
    or g288(n1492 ,n1356 ,n1456);
    or g289(n1491 ,n1372 ,n1451);
    or g290(n1490 ,n1350 ,n1450);
    or g291(n1489 ,n1347 ,n1466);
    or g292(n1488 ,n1429 ,n1454);
    or g293(n1487 ,n1371 ,n1448);
    or g294(n1486 ,n1370 ,n1446);
    or g295(n1485 ,n744 ,n1447);
    or g296(n1484 ,n1326 ,n1453);
    or g297(n1483 ,n743 ,n1445);
    or g298(n1482 ,n1398 ,n1452);
    or g299(n1481 ,n1292 ,n1449);
    or g300(n1480 ,n1464 ,n1467);
    or g301(n1479 ,n1462 ,n1469);
    or g302(n1478 ,n1461 ,n1470);
    or g303(n1477 ,n1463 ,n1468);
    or g304(n1476 ,n1460 ,n1471);
    or g305(n1475 ,n1458 ,n1455);
    or g306(n1474 ,n1457 ,n1465);
    or g307(n1473 ,n1459 ,n1472);
    nor g308(n1472 ,n142 ,n1443);
    nor g309(n1471 ,n148 ,n1443);
    nor g310(n1470 ,n265 ,n1443);
    nor g311(n1469 ,n145 ,n1443);
    nor g312(n1468 ,n268 ,n1443);
    nor g313(n1467 ,n269 ,n1443);
    or g314(n1466 ,n1432 ,n1431);
    nor g315(n1465 ,n274 ,n1443);
    nor g316(n1464 ,n307 ,n1444);
    nor g317(n1463 ,n194 ,n1444);
    nor g318(n1462 ,n388 ,n1444);
    nor g319(n1461 ,n308 ,n1444);
    nor g320(n1460 ,n213 ,n1444);
    nor g321(n1459 ,n303 ,n1444);
    nor g322(n1458 ,n369 ,n1444);
    nor g323(n1457 ,n286 ,n1444);
    or g324(n1456 ,n1442 ,n1433);
    nor g325(n1455 ,n144 ,n1443);
    or g326(n1454 ,n1337 ,n1435);
    or g327(n1453 ,n1438 ,n1439);
    or g328(n1452 ,n1441 ,n1440);
    or g329(n1451 ,n1260 ,n1416);
    or g330(n1450 ,n1243 ,n1427);
    or g331(n1449 ,n1246 ,n1426);
    or g332(n1448 ,n1219 ,n1423);
    or g333(n1447 ,n1301 ,n1420);
    or g334(n1446 ,n1207 ,n1421);
    or g335(n1445 ,n1285 ,n1419);
    not g336(n1443 ,n1444);
    or g337(n1442 ,n1355 ,n1354);
    or g338(n1441 ,n1399 ,n1400);
    or g339(n1440 ,n1401 ,n1402);
    or g340(n1439 ,n1323 ,n1396);
    or g341(n1438 ,n1325 ,n1324);
    or g342(n1437 ,n1331 ,n1330);
    or g343(n1436 ,n1335 ,n1334);
    or g344(n1435 ,n735 ,n1336);
    or g345(n1434 ,n1359 ,n1358);
    or g346(n1433 ,n1353 ,n1352);
    or g347(n1432 ,n1346 ,n1345);
    or g348(n1431 ,n1344 ,n1343);
    or g349(n1430 ,n1342 ,n1341);
    or g350(n1429 ,n1339 ,n1338);
    nor g351(n1444 ,n403 ,n1373);
    or g352(n1428 ,n612 ,n1394);
    or g353(n1427 ,n1251 ,n1349);
    or g354(n1426 ,n1302 ,n1348);
    or g355(n1425 ,n1235 ,n1340);
    or g356(n1424 ,n1222 ,n1333);
    or g357(n1423 ,n1218 ,n1332);
    or g358(n1422 ,n1211 ,n1329);
    or g359(n1421 ,n1206 ,n1328);
    or g360(n1420 ,n1228 ,n1327);
    or g361(n1419 ,n1254 ,n1397);
    nor g362(n1418 ,n123 ,n1364);
    or g363(n1417 ,n603 ,n1395);
    or g364(n1416 ,n1259 ,n1351);
    or g365(n1415 ,n602 ,n1393);
    or g366(n1414 ,n1381 ,n1389);
    or g367(n1413 ,n1380 ,n1388);
    or g368(n1412 ,n1379 ,n1387);
    or g369(n1411 ,n1378 ,n1386);
    or g370(n1410 ,n1377 ,n1385);
    or g371(n1409 ,n1376 ,n1384);
    or g372(n1408 ,n1375 ,n1383);
    or g373(n1407 ,n1374 ,n1382);
    or g374(n1406 ,n1299 ,n1392);
    or g375(n1405 ,n1297 ,n1390);
    or g376(n1404 ,n1298 ,n1391);
    or g377(n1403 ,n525 ,n1308);
    or g378(n1402 ,n1232 ,n1187);
    or g379(n1401 ,n1188 ,n1189);
    or g380(n1400 ,n1303 ,n1190);
    or g381(n1399 ,n1283 ,n1248);
    or g382(n1398 ,n1192 ,n1191);
    or g383(n1397 ,n1194 ,n1274);
    or g384(n1396 ,n1261 ,n1195);
    nor g385(n1395 ,n244 ,n1320);
    nor g386(n1394 ,n230 ,n1320);
    nor g387(n1393 ,n256 ,n1320);
    nor g388(n1392 ,n242 ,n1319);
    nor g389(n1391 ,n235 ,n1319);
    nor g390(n1390 ,n259 ,n1319);
    nor g391(n1389 ,n269 ,n1317);
    nor g392(n1388 ,n268 ,n1317);
    nor g393(n1387 ,n145 ,n1317);
    nor g394(n1386 ,n265 ,n1317);
    nor g395(n1385 ,n148 ,n1317);
    nor g396(n1384 ,n142 ,n1317);
    nor g397(n1383 ,n144 ,n1317);
    nor g398(n1382 ,n274 ,n1317);
    nor g399(n1381 ,n218 ,n1318);
    nor g400(n1380 ,n391 ,n1318);
    nor g401(n1379 ,n322 ,n1318);
    nor g402(n1378 ,n167 ,n1318);
    nor g403(n1377 ,n177 ,n1318);
    nor g404(n1376 ,n287 ,n1318);
    nor g405(n1375 ,n396 ,n1318);
    nor g406(n1374 ,n394 ,n1318);
    or g407(n1373 ,n24[3] ,n1322);
    or g408(n1372 ,n707 ,n1109);
    or g409(n1371 ,n702 ,n1100);
    or g410(n1370 ,n703 ,n1097);
    nor g411(n1369 ,n127 ,n1099);
    nor g412(n1368 ,n126 ,n1096);
    nor g413(n1367 ,n123 ,n1090);
    nor g414(n1366 ,n123 ,n1087);
    nor g415(n1365 ,n124 ,n1083);
    nor g416(n1364 ,n1186 ,n1309);
    or g417(n1363 ,n1300 ,n1321);
    or g418(n1362 ,n524 ,n1307);
    or g419(n1361 ,n523 ,n1306);
    or g420(n1360 ,n564 ,n1305);
    or g421(n1359 ,n1295 ,n1294);
    or g422(n1358 ,n1293 ,n1304);
    or g423(n1357 ,n1273 ,n727);
    or g424(n1356 ,n1271 ,n1270);
    or g425(n1355 ,n1269 ,n1268);
    or g426(n1354 ,n1267 ,n1266);
    or g427(n1353 ,n1265 ,n1264);
    or g428(n1352 ,n1263 ,n1262);
    or g429(n1351 ,n1257 ,n1258);
    or g430(n1350 ,n1252 ,n1253);
    or g431(n1349 ,n1250 ,n1249);
    or g432(n1348 ,n1245 ,n1244);
    or g433(n1347 ,n1242 ,n1241);
    or g434(n1346 ,n1240 ,n1239);
    or g435(n1345 ,n1279 ,n1277);
    or g436(n1344 ,n1290 ,n1278);
    or g437(n1343 ,n1289 ,n1238);
    or g438(n1342 ,n1288 ,n1296);
    or g439(n1341 ,n1237 ,n1236);
    or g440(n1340 ,n1234 ,n1233);
    or g441(n1339 ,n1230 ,n1231);
    or g442(n1338 ,n1282 ,n1229);
    or g443(n1337 ,n1281 ,n1227);
    or g444(n1336 ,n1226 ,n729);
    or g445(n1335 ,n1224 ,n1225);
    or g446(n1334 ,n1280 ,n1223);
    or g447(n1333 ,n1221 ,n1220);
    or g448(n1332 ,n1216 ,n1217);
    or g449(n1331 ,n1215 ,n1214);
    or g450(n1330 ,n1213 ,n1212);
    or g451(n1329 ,n1210 ,n1209);
    or g452(n1328 ,n1205 ,n1276);
    or g453(n1327 ,n1287 ,n1203);
    or g454(n1326 ,n1286 ,n1200);
    or g455(n1325 ,n1199 ,n1204);
    or g456(n1324 ,n1291 ,n1198);
    or g457(n1323 ,n1197 ,n1196);
    not g458(n1322 ,n1321);
    not g459(n1317 ,n1318);
    nor g460(n1316 ,n125 ,n750);
    nor g461(n1315 ,n125 ,n749);
    nor g462(n1314 ,n127 ,n747);
    nor g463(n1313 ,n126 ,n738);
    nor g464(n1312 ,n125 ,n746);
    nor g465(n1311 ,n125 ,n745);
    nor g466(n1310 ,n127 ,n734);
    nor g467(n1309 ,n360 ,n896);
    nor g468(n1308 ,n231 ,n891);
    nor g469(n1307 ,n225 ,n891);
    nor g470(n1306 ,n224 ,n891);
    nor g471(n1305 ,n233 ,n891);
    nor g472(n1304 ,n354 ,n893);
    nor g473(n1303 ,n331 ,n893);
    nor g474(n1302 ,n325 ,n893);
    nor g475(n1301 ,n321 ,n893);
    nor g476(n1300 ,n143 ,n892);
    nor g477(n1299 ,n266 ,n892);
    nor g478(n1298 ,n270 ,n892);
    nor g479(n1297 ,n267 ,n892);
    nor g480(n1296 ,n279 ,n889);
    nor g481(n1295 ,n310 ,n888);
    nor g482(n1294 ,n168 ,n890);
    nor g483(n1293 ,n305 ,n889);
    nor g484(n1292 ,n208 ,n888);
    nor g485(n1291 ,n349 ,n890);
    nor g486(n1290 ,n329 ,n889);
    nor g487(n1289 ,n198 ,n890);
    nor g488(n1288 ,n294 ,n890);
    nor g489(n1287 ,n280 ,n889);
    nor g490(n1286 ,n219 ,n888);
    nor g491(n1285 ,n210 ,n890);
    nor g492(n1284 ,n380 ,n888);
    nor g493(n1283 ,n362 ,n889);
    nor g494(n1282 ,n393 ,n879);
    nor g495(n1281 ,n164 ,n876);
    nor g496(n1280 ,n299 ,n876);
    nor g497(n1279 ,n170 ,n886);
    nor g498(n1278 ,n327 ,n878);
    nor g499(n1277 ,n357 ,n875);
    nor g500(n1276 ,n277 ,n880);
    nor g501(n1275 ,n348 ,n883);
    nor g502(n1274 ,n173 ,n881);
    nor g503(n1273 ,n293 ,n883);
    nor g504(n1272 ,n203 ,n880);
    nor g505(n1271 ,n206 ,n881);
    nor g506(n1270 ,n342 ,n877);
    nor g507(n1269 ,n304 ,n882);
    nor g508(n1268 ,n184 ,n878);
    nor g509(n1267 ,n355 ,n876);
    nor g510(n1266 ,n165 ,n875);
    nor g511(n1265 ,n371 ,n879);
    nor g512(n1264 ,n281 ,n886);
    nor g513(n1263 ,n337 ,n884);
    nor g514(n1262 ,n155 ,n885);
    nor g515(n1261 ,n392 ,n886);
    nor g516(n1260 ,n166 ,n886);
    nor g517(n1259 ,n365 ,n885);
    nor g518(n1258 ,n161 ,n880);
    nor g519(n1257 ,n306 ,n875);
    nor g520(n1256 ,n328 ,n879);
    nor g521(n1255 ,n296 ,n878);
    nor g522(n1254 ,n159 ,n884);
    nor g523(n1253 ,n343 ,n876);
    nor g524(n1252 ,n200 ,n883);
    nor g525(n1251 ,n181 ,n884);
    nor g526(n1250 ,n358 ,n882);
    nor g527(n1249 ,n313 ,n877);
    nor g528(n1248 ,n163 ,n877);
    nor g529(n1247 ,n320 ,n877);
    nor g530(n1246 ,n372 ,n883);
    nor g531(n1245 ,n376 ,n879);
    nor g532(n1244 ,n366 ,n881);
    nor g533(n1243 ,n318 ,n881);
    nor g534(n1242 ,n323 ,n884);
    nor g535(n1241 ,n384 ,n880);
    nor g536(n1240 ,n202 ,n882);
    nor g537(n1239 ,n340 ,n876);
    nor g538(n1238 ,n330 ,n885);
    nor g539(n1237 ,n336 ,n881);
    nor g540(n1236 ,n332 ,n884);
    nor g541(n1235 ,n386 ,n877);
    nor g542(n1234 ,n178 ,n886);
    nor g543(n1233 ,n350 ,n875);
    nor g544(n1232 ,n383 ,n880);
    nor g545(n1231 ,n364 ,n880);
    nor g546(n1230 ,n215 ,n882);
    nor g547(n1229 ,n179 ,n885);
    nor g548(n1228 ,n187 ,n884);
    nor g549(n1227 ,n276 ,n878);
    nor g550(n1226 ,n395 ,n883);
    nor g551(n1225 ,n207 ,n881);
    nor g552(n1224 ,n284 ,n879);
    nor g553(n1223 ,n363 ,n880);
    nor g554(n1222 ,n344 ,n877);
    nor g555(n1221 ,n278 ,n882);
    nor g556(n1220 ,n189 ,n884);
    nor g557(n1219 ,n333 ,n875);
    nor g558(n1218 ,n367 ,n885);
    nor g559(n1217 ,n174 ,n878);
    nor g560(n1216 ,n382 ,n886);
    nor g561(n1215 ,n186 ,n883);
    nor g562(n1214 ,n341 ,n881);
    nor g563(n1213 ,n309 ,n878);
    nor g564(n1212 ,n353 ,n885);
    nor g565(n1211 ,n390 ,n875);
    nor g566(n1210 ,n214 ,n879);
    nor g567(n1209 ,n375 ,n886);
    nor g568(n1208 ,n335 ,n884);
    nor g569(n1207 ,n356 ,n882);
    nor g570(n1206 ,n211 ,n877);
    nor g571(n1205 ,n302 ,n876);
    nor g572(n1204 ,n205 ,n881);
    nor g573(n1203 ,n315 ,n879);
    nor g574(n1202 ,n387 ,n883);
    nor g575(n1201 ,n374 ,n875);
    nor g576(n1200 ,n379 ,n877);
    nor g577(n1199 ,n209 ,n882);
    nor g578(n1198 ,n385 ,n880);
    nor g579(n1197 ,n199 ,n876);
    nor g580(n1196 ,n285 ,n878);
    nor g581(n1195 ,n201 ,n885);
    nor g582(n1194 ,n217 ,n879);
    nor g583(n1193 ,n373 ,n886);
    nor g584(n1192 ,n301 ,n883);
    nor g585(n1191 ,n346 ,n878);
    nor g586(n1190 ,n191 ,n876);
    nor g587(n1189 ,n220 ,n875);
    nor g588(n1188 ,n298 ,n882);
    nor g589(n1187 ,n156 ,n885);
    nor g590(n1186 ,n136 ,n895);
    nor g591(n1321 ,n24[0] ,n894);
    or g592(n1320 ,n529 ,n887);
    nor g593(n1318 ,n467 ,n894);
    or g594(n1185 ,n1036 ,n761);
    nor g595(n1184 ,n126 ,n736);
    or g596(n1183 ,n947 ,n870);
    or g597(n1182 ,n1019 ,n1039);
    or g598(n1181 ,n1018 ,n1040);
    or g599(n1180 ,n1020 ,n1037);
    or g600(n1179 ,n1017 ,n1041);
    or g601(n1178 ,n1016 ,n1042);
    or g602(n1177 ,n1015 ,n874);
    or g603(n1176 ,n1014 ,n873);
    or g604(n1175 ,n1013 ,n872);
    or g605(n1174 ,n1012 ,n871);
    or g606(n1173 ,n1011 ,n869);
    or g607(n1172 ,n1010 ,n868);
    or g608(n1171 ,n1009 ,n864);
    or g609(n1170 ,n1008 ,n867);
    or g610(n1169 ,n1007 ,n866);
    or g611(n1168 ,n1005 ,n865);
    or g612(n1167 ,n1002 ,n1038);
    or g613(n1166 ,n1004 ,n863);
    or g614(n1165 ,n1003 ,n862);
    or g615(n1164 ,n1001 ,n861);
    or g616(n1163 ,n1000 ,n781);
    or g617(n1162 ,n999 ,n814);
    or g618(n1161 ,n998 ,n859);
    or g619(n1160 ,n995 ,n809);
    or g620(n1159 ,n996 ,n858);
    or g621(n1158 ,n994 ,n857);
    or g622(n1157 ,n733 ,n718);
    or g623(n1156 ,n993 ,n856);
    or g624(n1155 ,n939 ,n812);
    or g625(n1154 ,n997 ,n860);
    or g626(n1153 ,n988 ,n821);
    or g627(n1152 ,n992 ,n818);
    or g628(n1151 ,n991 ,n855);
    or g629(n1150 ,n989 ,n822);
    or g630(n1149 ,n1006 ,n819);
    or g631(n1148 ,n986 ,n854);
    or g632(n1147 ,n987 ,n853);
    or g633(n1146 ,n985 ,n852);
    or g634(n1145 ,n1028 ,n717);
    or g635(n1144 ,n984 ,n849);
    or g636(n1143 ,n948 ,n851);
    or g637(n1142 ,n983 ,n753);
    or g638(n1141 ,n981 ,n848);
    or g639(n1140 ,n951 ,n760);
    or g640(n1139 ,n980 ,n759);
    or g641(n1138 ,n979 ,n758);
    or g642(n1137 ,n978 ,n847);
    or g643(n1136 ,n977 ,n757);
    or g644(n1135 ,n976 ,n756);
    or g645(n1134 ,n958 ,n846);
    or g646(n1133 ,n957 ,n755);
    or g647(n1132 ,n975 ,n754);
    or g648(n1131 ,n973 ,n845);
    or g649(n1130 ,n974 ,n850);
    or g650(n1129 ,n972 ,n844);
    or g651(n1128 ,n971 ,n843);
    or g652(n1127 ,n969 ,n842);
    or g653(n1126 ,n968 ,n840);
    or g654(n1125 ,n982 ,n813);
    or g655(n1124 ,n967 ,n839);
    or g656(n1123 ,n966 ,n825);
    or g657(n1122 ,n965 ,n837);
    or g658(n1121 ,n963 ,n836);
    or g659(n1120 ,n962 ,n835);
    or g660(n1119 ,n1026 ,n716);
    or g661(n1118 ,n942 ,n834);
    or g662(n1117 ,n960 ,n832);
    or g663(n1116 ,n959 ,n786);
    or g664(n1115 ,n1027 ,n715);
    or g665(n1114 ,n938 ,n807);
    or g666(n1113 ,n911 ,n767);
    or g667(n1112 ,n956 ,n831);
    or g668(n1111 ,n955 ,n830);
    or g669(n1110 ,n954 ,n829);
    or g670(n1109 ,n712 ,n730);
    or g671(n1108 ,n934 ,n811);
    or g672(n1107 ,n952 ,n828);
    or g673(n1106 ,n950 ,n827);
    or g674(n1105 ,n943 ,n815);
    or g675(n1104 ,n923 ,n826);
    or g676(n1103 ,n946 ,n823);
    or g677(n1102 ,n953 ,n841);
    or g678(n1101 ,n945 ,n820);
    or g679(n1100 ,n711 ,n728);
    nor g680(n1099 ,n990 ,n1024);
    or g681(n1098 ,n944 ,n824);
    or g682(n1097 ,n713 ,n731);
    nor g683(n1096 ,n961 ,n1023);
    or g684(n1095 ,n940 ,n816);
    or g685(n1094 ,n970 ,n838);
    or g686(n1093 ,n949 ,n806);
    or g687(n1092 ,n1043 ,n810);
    or g688(n1091 ,n933 ,n833);
    nor g689(n1090 ,n936 ,n1025);
    or g690(n1089 ,n935 ,n794);
    or g691(n1088 ,n937 ,n808);
    nor g692(n1087 ,n932 ,n1022);
    or g693(n1086 ,n931 ,n805);
    or g694(n1085 ,n930 ,n804);
    or g695(n1084 ,n929 ,n803);
    nor g696(n1083 ,n927 ,n1021);
    or g697(n1082 ,n928 ,n802);
    or g698(n1081 ,n926 ,n801);
    or g699(n1080 ,n924 ,n799);
    or g700(n1079 ,n925 ,n800);
    or g701(n1078 ,n922 ,n798);
    or g702(n1077 ,n921 ,n797);
    or g703(n1076 ,n920 ,n796);
    or g704(n1075 ,n919 ,n795);
    or g705(n1074 ,n918 ,n793);
    or g706(n1073 ,n917 ,n792);
    or g707(n1072 ,n916 ,n791);
    or g708(n1071 ,n915 ,n790);
    or g709(n1070 ,n914 ,n789);
    or g710(n1069 ,n913 ,n788);
    or g711(n1068 ,n912 ,n787);
    or g712(n1067 ,n910 ,n785);
    or g713(n1066 ,n941 ,n817);
    or g714(n1065 ,n909 ,n784);
    or g715(n1064 ,n908 ,n783);
    or g716(n1063 ,n907 ,n782);
    or g717(n1062 ,n906 ,n780);
    or g718(n1061 ,n905 ,n779);
    or g719(n1060 ,n904 ,n778);
    or g720(n1059 ,n903 ,n777);
    or g721(n1058 ,n902 ,n776);
    or g722(n1057 ,n901 ,n775);
    or g723(n1056 ,n900 ,n774);
    or g724(n1055 ,n899 ,n773);
    or g725(n1054 ,n898 ,n772);
    or g726(n1053 ,n897 ,n771);
    or g727(n1052 ,n964 ,n770);
    or g728(n1051 ,n1029 ,n769);
    or g729(n1050 ,n1030 ,n768);
    or g730(n1049 ,n1031 ,n766);
    or g731(n1048 ,n1032 ,n765);
    or g732(n1047 ,n1033 ,n764);
    or g733(n1046 ,n1034 ,n763);
    or g734(n1045 ,n1035 ,n762);
    nor g735(n1044 ,n125 ,n752);
    nor g736(n1043 ,n341 ,n665);
    nor g737(n1042 ,n129 ,n654);
    nor g738(n1041 ,n132 ,n674);
    nor g739(n1040 ,n135 ,n674);
    nor g740(n1039 ,n134 ,n674);
    nor g741(n1038 ,n131 ,n656);
    nor g742(n1037 ,n133 ,n674);
    nor g743(n1036 ,n294 ,n675);
    nor g744(n1035 ,n198 ,n675);
    nor g745(n1034 ,n381 ,n675);
    nor g746(n1033 ,n168 ,n675);
    nor g747(n1032 ,n191 ,n671);
    nor g748(n1031 ,n199 ,n671);
    nor g749(n1030 ,n302 ,n671);
    nor g750(n1029 ,n299 ,n671);
    nor g751(n1028 ,n223 ,n688);
    nor g752(n1027 ,n232 ,n688);
    nor g753(n1026 ,n257 ,n688);
    nor g754(n1025 ,n237 ,n684);
    nor g755(n1024 ,n255 ,n684);
    nor g756(n1023 ,n246 ,n684);
    nor g757(n1022 ,n239 ,n684);
    nor g758(n1021 ,n229 ,n684);
    nor g759(n1020 ,n195 ,n675);
    nor g760(n1019 ,n314 ,n675);
    nor g761(n1018 ,n349 ,n675);
    nor g762(n1017 ,n210 ,n675);
    nor g763(n1016 ,n281 ,n655);
    nor g764(n1015 ,n166 ,n655);
    nor g765(n1014 ,n170 ,n655);
    nor g766(n1013 ,n178 ,n655);
    nor g767(n1012 ,n382 ,n655);
    nor g768(n1011 ,n375 ,n655);
    nor g769(n1010 ,n392 ,n655);
    nor g770(n1009 ,n155 ,n657);
    nor g771(n1008 ,n373 ,n655);
    nor g772(n1007 ,n293 ,n659);
    nor g773(n1006 ,n296 ,n669);
    nor g774(n1005 ,n200 ,n659);
    nor g775(n1004 ,n372 ,n659);
    nor g776(n1003 ,n395 ,n659);
    nor g777(n1002 ,n365 ,n657);
    nor g778(n1001 ,n387 ,n659);
    nor g779(n1000 ,n186 ,n659);
    nor g780(n999 ,n330 ,n657);
    nor g781(n998 ,n348 ,n659);
    nor g782(n997 ,n327 ,n669);
    nor g783(n996 ,n301 ,n659);
    nor g784(n995 ,n179 ,n657);
    nor g785(n994 ,n304 ,n661);
    nor g786(n993 ,n367 ,n657);
    nor g787(n992 ,n202 ,n661);
    nor g788(n991 ,n215 ,n661);
    nor g789(n990 ,n351 ,n685);
    nor g790(n989 ,n278 ,n661);
    nor g791(n988 ,n353 ,n657);
    nor g792(n987 ,n201 ,n657);
    nor g793(n986 ,n356 ,n661);
    nor g794(n985 ,n209 ,n661);
    nor g795(n984 ,n156 ,n657);
    nor g796(n983 ,n310 ,n653);
    nor g797(n982 ,n320 ,n673);
    nor g798(n981 ,n337 ,n667);
    nor g799(n980 ,n208 ,n653);
    nor g800(n979 ,n370 ,n653);
    nor g801(n978 ,n181 ,n667);
    nor g802(n977 ,n175 ,n653);
    nor g803(n976 ,n312 ,n653);
    nor g804(n975 ,n380 ,n653);
    nor g805(n974 ,n184 ,n669);
    nor g806(n973 ,n332 ,n667);
    nor g807(n972 ,n189 ,n667);
    nor g808(n971 ,n335 ,n667);
    nor g809(n970 ,n336 ,n665);
    nor g810(n969 ,n187 ,n667);
    nor g811(n968 ,n159 ,n667);
    nor g812(n967 ,n165 ,n663);
    nor g813(n966 ,n331 ,n681);
    nor g814(n965 ,n306 ,n663);
    nor g815(n964 ,n164 ,n671);
    nor g816(n963 ,n357 ,n663);
    nor g817(n962 ,n350 ,n663);
    nor g818(n961 ,n378 ,n685);
    nor g819(n960 ,n390 ,n663);
    nor g820(n959 ,n374 ,n663);
    nor g821(n958 ,n323 ,n667);
    nor g822(n957 ,n219 ,n653);
    nor g823(n956 ,n354 ,n681);
    nor g824(n955 ,n347 ,n681);
    nor g825(n954 ,n325 ,n681);
    nor g826(n953 ,n309 ,n669);
    nor g827(n952 ,n180 ,n681);
    nor g828(n951 ,n319 ,n653);
    nor g829(n950 ,n192 ,n681);
    nor g830(n949 ,n207 ,n665);
    nor g831(n948 ,n298 ,n661);
    nor g832(n947 ,n276 ,n669);
    nor g833(n946 ,n174 ,n669);
    nor g834(n945 ,n285 ,n669);
    nor g835(n944 ,n346 ,n669);
    nor g836(n943 ,n206 ,n665);
    nor g837(n942 ,n333 ,n663);
    nor g838(n941 ,n318 ,n665);
    nor g839(n940 ,n366 ,n665);
    nor g840(n939 ,n358 ,n661);
    nor g841(n938 ,n342 ,n673);
    nor g842(n937 ,n173 ,n665);
    nor g843(n936 ,n334 ,n685);
    nor g844(n935 ,n313 ,n673);
    nor g845(n934 ,n345 ,n681);
    nor g846(n933 ,n205 ,n665);
    nor g847(n932 ,n311 ,n685);
    nor g848(n931 ,n386 ,n673);
    nor g849(n930 ,n344 ,n673);
    nor g850(n929 ,n211 ,n673);
    nor g851(n928 ,n379 ,n673);
    nor g852(n927 ,n292 ,n685);
    nor g853(n926 ,n163 ,n673);
    nor g854(n925 ,n305 ,n677);
    nor g855(n924 ,n182 ,n677);
    nor g856(n923 ,n321 ,n681);
    nor g857(n922 ,n329 ,n677);
    nor g858(n921 ,n279 ,n677);
    nor g859(n920 ,n291 ,n677);
    nor g860(n919 ,n290 ,n677);
    nor g861(n918 ,n280 ,n677);
    nor g862(n917 ,n362 ,n677);
    nor g863(n916 ,n203 ,n679);
    nor g864(n915 ,n161 ,n679);
    nor g865(n914 ,n384 ,n679);
    nor g866(n913 ,n364 ,n679);
    nor g867(n912 ,n363 ,n679);
    nor g868(n911 ,n220 ,n663);
    nor g869(n910 ,n277 ,n679);
    nor g870(n909 ,n385 ,n679);
    nor g871(n908 ,n383 ,n679);
    nor g872(n907 ,n371 ,n683);
    nor g873(n906 ,n328 ,n683);
    nor g874(n905 ,n376 ,n683);
    nor g875(n904 ,n393 ,n683);
    nor g876(n903 ,n284 ,n683);
    nor g877(n902 ,n214 ,n683);
    nor g878(n901 ,n315 ,n683);
    nor g879(n900 ,n217 ,n683);
    nor g880(n899 ,n355 ,n671);
    nor g881(n898 ,n343 ,n671);
    nor g882(n897 ,n340 ,n671);
    not g883(n896 ,n895);
    not g884(n888 ,n887);
    nor g885(n874 ,n131 ,n654);
    nor g886(n873 ,n128 ,n654);
    nor g887(n872 ,n130 ,n654);
    nor g888(n871 ,n133 ,n654);
    nor g889(n870 ,n130 ,n668);
    nor g890(n869 ,n134 ,n654);
    nor g891(n868 ,n135 ,n654);
    nor g892(n867 ,n132 ,n654);
    nor g893(n866 ,n129 ,n658);
    nor g894(n865 ,n131 ,n658);
    nor g895(n864 ,n129 ,n656);
    nor g896(n863 ,n128 ,n658);
    nor g897(n862 ,n130 ,n658);
    nor g898(n861 ,n133 ,n658);
    nor g899(n860 ,n128 ,n668);
    nor g900(n859 ,n135 ,n658);
    nor g901(n858 ,n132 ,n658);
    nor g902(n857 ,n129 ,n660);
    nor g903(n856 ,n133 ,n656);
    nor g904(n855 ,n130 ,n660);
    nor g905(n854 ,n134 ,n660);
    nor g906(n853 ,n135 ,n656);
    nor g907(n852 ,n135 ,n660);
    nor g908(n851 ,n132 ,n660);
    nor g909(n850 ,n129 ,n668);
    nor g910(n849 ,n132 ,n656);
    nor g911(n848 ,n129 ,n666);
    nor g912(n847 ,n131 ,n666);
    nor g913(n846 ,n128 ,n666);
    nor g914(n845 ,n130 ,n666);
    nor g915(n844 ,n133 ,n666);
    nor g916(n843 ,n134 ,n666);
    nor g917(n842 ,n135 ,n666);
    nor g918(n841 ,n134 ,n668);
    nor g919(n840 ,n132 ,n666);
    nor g920(n839 ,n129 ,n662);
    nor g921(n838 ,n130 ,n664);
    nor g922(n837 ,n131 ,n662);
    nor g923(n836 ,n128 ,n662);
    nor g924(n835 ,n130 ,n662);
    nor g925(n834 ,n133 ,n662);
    nor g926(n833 ,n135 ,n664);
    nor g927(n832 ,n134 ,n662);
    nor g928(n831 ,n129 ,n680);
    nor g929(n830 ,n131 ,n680);
    nor g930(n829 ,n128 ,n680);
    nor g931(n828 ,n133 ,n680);
    nor g932(n827 ,n134 ,n680);
    nor g933(n826 ,n135 ,n680);
    nor g934(n825 ,n132 ,n680);
    nor g935(n824 ,n132 ,n668);
    nor g936(n823 ,n133 ,n668);
    nor g937(n822 ,n133 ,n660);
    nor g938(n821 ,n134 ,n656);
    nor g939(n820 ,n135 ,n668);
    nor g940(n819 ,n131 ,n668);
    nor g941(n818 ,n128 ,n660);
    nor g942(n817 ,n131 ,n664);
    nor g943(n816 ,n128 ,n664);
    nor g944(n815 ,n129 ,n664);
    nor g945(n814 ,n128 ,n656);
    nor g946(n813 ,n128 ,n672);
    nor g947(n812 ,n131 ,n660);
    nor g948(n811 ,n130 ,n680);
    nor g949(n810 ,n134 ,n664);
    nor g950(n809 ,n130 ,n656);
    nor g951(n808 ,n132 ,n664);
    nor g952(n807 ,n129 ,n672);
    nor g953(n806 ,n133 ,n664);
    nor g954(n805 ,n130 ,n672);
    nor g955(n804 ,n133 ,n672);
    nor g956(n803 ,n134 ,n672);
    nor g957(n802 ,n135 ,n672);
    nor g958(n801 ,n132 ,n672);
    nor g959(n800 ,n129 ,n676);
    nor g960(n799 ,n131 ,n676);
    nor g961(n798 ,n128 ,n676);
    nor g962(n797 ,n130 ,n676);
    nor g963(n796 ,n133 ,n676);
    nor g964(n795 ,n134 ,n676);
    nor g965(n794 ,n131 ,n672);
    nor g966(n793 ,n135 ,n676);
    nor g967(n792 ,n132 ,n676);
    nor g968(n791 ,n129 ,n678);
    nor g969(n790 ,n131 ,n678);
    nor g970(n789 ,n128 ,n678);
    nor g971(n788 ,n130 ,n678);
    nor g972(n787 ,n133 ,n678);
    nor g973(n786 ,n135 ,n662);
    nor g974(n785 ,n134 ,n678);
    nor g975(n784 ,n135 ,n678);
    nor g976(n783 ,n132 ,n678);
    nor g977(n782 ,n129 ,n682);
    nor g978(n781 ,n134 ,n658);
    nor g979(n780 ,n131 ,n682);
    nor g980(n779 ,n128 ,n682);
    nor g981(n778 ,n130 ,n682);
    nor g982(n777 ,n133 ,n682);
    nor g983(n776 ,n134 ,n682);
    nor g984(n775 ,n135 ,n682);
    nor g985(n774 ,n132 ,n682);
    nor g986(n773 ,n129 ,n670);
    nor g987(n772 ,n131 ,n670);
    nor g988(n771 ,n128 ,n670);
    nor g989(n770 ,n130 ,n670);
    nor g990(n769 ,n133 ,n670);
    nor g991(n768 ,n134 ,n670);
    nor g992(n767 ,n132 ,n662);
    nor g993(n766 ,n135 ,n670);
    nor g994(n765 ,n132 ,n670);
    nor g995(n764 ,n129 ,n674);
    nor g996(n763 ,n131 ,n674);
    nor g997(n762 ,n128 ,n674);
    nor g998(n761 ,n130 ,n674);
    nor g999(n760 ,n131 ,n652);
    nor g1000(n759 ,n128 ,n652);
    nor g1001(n758 ,n130 ,n652);
    nor g1002(n757 ,n133 ,n652);
    nor g1003(n756 ,n134 ,n652);
    nor g1004(n755 ,n135 ,n652);
    nor g1005(n754 ,n132 ,n652);
    nor g1006(n753 ,n129 ,n652);
    nor g1007(n752 ,n723 ,n694);
    or g1008(n751 ,n687 ,n587);
    nor g1009(n750 ,n724 ,n693);
    nor g1010(n749 ,n726 ,n695);
    nor g1011(n748 ,n565 ,n636);
    nor g1012(n747 ,n722 ,n696);
    nor g1013(n746 ,n692 ,n698);
    nor g1014(n745 ,n720 ,n699);
    or g1015(n744 ,n709 ,n704);
    or g1016(n743 ,n708 ,n701);
    nor g1017(n742 ,n562 ,n637);
    or g1018(n741 ,n710 ,n706);
    nor g1019(n740 ,n566 ,n651);
    nor g1020(n739 ,n536 ,n628);
    nor g1021(n738 ,n721 ,n697);
    nor g1022(n737 ,n569 ,n639);
    nor g1023(n736 ,n725 ,n700);
    or g1024(n735 ,n714 ,n705);
    nor g1025(n734 ,n634 ,n719);
    nor g1026(n733 ,n18[0] ,n688);
    nor g1027(n732 ,n127 ,n646);
    nor g1028(n731 ,n686 ,n614);
    nor g1029(n730 ,n686 ,n613);
    nor g1030(n729 ,n526 ,n686);
    nor g1031(n728 ,n686 ,n615);
    nor g1032(n895 ,n415 ,n685);
    or g1033(n894 ,n123 ,n684);
    or g1034(n893 ,n408 ,n686);
    or g1035(n892 ,n123 ,n685);
    or g1036(n890 ,n410 ,n686);
    or g1037(n889 ,n409 ,n686);
    nor g1038(n887 ,n407 ,n686);
    or g1039(n886 ,n407 ,n691);
    or g1040(n885 ,n408 ,n691);
    or g1041(n884 ,n408 ,n689);
    or g1042(n883 ,n407 ,n689);
    or g1043(n882 ,n407 ,n690);
    or g1044(n881 ,n409 ,n689);
    or g1045(n880 ,n410 ,n691);
    or g1046(n879 ,n410 ,n689);
    or g1047(n878 ,n409 ,n691);
    or g1048(n877 ,n409 ,n690);
    or g1049(n876 ,n410 ,n690);
    or g1050(n875 ,n408 ,n690);
    nor g1051(n727 ,n185 ,n593);
    nor g1052(n726 ,n148 ,n620);
    nor g1053(n725 ,n274 ,n620);
    nor g1054(n724 ,n144 ,n620);
    nor g1055(n723 ,n142 ,n620);
    nor g1056(n722 ,n265 ,n620);
    nor g1057(n721 ,n145 ,n620);
    nor g1058(n720 ,n269 ,n620);
    nor g1059(n719 ,n324 ,n601);
    nor g1060(n718 ,n272 ,n597);
    nor g1061(n717 ,n150 ,n597);
    nor g1062(n716 ,n151 ,n597);
    nor g1063(n715 ,n152 ,n597);
    nor g1064(n714 ,n297 ,n594);
    nor g1065(n713 ,n160 ,n594);
    nor g1066(n712 ,n185 ,n594);
    nor g1067(n711 ,n288 ,n594);
    nor g1068(n710 ,n295 ,n594);
    nor g1069(n709 ,n326 ,n594);
    nor g1070(n708 ,n283 ,n594);
    nor g1071(n707 ,n295 ,n593);
    nor g1072(n706 ,n297 ,n593);
    nor g1073(n705 ,n288 ,n593);
    nor g1074(n704 ,n283 ,n593);
    nor g1075(n703 ,n326 ,n593);
    nor g1076(n702 ,n160 ,n593);
    nor g1077(n701 ,n316 ,n593);
    nor g1078(n700 ,n144 ,n619);
    nor g1079(n699 ,n1516 ,n619);
    nor g1080(n698 ,n269 ,n619);
    nor g1081(n697 ,n268 ,n619);
    nor g1082(n696 ,n145 ,n619);
    nor g1083(n695 ,n265 ,n619);
    nor g1084(n694 ,n148 ,n619);
    nor g1085(n693 ,n142 ,n619);
    nor g1086(n692 ,n268 ,n620);
    not g1087(n688 ,n687);
    not g1088(n684 ,n685);
    not g1089(n682 ,n683);
    not g1090(n680 ,n681);
    not g1091(n678 ,n679);
    not g1092(n676 ,n677);
    not g1093(n674 ,n675);
    not g1094(n672 ,n673);
    not g1095(n670 ,n671);
    not g1096(n668 ,n669);
    not g1097(n666 ,n667);
    not g1098(n664 ,n665);
    not g1099(n662 ,n663);
    not g1100(n660 ,n661);
    not g1101(n658 ,n659);
    not g1102(n656 ,n657);
    not g1103(n654 ,n655);
    not g1104(n652 ,n653);
    nor g1105(n651 ,n17[0] ,n622);
    or g1106(n650 ,n455 ,n607);
    or g1107(n649 ,n475 ,n611);
    or g1108(n648 ,n474 ,n608);
    or g1109(n647 ,n472 ,n610);
    nor g1110(n646 ,n604 ,n609);
    or g1111(n645 ,n605 ,n598);
    nor g1112(n644 ,n126 ,n572);
    nor g1113(n643 ,n127 ,n586);
    nor g1114(n642 ,n125 ,n571);
    nor g1115(n641 ,n126 ,n573);
    nor g1116(n640 ,n127 ,n574);
    nor g1117(n639 ,n17[1] ,n622);
    or g1118(n638 ,n621 ,n528);
    nor g1119(n637 ,n17[3] ,n622);
    nor g1120(n636 ,n17[2] ,n622);
    or g1121(n635 ,n549 ,n589);
    nor g1122(n634 ,n136 ,n600);
    or g1123(n633 ,n547 ,n588);
    or g1124(n632 ,n559 ,n592);
    or g1125(n631 ,n556 ,n576);
    or g1126(n630 ,n554 ,n577);
    or g1127(n629 ,n550 ,n591);
    nor g1128(n628 ,n496 ,n575);
    or g1129(n627 ,n551 ,n585);
    or g1130(n626 ,n546 ,n590);
    or g1131(n691 ,n44[1] ,n599);
    or g1132(n690 ,n138 ,n599);
    or g1133(n689 ,n44[1] ,n625);
    nor g1134(n687 ,n123 ,n619);
    or g1135(n686 ,n138 ,n625);
    nor g1136(n685 ,n470 ,n619);
    nor g1137(n683 ,n413 ,n623);
    nor g1138(n681 ,n412 ,n624);
    nor g1139(n679 ,n413 ,n595);
    nor g1140(n677 ,n414 ,n624);
    nor g1141(n675 ,n412 ,n623);
    nor g1142(n673 ,n414 ,n596);
    nor g1143(n671 ,n412 ,n595);
    nor g1144(n669 ,n411 ,n596);
    nor g1145(n667 ,n413 ,n624);
    nor g1146(n665 ,n411 ,n624);
    nor g1147(n663 ,n412 ,n596);
    nor g1148(n661 ,n414 ,n595);
    nor g1149(n659 ,n411 ,n623);
    nor g1150(n657 ,n413 ,n596);
    nor g1151(n655 ,n411 ,n595);
    nor g1152(n653 ,n414 ,n623);
    not g1153(n622 ,n621);
    not g1154(n619 ,n620);
    nor g1155(n618 ,n127 ,n518);
    nor g1156(n617 ,n124 ,n519);
    nor g1157(n616 ,n124 ,n568);
    nor g1158(n615 ,n504 ,n503);
    nor g1159(n614 ,n499 ,n508);
    nor g1160(n613 ,n517 ,n516);
    nor g1161(n612 ,n262 ,n527);
    nor g1162(n611 ,n227 ,n532);
    nor g1163(n610 ,n245 ,n532);
    nor g1164(n609 ,n316 ,n531);
    nor g1165(n608 ,n254 ,n532);
    nor g1166(n607 ,n248 ,n532);
    nor g1167(n606 ,n1517 ,n515);
    nor g1168(n605 ,n271 ,n527);
    nor g1169(n604 ,n158 ,n530);
    nor g1170(n603 ,n138 ,n527);
    nor g1171(n602 ,n264 ,n527);
    or g1172(n625 ,n271 ,n529);
    or g1173(n624 ,n141 ,n533);
    or g1174(n623 ,n141 ,n570);
    nor g1175(n621 ,n136 ,n536);
    nor g1176(n620 ,n136 ,n535);
    not g1177(n601 ,n600);
    not g1178(n599 ,n598);
    or g1179(n592 ,n480 ,n558);
    or g1180(n591 ,n450 ,n552);
    or g1181(n590 ,n478 ,n545);
    or g1182(n589 ,n451 ,n548);
    or g1183(n588 ,n452 ,n560);
    nor g1184(n587 ,n462 ,n561);
    nor g1185(n586 ,n539 ,n540);
    or g1186(n585 ,n497 ,n557);
    nor g1187(n584 ,n124 ,n502);
    nor g1188(n583 ,n124 ,n501);
    nor g1189(n582 ,n127 ,n500);
    nor g1190(n581 ,n126 ,n512);
    nor g1191(n580 ,n125 ,n514);
    nor g1192(n579 ,n123 ,n509);
    nor g1193(n578 ,n126 ,n567);
    or g1194(n577 ,n481 ,n555);
    or g1195(n576 ,n454 ,n553);
    or g1196(n575 ,n26[0] ,n520);
    nor g1197(n574 ,n563 ,n544);
    nor g1198(n573 ,n537 ,n543);
    nor g1199(n572 ,n521 ,n541);
    nor g1200(n571 ,n538 ,n542);
    nor g1201(n600 ,n415 ,n522);
    nor g1202(n598 ,n44[0] ,n529);
    or g1203(n597 ,n461 ,n534);
    or g1204(n596 ,n45[0] ,n533);
    or g1205(n595 ,n45[0] ,n570);
    or g1206(n594 ,n124 ,n531);
    or g1207(n593 ,n527 ,n530);
    nor g1208(n569 ,n234 ,n460);
    or g1209(n568 ,n197 ,n465);
    or g1210(n567 ,n153 ,n471);
    nor g1211(n566 ,n250 ,n460);
    nor g1212(n565 ,n258 ,n460);
    nor g1213(n564 ,n154 ,n459);
    nor g1214(n563 ,n389 ,n457);
    nor g1215(n562 ,n221 ,n460);
    or g1216(n561 ,n146 ,n461);
    nor g1217(n560 ,n194 ,n458);
    nor g1218(n559 ,n287 ,n498);
    nor g1219(n558 ,n303 ,n458);
    nor g1220(n557 ,n218 ,n498);
    nor g1221(n556 ,n286 ,n458);
    nor g1222(n555 ,n369 ,n458);
    nor g1223(n554 ,n396 ,n498);
    nor g1224(n553 ,n394 ,n498);
    nor g1225(n552 ,n213 ,n458);
    nor g1226(n551 ,n307 ,n458);
    nor g1227(n550 ,n177 ,n498);
    nor g1228(n549 ,n308 ,n458);
    nor g1229(n548 ,n167 ,n498);
    nor g1230(n547 ,n391 ,n498);
    nor g1231(n546 ,n322 ,n498);
    nor g1232(n545 ,n388 ,n458);
    nor g1233(n544 ,n252 ,n456);
    nor g1234(n543 ,n228 ,n456);
    nor g1235(n542 ,n253 ,n456);
    nor g1236(n541 ,n240 ,n456);
    nor g1237(n540 ,n236 ,n456);
    nor g1238(n539 ,n338 ,n457);
    nor g1239(n538 ,n275 ,n457);
    nor g1240(n537 ,n162 ,n457);
    or g1241(n570 ,n154 ,n464);
    not g1242(n535 ,n534);
    not g1243(n531 ,n530);
    not g1244(n529 ,n528);
    nor g1245(n526 ,n489 ,n488);
    nor g1246(n525 ,n141 ,n459);
    nor g1247(n524 ,n139 ,n459);
    nor g1248(n523 ,n140 ,n459);
    nor g1249(n522 ,n136 ,n469);
    nor g1250(n521 ,n216 ,n457);
    nor g1251(n520 ,n439 ,n470);
    or g1252(n519 ,n22[4] ,n465);
    or g1253(n518 ,n43[4] ,n471);
    or g1254(n517 ,n484 ,n494);
    or g1255(n516 ,n491 ,n485);
    nor g1256(n514 ,n423 ,n438);
    nor g1257(n513 ,n19[0] ,n461);
    nor g1258(n512 ,n447 ,n476);
    nor g1259(n511 ,n123 ,n441);
    nor g1260(n510 ,n123 ,n440);
    nor g1261(n509 ,n446 ,n473);
    or g1262(n508 ,n486 ,n483);
    nor g1263(n507 ,n123 ,n444);
    nor g1264(n506 ,n123 ,n442);
    nor g1265(n505 ,n124 ,n443);
    or g1266(n504 ,n482 ,n492);
    or g1267(n503 ,n490 ,n487);
    nor g1268(n502 ,n449 ,n453);
    nor g1269(n501 ,n448 ,n477);
    nor g1270(n500 ,n445 ,n479);
    or g1271(n499 ,n495 ,n493);
    or g1272(n536 ,n124 ,n468);
    nor g1273(n534 ,n15 ,n463);
    or g1274(n533 ,n45[3] ,n464);
    nor g1275(n530 ,n424 ,n463);
    nor g1276(n528 ,n125 ,n456);
    or g1277(n527 ,n123 ,n457);
    nor g1278(n497 ,n282 ,n406);
    nor g1279(n496 ,n1518 ,n420);
    nor g1280(n495 ,n314 ,n410);
    nor g1281(n494 ,n182 ,n409);
    nor g1282(n493 ,n290 ,n409);
    nor g1283(n492 ,n291 ,n409);
    nor g1284(n491 ,n381 ,n410);
    nor g1285(n490 ,n195 ,n410);
    nor g1286(n489 ,n370 ,n407);
    nor g1287(n488 ,n345 ,n408);
    nor g1288(n487 ,n180 ,n408);
    nor g1289(n486 ,n312 ,n407);
    nor g1290(n485 ,n347 ,n408);
    nor g1291(n484 ,n319 ,n407);
    nor g1292(n483 ,n192 ,n408);
    nor g1293(n482 ,n175 ,n407);
    nor g1294(n481 ,n377 ,n406);
    nor g1295(n480 ,n289 ,n406);
    nor g1296(n479 ,n243 ,n434);
    nor g1297(n478 ,n359 ,n406);
    nor g1298(n477 ,n247 ,n434);
    nor g1299(n476 ,n251 ,n434);
    nor g1300(n475 ,n193 ,n406);
    nor g1301(n474 ,n188 ,n406);
    nor g1302(n473 ,n261 ,n434);
    nor g1303(n472 ,n183 ,n406);
    or g1304(n498 ,n147 ,n416);
    not g1305(n469 ,n468);
    not g1306(n467 ,n466);
    not g1307(n463 ,n462);
    not g1308(n456 ,n457);
    nor g1309(n455 ,n147 ,n406);
    nor g1310(n454 ,n352 ,n406);
    nor g1311(n453 ,n226 ,n434);
    nor g1312(n452 ,n212 ,n406);
    nor g1313(n451 ,n204 ,n406);
    nor g1314(n450 ,n190 ,n406);
    nor g1315(n449 ,n300 ,n435);
    nor g1316(n448 ,n339 ,n435);
    nor g1317(n447 ,n172 ,n435);
    nor g1318(n445 ,n361 ,n435);
    nor g1319(n444 ,n428 ,n419);
    nor g1320(n443 ,n427 ,n404);
    nor g1321(n442 ,n425 ,n397);
    nor g1322(n441 ,n426 ,n431);
    nor g1323(n440 ,n429 ,n421);
    or g1324(n439 ,n136 ,n437);
    or g1325(n471 ,n400 ,n399);
    or g1326(n470 ,n430 ,n418);
    nor g1327(n468 ,n263 ,n437);
    nor g1328(n466 ,n432 ,n433);
    or g1329(n465 ,n401 ,n398);
    or g1330(n464 ,n124 ,n434);
    nor g1331(n462 ,n26[0] ,n437);
    or g1332(n461 ,n123 ,n415);
    or g1333(n460 ,n124 ,n417);
    or g1334(n459 ,n124 ,n435);
    or g1335(n458 ,n23[3] ,n416);
    nor g1336(n457 ,n437 ,n417);
    not g1337(n437 ,n436);
    not g1338(n434 ,n435);
    or g1339(n433 ,n270 ,n267);
    or g1340(n432 ,n143 ,n266);
    nor g1341(n431 ,n317 ,n1548);
    or g1342(n430 ,n272 ,n150);
    nor g1343(n429 ,n137 ,n222);
    nor g1344(n428 ,n137 ,n238);
    nor g1345(n427 ,n137 ,n249);
    nor g1346(n426 ,n137 ,n260);
    nor g1347(n425 ,n137 ,n241);
    or g1348(n424 ,n146 ,n136);
    nor g1349(n423 ,n273 ,n136);
    nor g1350(n422 ,n273 ,n126);
    nor g1351(n421 ,n169 ,n1548);
    or g1352(n420 ,n196 ,n26[1]);
    nor g1353(n419 ,n368 ,n1548);
    or g1354(n418 ,n151 ,n18[3]);
    nor g1355(n436 ,n149 ,n157);
    nor g1356(n435 ,n196 ,n43[4]);
    nor g1357(n405 ,n136 ,n123);
    nor g1358(n404 ,n176 ,n1548);
    or g1359(n403 ,n24[1] ,n24[2]);
    nor g1360(n402 ,n263 ,n123);
    or g1361(n401 ,n22[0] ,n22[3]);
    or g1362(n400 ,n43[0] ,n43[3]);
    or g1363(n399 ,n43[2] ,n43[1]);
    or g1364(n398 ,n22[2] ,n22[1]);
    nor g1365(n397 ,n171 ,n1548);
    or g1366(n417 ,n263 ,n26[1]);
    or g1367(n416 ,n124 ,n137);
    nor g1368(n415 ,n26[0] ,n26[1]);
    or g1369(n414 ,n140 ,n139);
    or g1370(n413 ,n45[2] ,n45[1]);
    or g1371(n412 ,n139 ,n45[2]);
    or g1372(n411 ,n140 ,n45[1]);
    or g1373(n410 ,n264 ,n44[2]);
    or g1374(n409 ,n262 ,n44[3]);
    or g1375(n408 ,n44[2] ,n44[3]);
    or g1376(n407 ,n262 ,n264);
    or g1377(n406 ,n124 ,n1548);
    not g1378(n396 ,n21[6]);
    not g1379(n395 ,n40[3]);
    not g1380(n394 ,n21[7]);
    not g1381(n393 ,n36[3]);
    not g1382(n392 ,n39[6]);
    not g1383(n391 ,n21[1]);
    not g1384(n390 ,n29[5]);
    not g1385(n389 ,n43[0]);
    not g1386(n388 ,n20[2]);
    not g1387(n387 ,n40[4]);
    not g1388(n386 ,n33[3]);
    not g1389(n385 ,n35[6]);
    not g1390(n384 ,n35[2]);
    not g1391(n383 ,n35[7]);
    not g1392(n382 ,n39[4]);
    not g1393(n381 ,n38[1]);
    not g1394(n380 ,n42[7]);
    not g1395(n379 ,n33[6]);
    not g1396(n378 ,n22[1]);
    not g1397(n377 ,n6[6]);
    not g1398(n376 ,n36[2]);
    not g1399(n375 ,n39[5]);
    not g1400(n374 ,n29[6]);
    not g1401(n373 ,n39[7]);
    not g1402(n372 ,n40[2]);
    not g1403(n371 ,n36[0]);
    not g1404(n370 ,n42[3]);
    not g1405(n369 ,n20[6]);
    not g1406(n368 ,n22[0]);
    not g1407(n367 ,n27[4]);
    not g1408(n366 ,n32[2]);
    not g1409(n365 ,n27[1]);
    not g1410(n364 ,n35[3]);
    not g1411(n363 ,n35[4]);
    not g1412(n362 ,n34[7]);
    not g1413(n361 ,n43[3]);
    not g1414(n360 ,n12);
    not g1415(n359 ,n6[2]);
    not g1416(n358 ,n41[1]);
    not g1417(n357 ,n29[2]);
    not g1418(n356 ,n41[5]);
    not g1419(n355 ,n37[0]);
    not g1420(n354 ,n30[0]);
    not g1421(n353 ,n27[5]);
    not g1422(n352 ,n6[7]);
    not g1423(n351 ,n22[0]);
    not g1424(n350 ,n29[3]);
    not g1425(n349 ,n38[6]);
    not g1426(n348 ,n40[6]);
    not g1427(n347 ,n30[1]);
    not g1428(n346 ,n31[7]);
    not g1429(n345 ,n30[3]);
    not g1430(n344 ,n33[4]);
    not g1431(n343 ,n37[1]);
    not g1432(n342 ,n33[0]);
    not g1433(n341 ,n32[5]);
    not g1434(n340 ,n37[2]);
    not g1435(n339 ,n43[2]);
    not g1436(n338 ,n43[3]);
    not g1437(n337 ,n28[0]);
    not g1438(n336 ,n32[3]);
    not g1439(n335 ,n28[5]);
    not g1440(n334 ,n22[2]);
    not g1441(n333 ,n29[4]);
    not g1442(n332 ,n28[3]);
    not g1443(n331 ,n30[7]);
    not g1444(n330 ,n27[2]);
    not g1445(n329 ,n34[2]);
    not g1446(n328 ,n36[1]);
    not g1447(n327 ,n31[2]);
    not g1448(n326 ,n46[5]);
    not g1449(n325 ,n30[2]);
    not g1450(n324 ,n11);
    not g1451(n323 ,n28[2]);
    not g1452(n322 ,n21[2]);
    not g1453(n321 ,n30[6]);
    not g1454(n320 ,n33[2]);
    not g1455(n319 ,n42[1]);
    not g1456(n318 ,n32[1]);
    not g1457(n317 ,n22[1]);
    not g1458(n316 ,n46[7]);
    not g1459(n315 ,n36[6]);
    not g1460(n314 ,n38[5]);
    not g1461(n313 ,n33[1]);
    not g1462(n312 ,n42[5]);
    not g1463(n311 ,n22[3]);
    not g1464(n310 ,n42[0]);
    not g1465(n309 ,n31[5]);
    not g1466(n308 ,n20[3]);
    not g1467(n307 ,n20[0]);
    not g1468(n306 ,n29[1]);
    not g1469(n305 ,n34[0]);
    not g1470(n304 ,n41[0]);
    not g1471(n303 ,n20[5]);
    not g1472(n302 ,n37[5]);
    not g1473(n301 ,n40[7]);
    not g1474(n300 ,n43[1]);
    not g1475(n299 ,n37[4]);
    not g1476(n298 ,n41[7]);
    not g1477(n297 ,n46[2]);
    not g1478(n296 ,n31[1]);
    not g1479(n295 ,n46[1]);
    not g1480(n294 ,n38[3]);
    not g1481(n293 ,n40[0]);
    not g1482(n292 ,n22[4]);
    not g1483(n291 ,n34[4]);
    not g1484(n290 ,n34[5]);
    not g1485(n289 ,n6[5]);
    not g1486(n288 ,n46[3]);
    not g1487(n287 ,n21[5]);
    not g1488(n286 ,n20[7]);
    not g1489(n285 ,n31[6]);
    not g1490(n284 ,n36[4]);
    not g1491(n283 ,n46[6]);
    not g1492(n282 ,n6[0]);
    not g1493(n281 ,n39[0]);
    not g1494(n280 ,n34[6]);
    not g1495(n279 ,n34[3]);
    not g1496(n278 ,n41[4]);
    not g1497(n277 ,n35[5]);
    not g1498(n276 ,n31[3]);
    not g1499(n275 ,n43[2]);
    not g1500(n274 ,n25[7]);
    not g1501(n273 ,n13);
    not g1502(n272 ,n18[0]);
    not g1503(n271 ,n44[0]);
    not g1504(n270 ,n24[2]);
    not g1505(n269 ,n25[0]);
    not g1506(n268 ,n25[1]);
    not g1507(n267 ,n24[3]);
    not g1508(n266 ,n24[1]);
    not g1509(n265 ,n25[3]);
    not g1510(n264 ,n44[3]);
    not g1511(n263 ,n26[0]);
    not g1512(n262 ,n44[2]);
    not g1513(n261 ,n1554);
    not g1514(n260 ,n1541);
    not g1515(n259 ,n1524);
    not g1516(n258 ,n5[2]);
    not g1517(n257 ,n1535);
    not g1518(n256 ,n1521);
    not g1519(n255 ,n1553);
    not g1520(n254 ,n1530);
    not g1521(n253 ,n1545);
    not g1522(n252 ,n1547);
    not g1523(n251 ,n1558);
    not g1524(n250 ,n5[0]);
    not g1525(n249 ,n1538);
    not g1526(n248 ,n1532);
    not g1527(n247 ,n1556);
    not g1528(n246 ,n1552);
    not g1529(n245 ,n1529);
    not g1530(n244 ,n1519);
    not g1531(n243 ,n1555);
    not g1532(n242 ,n1522);
    not g1533(n241 ,n1539);
    not g1534(n240 ,n1543);
    not g1535(n239 ,n1550);
    not g1536(n238 ,n1542);
    not g1537(n237 ,n1551);
    not g1538(n236 ,n1544);
    not g1539(n235 ,n1523);
    not g1540(n234 ,n5[1]);
    not g1541(n233 ,n1528);
    not g1542(n232 ,n1536);
    not g1543(n231 ,n1525);
    not g1544(n230 ,n1520);
    not g1545(n229 ,n1549);
    not g1546(n228 ,n1546);
    not g1547(n227 ,n1531);
    not g1548(n226 ,n1557);
    not g1549(n225 ,n1526);
    not g1550(n224 ,n1527);
    not g1551(n223 ,n1534);
    not g1552(n222 ,n1540);
    not g1553(n221 ,n5[3]);
    not g1554(n220 ,n29[7]);
    not g1555(n219 ,n42[6]);
    not g1556(n218 ,n21[0]);
    not g1557(n217 ,n36[7]);
    not g1558(n216 ,n43[4]);
    not g1559(n215 ,n41[3]);
    not g1560(n214 ,n36[5]);
    not g1561(n213 ,n20[4]);
    not g1562(n212 ,n6[1]);
    not g1563(n211 ,n33[5]);
    not g1564(n210 ,n38[7]);
    not g1565(n209 ,n41[6]);
    not g1566(n208 ,n42[2]);
    not g1567(n207 ,n32[4]);
    not g1568(n206 ,n32[0]);
    not g1569(n205 ,n32[6]);
    not g1570(n204 ,n6[3]);
    not g1571(n203 ,n35[0]);
    not g1572(n202 ,n41[2]);
    not g1573(n201 ,n27[6]);
    not g1574(n200 ,n40[1]);
    not g1575(n199 ,n37[6]);
    not g1576(n198 ,n38[2]);
    not g1577(n197 ,n22[4]);
    not g1578(n196 ,n2);
    not g1579(n195 ,n38[4]);
    not g1580(n194 ,n20[1]);
    not g1581(n193 ,n23[2]);
    not g1582(n192 ,n30[5]);
    not g1583(n191 ,n37[7]);
    not g1584(n190 ,n6[4]);
    not g1585(n189 ,n28[4]);
    not g1586(n188 ,n23[1]);
    not g1587(n187 ,n28[6]);
    not g1588(n186 ,n40[5]);
    not g1589(n185 ,n46[0]);
    not g1590(n184 ,n31[0]);
    not g1591(n183 ,n23[0]);
    not g1592(n182 ,n34[1]);
    not g1593(n181 ,n28[1]);
    not g1594(n180 ,n30[4]);
    not g1595(n179 ,n27[3]);
    not g1596(n178 ,n39[3]);
    not g1597(n177 ,n21[4]);
    not g1598(n176 ,n22[4]);
    not g1599(n175 ,n42[4]);
    not g1600(n174 ,n31[4]);
    not g1601(n173 ,n32[7]);
    not g1602(n172 ,n43[0]);
    not g1603(n171 ,n22[3]);
    not g1604(n170 ,n39[2]);
    not g1605(n169 ,n22[2]);
    not g1606(n168 ,n38[0]);
    not g1607(n167 ,n21[3]);
    not g1608(n166 ,n39[1]);
    not g1609(n165 ,n29[0]);
    not g1610(n164 ,n37[3]);
    not g1611(n163 ,n33[7]);
    not g1612(n162 ,n43[1]);
    not g1613(n161 ,n35[1]);
    not g1614(n160 ,n46[4]);
    not g1615(n159 ,n28[7]);
    not g1616(n158 ,n16);
    not g1617(n157 ,n19[1]);
    not g1618(n156 ,n27[7]);
    not g1619(n155 ,n27[0]);
    not g1620(n154 ,n45[3]);
    not g1621(n153 ,n43[4]);
    not g1622(n152 ,n18[3]);
    not g1623(n151 ,n18[2]);
    not g1624(n150 ,n18[1]);
    not g1625(n149 ,n19[0]);
    not g1626(n148 ,n25[4]);
    not g1627(n147 ,n23[3]);
    not g1628(n146 ,n15);
    not g1629(n145 ,n25[2]);
    not g1630(n144 ,n25[6]);
    not g1631(n143 ,n24[0]);
    not g1632(n142 ,n25[5]);
    not g1633(n141 ,n45[0]);
    not g1634(n140 ,n45[2]);
    not g1635(n139 ,n45[1]);
    not g1636(n138 ,n44[1]);
    not g1637(n137 ,n1548);
    not g1638(n136 ,n26[1]);
    not g1639(n135 ,n4[6]);
    not g1640(n134 ,n4[5]);
    not g1641(n133 ,n4[4]);
    not g1642(n132 ,n4[7]);
    not g1643(n131 ,n4[1]);
    not g1644(n130 ,n4[3]);
    not g1645(n129 ,n4[0]);
    not g1646(n128 ,n4[2]);
    not g1647(n127 ,n1);
    not g1648(n126 ,n1);
    not g1649(n125 ,n1);
    not g1650(n124 ,n1);
    not g1651(n123 ,n1);
    xor g1652(n1543 ,n43[4] ,n51);
    xor g1653(n1544 ,n43[3] ,n49);
    nor g1654(n51 ,n43[3] ,n50);
    xor g1655(n1545 ,n43[2] ,n47);
    not g1656(n50 ,n49);
    nor g1657(n49 ,n43[2] ,n48);
    xnor g1658(n1546 ,n43[1] ,n43[0]);
    not g1659(n48 ,n47);
    nor g1660(n47 ,n43[1] ,n43[0]);
    not g1661(n1547 ,n43[0]);
    xor g1662(n1538 ,n22[4] ,n56);
    xor g1663(n1539 ,n22[3] ,n54);
    nor g1664(n56 ,n22[3] ,n55);
    xor g1665(n1540 ,n22[2] ,n52);
    not g1666(n55 ,n54);
    nor g1667(n54 ,n22[2] ,n53);
    xnor g1668(n1541 ,n22[1] ,n22[0]);
    not g1669(n53 ,n52);
    nor g1670(n52 ,n22[1] ,n22[0]);
    not g1671(n1542 ,n22[0]);
    or g1672(n1537 ,n58 ,n59);
    or g1673(n59 ,n43[3] ,n57);
    or g1674(n58 ,n43[2] ,n43[0]);
    or g1675(n57 ,n43[4] ,n43[1]);
    or g1676(n1548 ,n61 ,n62);
    or g1677(n62 ,n22[3] ,n60);
    or g1678(n61 ,n22[2] ,n22[0]);
    or g1679(n60 ,n22[4] ,n22[1]);
    xor g1680(n1521 ,n44[3] ,n70);
    nor g1681(n1520 ,n69 ,n70);
    nor g1682(n70 ,n65 ,n68);
    nor g1683(n69 ,n44[2] ,n67);
    nor g1684(n1519 ,n67 ,n66);
    not g1685(n68 ,n67);
    nor g1686(n67 ,n63 ,n64);
    nor g1687(n66 ,n44[1] ,n44[0]);
    not g1688(n65 ,n44[2]);
    not g1689(n64 ,n44[0]);
    not g1690(n63 ,n44[1]);
    xor g1691(n1533 ,n19[1] ,n19[0]);
    xor g1692(n1524 ,n24[3] ,n78);
    nor g1693(n1523 ,n77 ,n78);
    nor g1694(n78 ,n73 ,n76);
    nor g1695(n77 ,n24[2] ,n75);
    nor g1696(n1522 ,n75 ,n74);
    not g1697(n76 ,n75);
    nor g1698(n75 ,n71 ,n72);
    nor g1699(n74 ,n24[1] ,n24[0]);
    not g1700(n73 ,n24[2]);
    not g1701(n72 ,n24[0]);
    not g1702(n71 ,n24[1]);
    xor g1703(n1549 ,n22[4] ,n89);
    nor g1704(n1550 ,n88 ,n89);
    nor g1705(n89 ,n80 ,n87);
    nor g1706(n88 ,n22[3] ,n86);
    nor g1707(n1551 ,n85 ,n86);
    not g1708(n87 ,n86);
    nor g1709(n86 ,n81 ,n84);
    nor g1710(n85 ,n22[2] ,n83);
    nor g1711(n1552 ,n83 ,n82);
    not g1712(n84 ,n83);
    nor g1713(n83 ,n79 ,n1553);
    nor g1714(n82 ,n22[1] ,n22[0]);
    not g1715(n81 ,n22[2]);
    not g1716(n1553 ,n22[0]);
    not g1717(n80 ,n22[3]);
    not g1718(n79 ,n22[1]);
    xor g1719(n1536 ,n18[3] ,n97);
    nor g1720(n1535 ,n96 ,n97);
    nor g1721(n97 ,n92 ,n95);
    nor g1722(n96 ,n18[2] ,n94);
    nor g1723(n1534 ,n94 ,n93);
    not g1724(n95 ,n94);
    nor g1725(n94 ,n90 ,n91);
    nor g1726(n93 ,n18[1] ,n18[0]);
    not g1727(n92 ,n18[2]);
    not g1728(n91 ,n18[0]);
    not g1729(n90 ,n18[1]);
    xor g1730(n1528 ,n104 ,n45[3]);
    nor g1731(n1527 ,n103 ,n104);
    nor g1732(n104 ,n99 ,n102);
    nor g1733(n103 ,n45[2] ,n101);
    nor g1734(n1526 ,n101 ,n100);
    not g1735(n102 ,n101);
    nor g1736(n101 ,n98 ,n1525);
    nor g1737(n100 ,n45[1] ,n45[0]);
    not g1738(n99 ,n45[2]);
    not g1739(n1525 ,n45[0]);
    not g1740(n98 ,n45[1]);
    nor g1741(n1555 ,n114 ,n115);
    nor g1742(n115 ,n106 ,n113);
    nor g1743(n114 ,n43[3] ,n112);
    nor g1744(n1556 ,n111 ,n112);
    not g1745(n113 ,n112);
    nor g1746(n112 ,n107 ,n110);
    nor g1747(n111 ,n43[2] ,n109);
    nor g1748(n1557 ,n109 ,n108);
    not g1749(n110 ,n109);
    nor g1750(n109 ,n105 ,n1558);
    nor g1751(n108 ,n43[1] ,n43[0]);
    not g1752(n107 ,n43[2]);
    not g1753(n1558 ,n43[0]);
    not g1754(n106 ,n43[3]);
    not g1755(n105 ,n43[1]);
    xor g1756(n1532 ,n122 ,n23[3]);
    nor g1757(n1531 ,n121 ,n122);
    nor g1758(n122 ,n117 ,n120);
    nor g1759(n121 ,n23[2] ,n119);
    nor g1760(n1530 ,n119 ,n118);
    not g1761(n120 ,n119);
    nor g1762(n119 ,n116 ,n1529);
    nor g1763(n118 ,n23[1] ,n23[0]);
    not g1764(n117 ,n23[2]);
    not g1765(n1529 ,n23[0]);
    not g1766(n116 ,n23[1]);
    buf g1767(n446 ,n43[4]);
    buf g1768(n515 ,n461);
    not g1769(n438 ,n417);
    buf g1770(n891 ,n464);
    buf g1771(n532 ,n416);
    buf g1772(n1554 ,n115);
    buf g1773(n1319 ,n894);
endmodule
