module top (n0, n1, n5, n6, n2, n3, n9, n14, n15, n7, n8, n4, n16, n17, n10, n11, n12, n13);
    input n0, n1, n2, n3, n4;
    input [31:0] n5, n6;
    input [3:0] n7;
    input [1:0] n8;
    output [31:0] n9, n10, n11, n12, n13;
    output n14, n15, n16;
    output [7:0] n17;
    wire n0, n1, n2, n3, n4;
    wire [31:0] n5, n6;
    wire [3:0] n7;
    wire [1:0] n8;
    wire [31:0] n9, n10, n11, n12, n13;
    wire n14, n15, n16;
    wire [7:0] n17;
    wire [2:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [7:0] n25;
    wire [15:0] n26;
    wire [1:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [7:0] n30;
    wire [15:0] n31;
    wire [15:0] n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526, n527, n528;
    wire n529, n530, n531, n532, n533, n534, n535, n536;
    wire n537, n538, n539, n540, n541, n542, n543, n544;
    wire n545, n546, n547, n548, n549, n550, n551, n552;
    wire n553, n554, n555, n556, n557, n558, n559, n560;
    wire n561, n562, n563, n564, n565, n566, n567, n568;
    wire n569, n570, n571, n572, n573, n574, n575, n576;
    wire n577, n578, n579, n580, n581, n582, n583, n584;
    wire n585, n586, n587, n588, n589, n590, n591, n592;
    wire n593, n594, n595, n596, n597, n598, n599, n600;
    wire n601, n602, n603, n604, n605, n606, n607, n608;
    wire n609, n610, n611, n612, n613, n614, n615, n616;
    wire n617, n618, n619, n620, n621, n622, n623, n624;
    wire n625, n626, n627, n628, n629, n630, n631, n632;
    wire n633, n634, n635, n636, n637, n638, n639, n640;
    wire n641, n642, n643, n644, n645, n646, n647, n648;
    wire n649, n650, n651, n652, n653, n654, n655, n656;
    wire n657, n658, n659, n660, n661, n662, n663, n664;
    wire n665, n666, n667, n668, n669, n670, n671, n672;
    wire n673, n674, n675, n676, n677, n678, n679, n680;
    wire n681, n682, n683, n684, n685, n686, n687, n688;
    wire n689, n690, n691, n692, n693, n694, n695, n696;
    wire n697, n698, n699, n700, n701, n702, n703, n704;
    wire n705, n706, n707, n708, n709, n710, n711, n712;
    wire n713, n714, n715, n716, n717, n718, n719, n720;
    wire n721, n722, n723, n724, n725, n726, n727, n728;
    wire n729, n730, n731, n732, n733, n734, n735, n736;
    wire n737, n738, n739, n740, n741, n742, n743, n744;
    wire n745, n746, n747, n748, n749, n750, n751, n752;
    wire n753, n754, n755, n756, n757, n758, n759, n760;
    wire n761, n762, n763, n764, n765, n766, n767, n768;
    wire n769, n770, n771, n772, n773, n774, n775, n776;
    wire n777, n778, n779, n780, n781, n782, n783, n784;
    wire n785, n786, n787, n788, n789, n790, n791, n792;
    wire n793, n794, n795, n796, n797, n798, n799, n800;
    wire n801, n802, n803, n804, n805, n806, n807, n808;
    wire n809, n810, n811, n812, n813, n814, n815, n816;
    wire n817, n818, n819, n820, n821, n822, n823, n824;
    wire n825, n826, n827, n828, n829, n830, n831, n832;
    wire n833, n834, n835, n836, n837, n838, n839, n840;
    wire n841, n842, n843, n844, n845, n846, n847, n848;
    wire n849, n850, n851, n852, n853, n854, n855, n856;
    wire n857, n858, n859, n860, n861, n862, n863, n864;
    wire n865, n866, n867, n868, n869, n870, n871, n872;
    wire n873, n874, n875, n876, n877, n878, n879, n880;
    wire n881, n882, n883, n884, n885, n886, n887, n888;
    wire n889, n890, n891, n892, n893, n894, n895, n896;
    wire n897, n898, n899, n900, n901, n902, n903, n904;
    wire n905, n906, n907, n908, n909, n910, n911, n912;
    wire n913, n914, n915, n916, n917, n918, n919, n920;
    wire n921, n922, n923, n924, n925, n926, n927, n928;
    wire n929, n930, n931, n932, n933, n934, n935, n936;
    wire n937, n938, n939, n940, n941, n942, n943, n944;
    wire n945, n946, n947, n948, n949, n950, n951, n952;
    wire n953, n954, n955, n956, n957, n958, n959, n960;
    wire n961, n962, n963, n964, n965, n966, n967, n968;
    wire n969, n970, n971, n972, n973, n974, n975, n976;
    wire n977, n978, n979, n980, n981, n982, n983, n984;
    wire n985, n986, n987, n988, n989, n990, n991, n992;
    wire n993, n994, n995, n996, n997, n998, n999, n1000;
    wire n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
    wire n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
    wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
    wire n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
    wire n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
    wire n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
    wire n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
    wire n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064;
    wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
    wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
    wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
    wire n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096;
    wire n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
    wire n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;
    wire n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120;
    wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
    wire n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136;
    wire n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
    wire n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152;
    wire n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
    wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168;
    wire n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176;
    wire n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184;
    wire n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192;
    wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
    wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
    wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
    wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
    wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
    wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
    wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
    wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
    wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
    wire n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
    wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
    wire n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288;
    wire n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;
    wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;
    wire n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;
    wire n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;
    wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
    wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
    wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;
    wire n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;
    wire n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;
    wire n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368;
    wire n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;
    wire n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384;
    wire n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392;
    wire n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400;
    wire n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408;
    wire n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416;
    wire n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424;
    wire n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432;
    wire n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440;
    wire n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448;
    wire n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456;
    wire n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464;
    wire n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472;
    wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480;
    wire n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488;
    wire n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496;
    wire n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504;
    wire n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512;
    wire n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520;
    wire n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528;
    wire n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536;
    wire n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544;
    wire n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552;
    wire n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560;
    wire n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568;
    wire n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576;
    wire n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584;
    wire n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592;
    wire n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600;
    wire n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608;
    wire n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616;
    wire n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624;
    wire n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632;
    wire n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640;
    wire n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648;
    wire n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656;
    wire n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664;
    wire n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672;
    wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
    wire n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688;
    wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
    wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
    wire n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712;
    wire n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720;
    wire n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728;
    wire n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736;
    wire n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744;
    wire n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752;
    wire n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760;
    wire n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768;
    wire n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776;
    wire n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;
    wire n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792;
    wire n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800;
    wire n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808;
    wire n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816;
    wire n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824;
    wire n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832;
    wire n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840;
    wire n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848;
    wire n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856;
    wire n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864;
    wire n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872;
    wire n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880;
    wire n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888;
    wire n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896;
    wire n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904;
    wire n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912;
    wire n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920;
    wire n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928;
    wire n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936;
    wire n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944;
    wire n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952;
    wire n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960;
    wire n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968;
    wire n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976;
    wire n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984;
    wire n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992;
    wire n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000;
    wire n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008;
    wire n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016;
    wire n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024;
    wire n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032;
    wire n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040;
    wire n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048;
    wire n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056;
    wire n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064;
    wire n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072;
    wire n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080;
    wire n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088;
    wire n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096;
    wire n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104;
    wire n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112;
    wire n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120;
    wire n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128;
    wire n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136;
    wire n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144;
    wire n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152;
    wire n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160;
    wire n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168;
    wire n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176;
    wire n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184;
    wire n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192;
    wire n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200;
    wire n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208;
    wire n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216;
    wire n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224;
    wire n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232;
    wire n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240;
    wire n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248;
    wire n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256;
    wire n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264;
    wire n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272;
    wire n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280;
    wire n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288;
    wire n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296;
    wire n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304;
    wire n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312;
    wire n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320;
    wire n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328;
    wire n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336;
    wire n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344;
    wire n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352;
    wire n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360;
    wire n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368;
    wire n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376;
    wire n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384;
    wire n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392;
    wire n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400;
    wire n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408;
    wire n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416;
    wire n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424;
    wire n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432;
    wire n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440;
    wire n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448;
    wire n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456;
    wire n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464;
    wire n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472;
    wire n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480;
    wire n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488;
    wire n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496;
    wire n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504;
    wire n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512;
    wire n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520;
    wire n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528;
    wire n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536;
    wire n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544;
    wire n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552;
    wire n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560;
    wire n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568;
    wire n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576;
    wire n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584;
    wire n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592;
    wire n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600;
    wire n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608;
    wire n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616;
    wire n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624;
    wire n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632;
    wire n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640;
    wire n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648;
    wire n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656;
    wire n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664;
    wire n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672;
    wire n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680;
    wire n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688;
    wire n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696;
    wire n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704;
    wire n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712;
    wire n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720;
    wire n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728;
    wire n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736;
    wire n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744;
    wire n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752;
    wire n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760;
    wire n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768;
    wire n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776;
    wire n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784;
    wire n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792;
    wire n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800;
    wire n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808;
    wire n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816;
    wire n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824;
    wire n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832;
    wire n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840;
    wire n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848;
    wire n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856;
    wire n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864;
    wire n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872;
    wire n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880;
    wire n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888;
    wire n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896;
    wire n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904;
    wire n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912;
    wire n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920;
    wire n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928;
    wire n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936;
    wire n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944;
    wire n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952;
    wire n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960;
    wire n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968;
    wire n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976;
    wire n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984;
    wire n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992;
    wire n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000;
    wire n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008;
    wire n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016;
    wire n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024;
    wire n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032;
    wire n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040;
    wire n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048;
    wire n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056;
    wire n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064;
    wire n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072;
    wire n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080;
    wire n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088;
    wire n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096;
    wire n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104;
    wire n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112;
    wire n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120;
    wire n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128;
    wire n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136;
    wire n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144;
    wire n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152;
    wire n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160;
    wire n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168;
    wire n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176;
    wire n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184;
    wire n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192;
    wire n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200;
    wire n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208;
    wire n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216;
    wire n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224;
    wire n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232;
    wire n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240;
    wire n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248;
    wire n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256;
    wire n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264;
    wire n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272;
    wire n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280;
    wire n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288;
    wire n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296;
    wire n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304;
    wire n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312;
    wire n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320;
    wire n3321, n3322, n3323;
    nor g0(n1745 ,n1697 ,n1721);
    not g1(n2657 ,n2656);
    nor g2(n791 ,n128 ,n655);
    not g3(n161 ,n10[3]);
    not g4(n1716 ,n1715);
    dff g5(.RN(n1), .SN(1'b1), .CK(n0), .D(n844), .Q(n20[4]));
    dff g6(.RN(n1), .SN(1'b1), .CK(n0), .D(n848), .Q(n20[0]));
    xnor g7(n3315 ,n3024 ,n3051);
    nor g8(n1537 ,n1523 ,n1512);
    nor g9(n674 ,n107 ,n661);
    xnor g10(n1486 ,n1463 ,n1435);
    nor g11(n2952 ,n2951 ,n2915);
    nor g12(n1136 ,n1049 ,n1102);
    xor g13(n3284 ,n2930 ,n2949);
    buf g14(n9[28], 1'b0);
    nor g15(n3176 ,n3087 ,n3141);
    or g16(n3163 ,n3154 ,n3138);
    nor g17(n1116 ,n958 ,n1064);
    nor g18(n456 ,n163 ,n102);
    nor g19(n2172 ,n2025 ,n2077);
    nor g20(n1361 ,n1329 ,n1322);
    nor g21(n2010 ,n1869 ,n1891);
    nor g22(n1095 ,n1012 ,n1069);
    nor g23(n2951 ,n2924 ,n2950);
    nor g24(n2681 ,n2580 ,n2629);
    not g25(n1734 ,n1733);
    nor g26(n727 ,n125 ,n649);
    nor g27(n989 ,n961 ,n971);
    or g28(n605 ,n379 ,n356);
    not g29(n191 ,n20[4]);
    not g30(n1232 ,n942);
    nor g31(n1102 ,n949 ,n1062);
    not g32(n1756 ,n1755);
    nor g33(n1449 ,n1416 ,n1422);
    nor g34(n415 ,n258 ,n349);
    nor g35(n1614 ,n1521 ,n1558);
    nor g36(n1114 ,n960 ,n1064);
    nor g37(n1618 ,n1520 ,n1551);
    nor g38(n520 ,n168 ,n348);
    nor g39(n3183 ,n3095 ,n3141);
    not g40(n1874 ,n22[2]);
    xor g41(n931 ,n30[7] ,n77);
    dff g42(.RN(n1), .SN(1'b1), .CK(n0), .D(n581), .Q(n25[5]));
    not g43(n154 ,n9[1]);
    buf g44(n9[21], 1'b0);
    xnor g45(n1788 ,n1747 ,n1700);
    xnor g46(n1293 ,n1213 ,n1212);
    nor g47(n2095 ,n1882 ,n1891);
    buf g48(n360 ,n347);
    nor g49(n937 ,n62 ,n61);
    or g50(n556 ,n396 ,n484);
    xnor g51(n1217 ,n1159 ,n1028);
    xor g52(n924 ,n25[7] ,n101);
    xnor g53(n2477 ,n2181 ,n2379);
    xnor g54(n3037 ,n3301 ,n3285);
    or g55(n535 ,n376 ,n453);
    xnor g56(n3028 ,n3290 ,n3274);
    nor g57(n2153 ,n1905 ,n1929);
    not g58(n75 ,n74);
    nor g59(n2510 ,n2368 ,n2396);
    buf g60(n12[23], n10[15]);
    xnor g61(n2654 ,n2536 ,n2459);
    nor g62(n2025 ,n1869 ,n1878);
    buf g63(n13[29], n10[5]);
    nor g64(n426 ,n282 ,n347);
    dff g65(.RN(n1), .SN(1'b1), .CK(n0), .D(n847), .Q(n20[1]));
    nor g66(n698 ,n111 ,n659);
    not g67(n3126 ,n3285);
    xnor g68(n1735 ,n1673 ,n1669);
    xnor g69(n1552 ,n3266 ,n23[2]);
    nor g70(n2628 ,n2524 ,n2567);
    not g71(n66 ,n65);
    buf g72(n12[7], 1'b0);
    nor g73(n480 ,n173 ,n104);
    not g74(n998 ,n997);
    not g75(n1718 ,n1717);
    buf g76(n11[19], n10[3]);
    dff g77(.RN(n1), .SN(1'b1), .CK(n0), .D(n571), .Q(n26[5]));
    nor g78(n1698 ,n1586 ,n1649);
    nor g79(n1495 ,n1454 ,n1494);
    nor g80(n70 ,n30[4] ,n68);
    not g81(n3058 ,n3057);
    or g82(n1064 ,n1021 ,n1035);
    xnor g83(n2690 ,n2612 ,n2634);
    not g84(n2134 ,n2133);
    not g85(n3115 ,n3298);
    or g86(n557 ,n438 ,n513);
    dff g87(.RN(n1), .SN(1'b1), .CK(n0), .D(n565), .Q(n26[9]));
    buf g88(n10[19], 1'b0);
    or g89(n641 ,n5[4] ,n639);
    xnor g90(n2394 ,n2260 ,n1997);
    nor g91(n1391 ,n1353 ,n1351);
    xor g92(n3270 ,n20[6] ,n21[6]);
    not g93(n648 ,n649);
    nor g94(n2323 ,n2281 ,n2278);
    or g95(n46 ,n30[7] ,n45);
    not g96(n1511 ,n23[5]);
    not g97(n2013 ,n2012);
    nor g98(n614 ,n231 ,n524);
    xnor g99(n1719 ,n1642 ,n1628);
    not g100(n1777 ,n1776);
    not g101(n1025 ,n1026);
    xnor g102(n2585 ,n2416 ,n2502);
    not g103(n1916 ,n1915);
    or g104(n846 ,n740 ,n697);
    nor g105(n501 ,n135 ,n346);
    xnor g106(n1419 ,n1379 ,n1356);
    not g107(n286 ,n30[2]);
    nor g108(n1452 ,n1413 ,n1424);
    not g109(n2421 ,n2420);
    nor g110(n1007 ,n976 ,n988);
    not g111(n1341 ,n1340);
    nor g112(n1466 ,n1441 ,n1447);
    xnor g113(n2410 ,n2259 ,n2010);
    nor g114(n1342 ,n1277 ,n1311);
    nor g115(n797 ,n217 ,n655);
    nor g116(n2941 ,n2914 ,n2931);
    or g117(n569 ,n405 ,n476);
    nor g118(n1369 ,n1255 ,n1323);
    not g119(n152 ,n31[10]);
    xnor g120(n1228 ,n1028 ,n1145);
    xor g121(n3286 ,n2882 ,n2953);
    nor g122(n813 ,n192 ,n665);
    not g123(n1811 ,n1810);
    not g124(n227 ,n10[15]);
    nor g125(n507 ,n149 ,n346);
    xnor g126(n1173 ,n1017 ,n1098);
    nor g127(n2565 ,n2467 ,n2492);
    not g128(n3084 ,n3286);
    xnor g129(n328 ,n208 ,n186);
    nor g130(n2811 ,n2733 ,n2765);
    not g131(n2919 ,n2918);
    xnor g132(n2249 ,n2055 ,n2079);
    nor g133(n611 ,n320 ,n351);
    not g134(n1912 ,n1911);
    not g135(n2417 ,n2416);
    nor g136(n1682 ,n1663 ,n1630);
    nor g137(n1810 ,n1783 ,n1800);
    not g138(n69 ,n68);
    or g139(n895 ,n886 ,n884);
    nor g140(n1683 ,n1627 ,n1648);
    or g141(n43 ,n30[1] ,n41);
    xnor g142(n1295 ,n1203 ,n1220);
    nor g143(n3186 ,n3079 ,n3141);
    nor g144(n464 ,n142 ,n104);
    nor g145(n812 ,n122 ,n654);
    xnor g146(n1795 ,n1729 ,n1759);
    nor g147(n719 ,n195 ,n651);
    nor g148(n1919 ,n1885 ,n1889);
    nor g149(n370 ,n237 ,n103);
    dff g150(.RN(n1), .SN(1'b1), .CK(n0), .D(n528), .Q(n29[9]));
    nor g151(n1406 ,n1370 ,n1376);
    not g152(n174 ,n927);
    or g153(n1536 ,n1516 ,n1518);
    or g154(n599 ,n428 ,n508);
    nor g155(n3063 ,n3037 ,n3062);
    nor g156(n1610 ,n1521 ,n1552);
    or g157(n870 ,n800 ,n799);
    nor g158(n1258 ,n1212 ,n1213);
    or g159(n299 ,n5[27] ,n5[26]);
    nor g160(n1050 ,n948 ,n1034);
    nor g161(n2325 ,n2190 ,n2317);
    nor g162(n720 ,n207 ,n651);
    nor g163(n759 ,n220 ,n658);
    nor g164(n1408 ,n943 ,n1382);
    nor g165(n1817 ,n1771 ,n1798);
    not g166(n2054 ,n2053);
    or g167(n842 ,n736 ,n693);
    nor g168(n1262 ,n1172 ,n1239);
    or g169(n886 ,n812 ,n811);
    nor g170(n3008 ,n3291 ,n3275);
    or g171(n652 ,n523 ,n647);
    nor g172(n476 ,n147 ,n102);
    not g173(n1525 ,n23[1]);
    dff g174(.RN(n1), .SN(1'b1), .CK(n0), .D(n540), .Q(n29[2]));
    xnor g175(n2918 ,n2883 ,n2870);
    buf g176(n17[5], 1'b0);
    dff g177(.RN(n1), .SN(1'b1), .CK(n0), .D(n917), .Q(n9[3]));
    nor g178(n2784 ,n2712 ,n2748);
    xnor g179(n1789 ,n1749 ,n1735);
    nor g180(n2897 ,n2775 ,n2872);
    nor g181(n1971 ,n1865 ,n1861);
    xnor g182(n2543 ,n2410 ,n2400);
    nor g183(n2367 ,n2204 ,n2290);
    buf g184(n11[7], 1'b0);
    nor g185(n2327 ,n2195 ,n2299);
    nor g186(n2866 ,n2792 ,n2851);
    nor g187(n2352 ,n2196 ,n2292);
    xnor g188(n2252 ,n2075 ,n1943);
    dff g189(.RN(n1), .SN(1'b1), .CK(n0), .D(n623), .Q(n26[1]));
    not g190(n1479 ,n1478);
    xnor g191(n1251 ,n1178 ,n1090);
    not g192(n3116 ,n3293);
    nor g193(n1164 ,n1050 ,n1119);
    not g194(n103 ,n104);
    nor g195(n455 ,n133 ,n102);
    xnor g196(n2398 ,n2258 ,n2104);
    nor g197(n621 ,n154 ,n524);
    dff g198(.RN(n1), .SN(1'b1), .CK(n0), .D(n534), .Q(n28[15]));
    not g199(n319 ,n318);
    nor g200(n1797 ,n1778 ,n1772);
    nor g201(n2573 ,n2432 ,n2485);
    nor g202(n1925 ,n1867 ,n1881);
    not g203(n2270 ,n2269);
    dff g204(.RN(n1), .SN(1'b1), .CK(n0), .D(n560), .Q(n26[14]));
    nor g205(n2778 ,n2707 ,n2741);
    xnor g206(n1457 ,n1423 ,n1413);
    or g207(n1063 ,n1024 ,n1033);
    nor g208(n357 ,n104 ,n334);
    not g209(n223 ,n17[4]);
    dff g210(.RN(n1), .SN(1'b1), .CK(n0), .D(n883), .Q(n23[7]));
    xnor g211(n2981 ,n22[3] ,n23[3]);
    nor g212(n1273 ,n1221 ,n1216);
    not g213(n2956 ,n23[2]);
    dff g214(.RN(n1), .SN(1'b1), .CK(n0), .D(n569), .Q(n26[6]));
    xor g215(n3262 ,n3036 ,n3064);
    not g216(n1422 ,n1421);
    nor g217(n2187 ,n1968 ,n1970);
    nor g218(n424 ,n235 ,n347);
    dff g219(.RN(n1), .SN(1'b1), .CK(n0), .D(n832), .Q(n21[6]));
    xnor g220(n2638 ,n2408 ,n2557);
    nor g221(n3044 ,n3026 ,n3043);
    not g222(n2887 ,n2886);
    nor g223(n1741 ,n1656 ,n1713);
    nor g224(n1277 ,n1223 ,n1217);
    not g225(n287 ,n10[14]);
    not g226(n1714 ,n1713);
    nor g227(n3199 ,n3125 ,n3142);
    nor g228(n1911 ,n1885 ,n1888);
    not g229(n2464 ,n2463);
    not g230(n1586 ,n1585);
    xnor g231(n1360 ,n1295 ,n1245);
    nor g232(n1383 ,n1191 ,n1362);
    nor g233(n1539 ,n1519 ,n1538);
    nor g234(n1565 ,n1519 ,n1533);
    nor g235(n1125 ,n956 ,n1089);
    nor g236(n2118 ,n1879 ,n1878);
    not g237(n1862 ,n23[7]);
    xnor g238(n527 ,n348 ,n25[0]);
    nor g239(n2437 ,n2180 ,n2349);
    nor g240(n770 ,n206 ,n655);
    nor g241(n2021 ,n1864 ,n1877);
    nor g242(n3188 ,n3086 ,n3142);
    nor g243(n1078 ,n958 ,n1040);
    not g244(n117 ,n27[0]);
    xnor g245(n2234 ,n1957 ,n1971);
    nor g246(n1190 ,n1017 ,n1171);
    xnor g247(n1225 ,n1030 ,n1138);
    buf g248(n12[12], n10[4]);
    not g249(n965 ,n20[4]);
    dff g250(.RN(n1), .SN(1'b1), .CK(n0), .D(n562), .Q(n26[11]));
    nor g251(n431 ,n277 ,n347);
    buf g252(n12[21], n10[13]);
    not g253(n1180 ,n1179);
    xnor g254(n1017 ,n997 ,n978);
    or g255(n606 ,n397 ,n488);
    not g256(n2072 ,n2071);
    dff g257(.RN(n1), .SN(1'b1), .CK(n0), .D(n588), .Q(n10[14]));
    nor g258(n1139 ,n1051 ,n1105);
    nor g259(n2310 ,n2002 ,n2165);
    nor g260(n817 ,n189 ,n656);
    or g261(n363 ,n26[12] ,n343);
    buf g262(n11[1], 1'b0);
    not g263(n167 ,n929);
    not g264(n2552 ,n2551);
    xnor g265(n1244 ,n1028 ,n1152);
    nor g266(n795 ,n130 ,n665);
    not g267(n2998 ,n3301);
    or g268(n337 ,n18[0] ,n319);
    nor g269(n3131 ,n3316 ,n32[9]);
    nor g270(n3180 ,n3113 ,n3142);
    nor g271(n2033 ,n1885 ,n1870);
    nor g272(n3045 ,n3013 ,n3044);
    nor g273(n1386 ,n1366 ,n1360);
    not g274(n283 ,n9[2]);
    nor g275(n3209 ,n3094 ,n3155);
    nor g276(n2443 ,n2378 ,n2360);
    xnor g277(n1733 ,n1675 ,n1648);
    nor g278(n784 ,n181 ,n652);
    not g279(n2272 ,n2271);
    nor g280(n1937 ,n1892 ,n1888);
    nor g281(n1130 ,n959 ,n1064);
    nor g282(n1168 ,n1080 ,n1123);
    or g283(n844 ,n738 ,n695);
    nor g284(n2439 ,n2328 ,n2326);
    nor g285(n450 ,n135 ,n104);
    not g286(n2659 ,n2658);
    not g287(n2431 ,n2430);
    nor g288(n1991 ,n1863 ,n1878);
    not g289(n271 ,n29[3]);
    not g290(n2589 ,n2588);
    nor g291(n2204 ,n2066 ,n1912);
    xnor g292(n1399 ,n1358 ,n1280);
    nor g293(n755 ,n150 ,n658);
    not g294(n1602 ,n1601);
    nor g295(n1642 ,n1548 ,n1589);
    nor g296(n800 ,n214 ,n654);
    nor g297(n1105 ,n946 ,n1062);
    xor g298(n3267 ,n20[3] ,n21[3]);
    nor g299(n3212 ,n3073 ,n3155);
    nor g300(n2636 ,n2509 ,n2566);
    nor g301(n474 ,n232 ,n102);
    xnor g302(n2385 ,n2273 ,n2226);
    not g303(n278 ,n29[13]);
    not g304(n2078 ,n2077);
    nor g305(n392 ,n204 ,n105);
    nor g306(n684 ,n113 ,n650);
    not g307(n1265 ,n1264);
    not g308(n141 ,n10[4]);
    nor g309(n2139 ,n1882 ,n1866);
    not g310(n1645 ,n1644);
    nor g311(n375 ,n261 ,n105);
    xnor g312(n1321 ,n1167 ,n1285);
    nor g313(n373 ,n291 ,n105);
    nor g314(n2881 ,n2782 ,n2844);
    nor g315(n1981 ,n1871 ,n1876);
    xnor g316(n2278 ,n2108 ,n1981);
    or g317(n2103 ,n1884 ,n1891);
    not g318(n1428 ,n1427);
    xor g319(n2470 ,n2264 ,n2115);
    nor g320(n1081 ,n959 ,n1038);
    not g321(n193 ,n23[7]);
    xnor g322(n326 ,n210 ,n188);
    nor g323(n2893 ,n2880 ,n2871);
    nor g324(n379 ,n271 ,n105);
    nor g325(n2820 ,n2747 ,n2779);
    nor g326(n2156 ,n1967 ,n1969);
    not g327(n139 ,n10[10]);
    or g328(n851 ,n747 ,n700);
    not g329(n2425 ,n2424);
    buf g330(n11[9], 1'b0);
    nor g331(n3150 ,n3106 ,n3101);
    nor g332(n2511 ,n2333 ,n2393);
    buf g333(n11[29], n10[13]);
    not g334(n183 ,n18[1]);
    nor g335(n1333 ,n1265 ,n1319);
    xnor g336(n1035 ,n938 ,n1008);
    xnor g337(n1806 ,n1770 ,n1757);
    nor g338(n664 ,n323 ,n646);
    nor g339(n3203 ,n3090 ,n3141);
    dff g340(.RN(n1), .SN(1'b1), .CK(n0), .D(n548), .Q(n28[8]));
    nor g341(n741 ,n194 ,n662);
    nor g342(n1084 ,n959 ,n1032);
    xnor g343(n980 ,n961 ,n21[3]);
    nor g344(n1115 ,n960 ,n1062);
    not g345(n3002 ,n3283);
    buf g346(n9[24], 1'b0);
    nor g347(n740 ,n192 ,n662);
    nor g348(n2163 ,n1907 ,n2063);
    buf g349(n11[26], n10[10]);
    or g350(n531 ,n443 ,n494);
    nor g351(n1011 ,n985 ,n981);
    nor g352(n1853 ,n1838 ,n1852);
    not g353(n2395 ,n2394);
    nor g354(n1121 ,n957 ,n1089);
    or g355(n312 ,n5[15] ,n5[14]);
    nor g356(n383 ,n233 ,n103);
    nor g357(n2154 ,n2067 ,n1933);
    nor g358(n1381 ,n1333 ,n1363);
    buf g359(n13[31], n10[7]);
    nor g360(n2718 ,n2604 ,n2655);
    not g361(n1036 ,n1035);
    nor g362(n1096 ,n1001 ,n1088);
    nor g363(n1401 ,n1330 ,n1387);
    nor g364(n2213 ,n1924 ,n2058);
    not g365(n1914 ,n1913);
    xnor g366(n1150 ,n1025 ,n1041);
    nor g367(n1773 ,n1723 ,n1759);
    nor g368(n514 ,n178 ,n348);
    nor g369(n3304 ,n2971 ,n2969);
    buf g370(n12[27], 1'b0);
    dff g371(.RN(n1), .SN(1'b1), .CK(n0), .D(n543), .Q(n28[14]));
    nor g372(n681 ,n114 ,n650);
    not g373(n1349 ,n1348);
    nor g374(n1763 ,n1732 ,n1734);
    xor g375(n3283 ,n2940 ,n2947);
    not g376(n1656 ,n1655);
    nor g377(n669 ,n106 ,n650);
    nor g378(n85 ,n25[1] ,n25[0]);
    not g379(n946 ,n3305);
    not g380(n290 ,n28[11]);
    xnor g381(n2978 ,n22[4] ,n23[4]);
    nor g382(n2555 ,n2434 ,n2490);
    or g383(n315 ,n7[3] ,n7[2]);
    nor g384(n1652 ,n1578 ,n1622);
    not g385(n1906 ,n1905);
    buf g386(n10[27], 1'b0);
    nor g387(n1670 ,n1564 ,n1611);
    nor g388(n1842 ,n1817 ,n1828);
    not g389(n957 ,n3309);
    nor g390(n728 ,n213 ,n649);
    or g391(n992 ,n978 ,n972);
    nor g392(n2983 ,n2966 ,n2982);
    nor g393(n2869 ,n2836 ,n2849);
    not g394(n2020 ,n2019);
    or g395(n314 ,n5[8] ,n5[7]);
    nor g396(n2320 ,n2042 ,n2221);
    xnor g397(n2687 ,n2615 ,n2555);
    nor g398(n1119 ,n957 ,n1063);
    buf g399(n9[18], 1'b0);
    nor g400(n2486 ,n2404 ,n2420);
    buf g401(n10[20], 1'b0);
    nor g402(n2666 ,n2556 ,n2591);
    nor g403(n1547 ,n1522 ,n1530);
    xnor g404(n1299 ,n1227 ,n1194);
    nor g405(n2498 ,n2356 ,n2441);
    nor g406(n1613 ,n1522 ,n1553);
    nor g407(n712 ,n112 ,n663);
    not g408(n122 ,n23[2]);
    not g409(n1960 ,n1959);
    dff g410(.RN(n1), .SN(1'b1), .CK(n0), .D(n582), .Q(n28[3]));
    not g411(n996 ,n995);
    nor g412(n785 ,n207 ,n655);
    xnor g413(n2243 ,n2087 ,n2081);
    not g414(n1436 ,n1435);
    not g415(n220 ,n24[1]);
    nor g416(n1507 ,n1506 ,n1467);
    nor g417(n2148 ,n1895 ,n2027);
    nor g418(n77 ,n54 ,n75);
    nor g419(n404 ,n202 ,n103);
    nor g420(n692 ,n111 ,n661);
    nor g421(n1256 ,n1220 ,n1203);
    nor g422(n1006 ,n977 ,n989);
    nor g423(n2876 ,n2818 ,n2845);
    not g424(n2795 ,n2794);
    dff g425(.RN(n1), .SN(1'b1), .CK(n0), .D(n611), .Q(n18[0]));
    nor g426(n1077 ,n960 ,n1034);
    not g427(n2846 ,n2845);
    xnor g428(n1211 ,n1029 ,n1154);
    nor g429(n2578 ,n2470 ,n2491);
    not g430(n113 ,n6[3]);
    not g431(n230 ,n28[9]);
    or g432(n923 ,n36 ,n39);
    buf g433(n12[24], 1'b0);
    not g434(n1869 ,n21[1]);
    nor g435(n2508 ,n2464 ,n2452);
    nor g436(n1051 ,n949 ,n1038);
    nor g437(n1364 ,n1335 ,n1344);
    xnor g438(n1456 ,n1422 ,n1415);
    not g439(n2853 ,n2852);
    nor g440(n2831 ,n2780 ,n2805);
    not g441(n964 ,n20[3]);
    nor g442(n2081 ,n1886 ,n1872);
    not g443(n1066 ,n1065);
    not g444(n255 ,n28[15]);
    nor g445(n708 ,n113 ,n657);
    not g446(n2965 ,n23[4]);
    buf g447(n17[0], n17[2]);
    nor g448(n715 ,n109 ,n663);
    not g449(n143 ,n31[9]);
    dff g450(.RN(n1), .SN(1'b1), .CK(n0), .D(n557), .Q(n17[4]));
    dff g451(.RN(n1), .SN(1'b1), .CK(n0), .D(n633), .Q(n18[1]));
    nor g452(n2577 ,n2431 ,n2486);
    or g453(n344 ,n18[2] ,n321);
    not g454(n2125 ,n2124);
    xnor g455(n2892 ,n2843 ,n2781);
    nor g456(n1387 ,n1326 ,n1348);
    xnor g457(n2269 ,n2130 ,n2124);
    buf g458(n11[11], 1'b0);
    not g459(n2921 ,n2920);
    nor g460(n44 ,n42 ,n43);
    or g461(n302 ,n26[13] ,n26[14]);
    buf g462(n13[10], 1'b0);
    nor g463(n1237 ,n1184 ,n1197);
    or g464(n1532 ,n1514 ,n1515);
    nor g465(n1189 ,n1028 ,n1147);
    buf g466(n10[17], 1'b0);
    or g467(n295 ,n26[4] ,n26[5]);
    or g468(n647 ,n323 ,n642);
    nor g469(n421 ,n254 ,n347);
    not g470(n125 ,n21[7]);
    xnor g471(n2723 ,n2646 ,n2498);
    not g472(n107 ,n6[0]);
    nor g473(n98 ,n83 ,n96);
    xnor g474(n2700 ,n2587 ,n2594);
    xnor g475(n2232 ,n2039 ,n1927);
    nor g476(n1316 ,n1269 ,n1282);
    nor g477(n1669 ,n1541 ,n1607);
    or g478(n868 ,n618 ,n795);
    nor g479(n1429 ,n1392 ,n1406);
    not g480(n1883 ,n20[0]);
    xnor g481(n1459 ,n1418 ,n1381);
    not g482(n2121 ,n2120);
    not g483(n1266 ,n945);
    or g484(n343 ,n303 ,n296);
    nor g485(n73 ,n30[5] ,n71);
    nor g486(n320 ,n184 ,n18[1]);
    xor g487(n2254 ,n2003 ,n2073);
    not g488(n106 ,n6[1]);
    not g489(n1968 ,n1967);
    nor g490(n2445 ,n2182 ,n2329);
    nor g491(n732 ,n127 ,n649);
    not g492(n216 ,n23[3]);
    xnor g493(n2457 ,n2262 ,n2071);
    not g494(n1176 ,n1175);
    not g495(n2136 ,n2135);
    xor g496(n943 ,n1183 ,n1241);
    xnor g497(n2382 ,n2275 ,n2228);
    or g498(n847 ,n741 ,n673);
    nor g499(n2359 ,n2227 ,n2273);
    nor g500(n709 ,n109 ,n657);
    not g501(n63 ,n62);
    nor g502(n2500 ,n2359 ,n2435);
    nor g503(n1739 ,n1680 ,n1722);
    nor g504(n330 ,n3 ,n293);
    nor g505(n391 ,n210 ,n105);
    nor g506(n2191 ,n2018 ,n2060);
    xnor g507(n2734 ,n2641 ,n2630);
    xnor g508(n2414 ,n2234 ,n2101);
    xnor g509(n1292 ,n1202 ,n1149);
    not g510(n121 ,n28[1]);
    nor g511(n3047 ,n3019 ,n3046);
    nor g512(n1308 ,n1166 ,n1263);
    nor g513(n805 ,n216 ,n654);
    not g514(n2797 ,n2796);
    dff g515(.RN(n1), .SN(1'b1), .CK(n0), .D(n603), .Q(n10[0]));
    nor g516(n2363 ,n1953 ,n2272);
    nor g517(n2990 ,n2972 ,n2989);
    nor g518(n2750 ,n2661 ,n2717);
    dff g519(.RN(n1), .SN(1'b1), .CK(n0), .D(n350), .Q(n17[2]));
    nor g520(n3148 ,n3109 ,n3071);
    nor g521(n2712 ,n2498 ,n2647);
    nor g522(n68 ,n57 ,n66);
    nor g523(n753 ,n256 ,n658);
    xnor g524(n3313 ,n3031 ,n3055);
    nor g525(n1100 ,n958 ,n1062);
    nor g526(n649 ,n324 ,n646);
    not g527(n1958 ,n1957);
    nor g528(n2166 ,n2037 ,n1939);
    nor g529(n2755 ,n2676 ,n2709);
    nor g530(n1832 ,n1804 ,n1806);
    xnor g531(n995 ,n20[3] ,n21[3]);
    nor g532(n1310 ,n1244 ,n1268);
    xnor g533(n1026 ,n1005 ,n984);
    not g534(n1319 ,n1318);
    xnor g535(n2586 ,n2426 ,n2496);
    buf g536(n12[25], 1'b0);
    xnor g537(n2473 ,n2333 ,n2374);
    not g538(n3127 ,n3273);
    nor g539(n2669 ,n2552 ,n2592);
    buf g540(n13[15], 1'b0);
    nor g541(n1740 ,n1696 ,n1727);
    not g542(n1091 ,n1090);
    xnor g543(n2594 ,n2482 ,n2406);
    xnor g544(n2765 ,n2687 ,n2590);
    dff g545(.RN(n1), .SN(1'b1), .CK(n0), .D(n826), .Q(n22[2]));
    nor g546(n1569 ,n1521 ,n1531);
    nor g547(n2037 ,n1880 ,n1872);
    nor g548(n64 ,n30[2] ,n62);
    xnor g549(n1347 ,n1250 ,n1305);
    not g550(n239 ,n10[0]);
    nor g551(n394 ,n208 ,n105);
    nor g552(n2948 ,n2947 ,n2937);
    nor g553(n651 ,n325 ,n646);
    dff g554(.RN(n1), .SN(1'b1), .CK(n0), .D(n555), .Q(n28[0]));
    nor g555(n478 ,n279 ,n102);
    nor g556(n1953 ,n1883 ,n1874);
    or g557(n830 ,n726 ,n670);
    or g558(n297 ,n5[5] ,n5[0]);
    buf g559(n11[23], n10[7]);
    not g560(n3122 ,n3278);
    not g561(n1884 ,n21[3]);
    not g562(n135 ,n31[11]);
    nor g563(n737 ,n130 ,n662);
    xnor g564(n2886 ,n2838 ,n2859);
    nor g565(n3061 ,n3035 ,n3060);
    not g566(n2772 ,n2771);
    nor g567(n686 ,n111 ,n648);
    buf g568(n13[7], 1'b0);
    nor g569(n3170 ,n3115 ,n3141);
    nor g570(n2099 ,n1869 ,n1888);
    nor g571(n1860 ,n1801 ,n1859);
    xnor g572(n3316 ,n3025 ,n3049);
    xnor g573(n1023 ,n1009 ,n984);
    nor g574(n694 ,n112 ,n661);
    not g575(n1633 ,n1632);
    xnor g576(n1823 ,n1791 ,n1768);
    nor g577(n2697 ,n2583 ,n2680);
    xnor g578(n2422 ,n2244 ,n2001);
    buf g579(n11[22], n10[6]);
    not g580(n2391 ,n2390);
    nor g581(n2533 ,n2357 ,n2443);
    nor g582(n929 ,n88 ,n89);
    xnor g583(n2247 ,n1933 ,n2067);
    nor g584(n2581 ,n2446 ,n2488);
    not g585(n2462 ,n2461);
    nor g586(n2760 ,n2664 ,n2697);
    nor g587(n1679 ,n1640 ,n1638);
    or g588(n3224 ,n3181 ,n3213);
    nor g589(n1058 ,n949 ,n1034);
    or g590(n528 ,n367 ,n449);
    nor g591(n1676 ,n1605 ,n1672);
    nor g592(n2548 ,n2469 ,n2487);
    not g593(n243 ,n9[3]);
    xnor g594(n3288 ,n1017 ,n1039);
    or g595(n903 ,n837 ,n834);
    or g596(n1089 ,n953 ,n1031);
    not g597(n259 ,n10[1]);
    nor g598(n1545 ,n1522 ,n1538);
    nor g599(n2906 ,n2862 ,n2896);
    nor g600(n2143 ,n2091 ,n1909);
    not g601(n956 ,n3307);
    xnor g602(n2740 ,n2639 ,n2592);
    not g603(n2048 ,n2047);
    or g604(n628 ,n473 ,n563);
    xnor g605(n1686 ,n1559 ,n1603);
    not g606(n211 ,n22[3]);
    nor g607(n3168 ,n3080 ,n3141);
    or g608(n890 ,n765 ,n714);
    nor g609(n484 ,n270 ,n102);
    nor g610(n2220 ,n2107 ,n2013);
    nor g611(n2972 ,n2957 ,n2965);
    nor g612(n2518 ,n2337 ,n2413);
    not g613(n2060 ,n2059);
    nor g614(n771 ,n215 ,n666);
    xnor g615(n1487 ,n1462 ,n1445);
    dff g616(.RN(n1), .SN(1'b1), .CK(n0), .D(n640), .Q(n16));
    xnor g617(n1301 ,n1240 ,n1148);
    xnor g618(n1375 ,n1342 ,n945);
    xor g619(n3260 ,n3035 ,n3060);
    or g620(n31[4] ,n3245 ,n3255);
    or g621(n852 ,n745 ,n717);
    nor g622(n1101 ,n948 ,n1062);
    nor g623(n2378 ,n2202 ,n2314);
    dff g624(.RN(n1), .SN(1'b1), .CK(n0), .D(n607), .Q(n29[5]));
    nor g625(n1126 ,n948 ,n1089);
    not g626(n1208 ,n1207);
    nor g627(n1097 ,n1004 ,n1075);
    nor g628(n1160 ,n1087 ,n1130);
    not g629(n1359 ,n1358);
    nor g630(n2783 ,n2718 ,n2750);
    xor g631(n2261 ,n2132 ,n2057);
    nor g632(n2932 ,n2908 ,n2922);
    nor g633(n2634 ,n2518 ,n2564);
    not g634(n2582 ,n2581);
    not g635(n1750 ,n1749);
    dff g636(.RN(n1), .SN(1'b1), .CK(n0), .D(n593), .Q(n10[10]));
    not g637(n1448 ,n1447);
    not g638(n3123 ,n3282);
    nor g639(n2953 ,n2901 ,n2952);
    buf g640(n9[29], 1'b0);
    nor g641(n1591 ,n1521 ,n1556);
    or g642(n31[2] ,n3228 ,n3251);
    not g643(n2591 ,n2590);
    xor g644(n3264 ,n20[0] ,n21[0]);
    not g645(n2219 ,n2218);
    nor g646(n1253 ,n1230 ,n1225);
    xnor g647(n2265 ,n1911 ,n2065);
    nor g648(n2680 ,n2495 ,n2631);
    dff g649(.RN(n1), .SN(1'b1), .CK(n0), .D(n890), .Q(n23[3]));
    nor g650(n3238 ,n3147 ,n3158);
    dff g651(.RN(n1), .SN(1'b1), .CK(n0), .D(n887), .Q(n23[5]));
    nor g652(n2879 ,n2801 ,n2855);
    nor g653(n1057 ,n947 ,n1038);
    or g654(n325 ,n118 ,n5[2]);
    dff g655(.RN(n1), .SN(1'b1), .CK(n0), .D(n820), .Q(n22[6]));
    nor g656(n707 ,n110 ,n657);
    dff g657(.RN(n1), .SN(1'b1), .CK(n0), .D(n573), .Q(n26[3]));
    dff g658(.RN(n1), .SN(1'b1), .CK(n0), .D(n547), .Q(n28[9]));
    not g659(n2752 ,n2751);
    xnor g660(n2250 ,n1925 ,n1917);
    nor g661(n658 ,n525 ,n644);
    not g662(n1872 ,n22[6]);
    not g663(n1966 ,n1965);
    xnor g664(n3275 ,n2723 ,n2722);
    not g665(n2100 ,n2099);
    nor g666(n971 ,n20[4] ,n20[3]);
    or g667(n306 ,n26[0] ,n26[1]);
    not g668(n1894 ,n1893);
    nor g669(n2748 ,n2722 ,n2719);
    not g670(n2058 ,n2057);
    not g671(n1538 ,n1537);
    not g672(n1471 ,n1470);
    xnor g673(n3305 ,n2977 ,n2971);
    nor g674(n2806 ,n2618 ,n2762);
    not g675(n1247 ,n1246);
    nor g676(n678 ,n107 ,n657);
    not g677(n58 ,n30[1]);
    nor g678(n2295 ,n2119 ,n2153);
    not g679(n2593 ,n2592);
    nor g680(n2381 ,n2201 ,n2313);
    nor g681(n749 ,n182 ,n660);
    not g682(n1578 ,n1577);
    dff g683(.RN(n1), .SN(1'b1), .CK(n0), .D(n584), .Q(n25[3]));
    nor g684(n2856 ,n2808 ,n2829);
    buf g685(n17[1], 1'b0);
    not g686(n3003 ,n3299);
    or g687(n530 ,n398 ,n493);
    buf g688(n13[27], n10[3]);
    xnor g689(n2233 ,n1963 ,n1955);
    buf g690(n13[6], 1'b0);
    nor g691(n1048 ,n949 ,n1036);
    dff g692(.RN(n1), .SN(1'b1), .CK(n0), .D(n527), .Q(n25[0]));
    not g693(n1166 ,n1167);
    xnor g694(n3281 ,n2938 ,n2943);
    nor g695(n3214 ,n3100 ,n3155);
    not g696(n3093 ,n3290);
    nor g697(n1080 ,n946 ,n1032);
    dff g698(.RN(n1), .SN(1'b1), .CK(n0), .D(n891), .Q(n23[2]));
    xnor g699(n2917 ,n2888 ,n2852);
    nor g700(n1087 ,n960 ,n1036);
    nor g701(n1437 ,n1393 ,n1407);
    not g702(n1169 ,n1168);
    nor g703(n2208 ,n1962 ,n2052);
    not g704(n136 ,n28[12]);
    dff g705(.RN(n1), .SN(1'b1), .CK(n0), .D(n566), .Q(n26[8]));
    nor g706(n1049 ,n956 ,n1038);
    nor g707(n1540 ,n1522 ,n1533);
    not g708(n321 ,n320);
    not g709(n2332 ,n2331);
    nor g710(n2814 ,n2752 ,n2768);
    nor g711(n3258 ,n1702 ,n1676);
    nor g712(n2186 ,n2044 ,n2062);
    not g713(n2119 ,n2118);
    nor g714(n2942 ,n2927 ,n2941);
    nor g715(n1772 ,n1700 ,n1747);
    not g716(n234 ,n30[6]);
    nor g717(n2108 ,n1864 ,n1875);
    xnor g718(n32[10] ,n1837 ,n1857);
    nor g719(n3143 ,n3104 ,n3069);
    nor g720(n2469 ,n2193 ,n2324);
    nor g721(n2348 ,n2185 ,n2302);
    nor g722(n3133 ,n3322 ,n32[3]);
    xnor g723(n1709 ,n1632 ,n1657);
    or g724(n3228 ,n3212 ,n3189);
    nor g725(n2296 ,n2113 ,n2170);
    or g726(n31[7] ,n3225 ,n3253);
    not g727(n920 ,n922);
    or g728(n646 ,n525 ,n641);
    xnor g729(n2259 ,n2033 ,n2053);
    nor g730(n1499 ,n1498 ,n1483);
    not g731(n245 ,n25[4]);
    nor g732(n700 ,n112 ,n659);
    not g733(n2791 ,n2790);
    nor g734(n1061 ,n948 ,n1038);
    nor g735(n2535 ,n2214 ,n2436);
    nor g736(n2710 ,n2633 ,n2674);
    not g737(n3074 ,n32[8]);
    xnor g738(n2637 ,n2388 ,n2549);
    not g739(n1654 ,n1653);
    nor g740(n1771 ,n1735 ,n1749);
    nor g741(n519 ,n167 ,n348);
    or g742(n552 ,n404 ,n487);
    not g743(n1954 ,n1953);
    not g744(n2805 ,n2804);
    xor g745(n3308 ,n2978 ,n2988);
    xnor g746(n2602 ,n2478 ,n2380);
    nor g747(n2571 ,n2409 ,n2500);
    nor g748(n1231 ,n1091 ,n1177);
    or g749(n820 ,n720 ,n681);
    buf g750(n13[8], 1'b0);
    not g751(n2423 ,n2422);
    not g752(n668 ,n667);
    nor g753(n1655 ,n1543 ,n1595);
    nor g754(n2448 ,n1931 ,n2346);
    nor g755(n3055 ,n3011 ,n3054);
    not g756(n55 ,n30[0]);
    nor g757(n2758 ,n2679 ,n2695);
    or g758(n549 ,n441 ,n492);
    xor g759(n2256 ,n2014 ,n2077);
    nor g760(n2493 ,n2379 ,n2447);
    nor g761(n2067 ,n1864 ,n1861);
    nor g762(n1973 ,n1887 ,n1876);
    not g763(n2062 ,n2061);
    or g764(n594 ,n423 ,n503);
    xnor g765(n3320 ,n3029 ,n3041);
    nor g766(n2487 ,n2410 ,n2400);
    nor g767(n1163 ,n1054 ,n1117);
    not g768(n1962 ,n1961);
    dff g769(.RN(n1), .SN(1'b1), .CK(n0), .D(n590), .Q(n30[6]));
    xor g770(n940 ,n967 ,n987);
    xor g771(n945 ,n1186 ,n1192);
    nor g772(n3244 ,n3151 ,n3164);
    not g773(n2009 ,n2008);
    or g774(n545 ,n374 ,n456);
    xnor g775(n1235 ,n1026 ,n1136);
    xnor g776(n1423 ,n1374 ,n1348);
    not g777(n2741 ,n2740);
    nor g778(n1568 ,n1521 ,n1534);
    nor g779(n1621 ,n1519 ,n1555);
    nor g780(n1094 ,n1002 ,n1078);
    nor g781(n1838 ,n1812 ,n1825);
    not g782(n172 ,n924);
    buf g783(n12[22], n10[14]);
    xnor g784(n1033 ,n940 ,n1018);
    nor g785(n2547 ,n2375 ,n2510);
    nor g786(n2008 ,n1887 ,n1875);
    not g787(n2964 ,n23[3]);
    not g788(n1703 ,n1702);
    xnor g789(n1776 ,n1707 ,n1745);
    nor g790(n2292 ,n2094 ,n2162);
    nor g791(n751 ,n180 ,n660);
    buf g792(n11[18], n10[2]);
    xnor g793(n1825 ,n1789 ,n1767);
    not g794(n3111 ,n3320);
    nor g795(n1003 ,n957 ,n992);
    nor g796(n470 ,n273 ,n102);
    nor g797(n1331 ,n1259 ,n1306);
    nor g798(n3046 ,n3032 ,n3045);
    or g799(n3229 ,n3190 ,n3211);
    or g800(n608 ,n445 ,n491);
    nor g801(n2284 ,n2041 ,n2220);
    nor g802(n2776 ,n2720 ,n2757);
    buf g803(n10[24], 1'b0);
    xnor g804(n1492 ,n1479 ,n1484);
    nor g805(n477 ,n156 ,n102);
    nor g806(n2515 ,n2344 ,n2418);
    not g807(n142 ,n31[1]);
    nor g808(n2532 ,n2455 ,n2453);
    not g809(n1900 ,n1899);
    nor g810(n1309 ,n1167 ,n1262);
    dff g811(.RN(n1), .SN(1'b1), .CK(n0), .D(n838), .Q(n21[2]));
    not g812(n82 ,n25[1]);
    nor g813(n489 ,n290 ,n102);
    xnor g814(n2888 ,n2821 ,n2847);
    nor g815(n1632 ,n1563 ,n1592);
    nor g816(n977 ,n965 ,n964);
    nor g817(n3149 ,n3076 ,n3100);
    or g818(n597 ,n426 ,n506);
    not g819(n2090 ,n2089);
    not g820(n1866 ,n23[0]);
    or g821(n604 ,n442 ,n490);
    or g822(n843 ,n737 ,n694);
    xnor g823(n2867 ,n2822 ,n2820);
    xnor g824(n2837 ,n2790 ,n2819);
    not g825(n1896 ,n1895);
    or g826(n3248 ,n3178 ,n3238);
    nor g827(n2862 ,n2781 ,n2843);
    xnor g828(n1707 ,n1549 ,n1653);
    nor g829(n713 ,n110 ,n663);
    not g830(n2871 ,n2870);
    nor g831(n2584 ,n2318 ,n2522);
    xnor g832(n1488 ,n1460 ,n1470);
    xnor g833(n2656 ,n2538 ,n2402);
    nor g834(n1850 ,n1834 ,n1849);
    nor g835(n2110 ,n1886 ,n1875);
    nor g836(n2668 ,n2579 ,n2628);
    nor g837(n2546 ,n2374 ,n2525);
    xnor g838(n1836 ,n1808 ,n1793);
    xnor g839(n2769 ,n2691 ,n2636);
    xnor g840(n1151 ,n1029 ,n1043);
    nor g841(n398 ,n253 ,n103);
    not g842(n1946 ,n1945);
    xor g843(n2538 ,n2433 ,n2371);
    or g844(n889 ,n622 ,n813);
    nor g845(n1969 ,n1890 ,n1878);
    nor g846(n2714 ,n2606 ,n2651);
    nor g847(n1678 ,n1657 ,n1632);
    nor g848(n733 ,n215 ,n649);
    or g849(n578 ,n410 ,n515);
    not g850(n127 ,n21[2]);
    nor g851(n510 ,n159 ,n346);
    or g852(n922 ,n30[6] ,n46);
    nor g853(n2924 ,n2886 ,n2906);
    nor g854(n402 ,n246 ,n103);
    or g855(n50 ,n25[6] ,n25[5]);
    buf g856(n13[12], 1'b0);
    not g857(n209 ,n21[5]);
    dff g858(.RN(n1), .SN(1'b1), .CK(n0), .D(n544), .Q(n28[13]));
    nor g859(n1648 ,n1571 ,n1617);
    nor g860(n2675 ,n2534 ,n2588);
    nor g861(n1608 ,n1522 ,n1552);
    nor g862(n1455 ,n1301 ,n1425);
    not g863(n2401 ,n2400);
    not g864(n2851 ,n2850);
    nor g865(n2282 ,n2085 ,n2217);
    not g866(n3082 ,n3300);
    not g867(n3071 ,n32[10]);
    nor g868(n1274 ,n1224 ,n1218);
    or g869(n845 ,n739 ,n696);
    not g870(n1938 ,n1937);
    nor g871(n3210 ,n3069 ,n3155);
    xnor g872(n2257 ,n1929 ,n1905);
    nor g873(n371 ,n265 ,n103);
    nor g874(n1476 ,n1445 ,n1461);
    xnor g875(n3277 ,n2839 ,n2858);
    not g876(n2397 ,n2396);
    xnor g877(n3029 ,n3291 ,n3275);
    xnor g878(n2689 ,n2600 ,n2598);
    nor g879(n1255 ,n1235 ,n1209);
    buf g880(n12[6], 1'b0);
    or g881(n853 ,n746 ,n718);
    nor g882(n1692 ,n1658 ,n1633);
    or g883(n543 ,n372 ,n454);
    nor g884(n1785 ,n1758 ,n1763);
    nor g885(n2228 ,n1978 ,n2009);
    not g886(n145 ,n31[8]);
    not g887(n99 ,n98);
    nor g888(n1800 ,n1768 ,n1774);
    dff g889(.RN(n1), .SN(1'b1), .CK(n0), .D(n549), .Q(n28[7]));
    nor g890(n725 ,n206 ,n651);
    nor g891(n2711 ,n2535 ,n2667);
    or g892(n3160 ,n3154 ,n3134);
    nor g893(n2982 ,n2971 ,n2977);
    xnor g894(n1400 ,n1327 ,n1354);
    nor g895(n1109 ,n948 ,n1064);
    or g896(n32[12] ,n1799 ,n1860);
    not g897(n275 ,n26[10]);
    nor g898(n1264 ,n1148 ,n1240);
    nor g899(n1093 ,n1003 ,n1072);
    nor g900(n2193 ,n1936 ,n1946);
    nor g901(n790 ,n185 ,n652);
    nor g902(n1783 ,n1699 ,n1756);
    nor g903(n1388 ,n1280 ,n1359);
    or g904(n341 ,n294 ,n299);
    not g905(n2405 ,n2404);
    nor g906(n1768 ,n1685 ,n1744);
    nor g907(n2524 ,n2341 ,n2466);
    nor g908(n3187 ,n3070 ,n3155);
    not g909(n1624 ,n1623);
    xnor g910(n2639 ,n2551 ,n2560);
    not g911(n1942 ,n1941);
    or g912(n838 ,n732 ,n691);
    nor g913(n419 ,n284 ,n105);
    xnor g914(n3292 ,n1399 ,n1384);
    nor g915(n1157 ,n1057 ,n1133);
    nor g916(n2358 ,n2226 ,n2274);
    dff g917(.RN(n1), .SN(1'b1), .CK(n0), .D(n839), .Q(n21[1]));
    nor g918(n1822 ,n1793 ,n1808);
    nor g919(n349 ,n108 ,n308);
    xnor g920(n3297 ,n1473 ,n1496);
    or g921(n905 ,n863 ,n862);
    buf g922(n11[8], 1'b0);
    nor g923(n2288 ,n1994 ,n2161);
    buf g924(n9[25], 1'b0);
    not g925(n657 ,n658);
    not g926(n2625 ,n2624);
    nor g927(n710 ,n111 ,n663);
    not g928(n1222 ,n1221);
    not g929(n249 ,n10[9]);
    nor g930(n757 ,n123 ,n658);
    or g931(n1531 ,n1513 ,n1527);
    nor g932(n1502 ,n1476 ,n1501);
    nor g933(n2757 ,n2668 ,n2721);
    xnor g934(n2786 ,n2736 ,n2738);
    nor g935(n2128 ,n1880 ,n1874);
    not g936(n1582 ,n1581);
    xnor g937(n2275 ,n2110 ,n1973);
    or g938(n3156 ,n3154 ,n3130);
    nor g939(n693 ,n114 ,n661);
    nor g940(n2039 ,n1871 ,n1874);
    not g941(n2731 ,n2730);
    or g942(n1040 ,n991 ,n1022);
    not g943(n1891 ,n23[4]);
    nor g944(n968 ,n20[5] ,n21[5]);
    not g945(n268 ,n26[4]);
    buf g946(n12[20], n10[12]);
    nor g947(n2150 ,n2017 ,n2059);
    or g948(n894 ,n768 ,n680);
    nor g949(n1329 ,n1270 ,n1314);
    or g950(n3221 ,n3174 ,n3170);
    nor g951(n471 ,n291 ,n104);
    not g952(n1699 ,n1698);
    xnor g953(n1213 ,n1153 ,n1028);
    nor g954(n440 ,n281 ,n103);
    nor g955(n620 ,n243 ,n524);
    dff g956(.RN(n1), .SN(1'b1), .CK(n0), .D(n892), .Q(n23[1]));
    nor g957(n3040 ,n3028 ,n3039);
    or g958(n3252 ,n3186 ,n3240);
    or g959(n596 ,n425 ,n505);
    dff g960(.RN(n1), .SN(1'b1), .CK(n0), .D(n833), .Q(n21[5]));
    xnor g961(n3294 ,n1439 ,n1472);
    nor g962(n62 ,n58 ,n55);
    or g963(n294 ,n5[29] ,n5[28]);
    nor g964(n1927 ,n1865 ,n1873);
    nor g965(n2516 ,n2372 ,n2402);
    not g966(n1643 ,n1642);
    not g967(n2000 ,n1999);
    not g968(n3001 ,n3272);
    not g969(n1631 ,n1630);
    nor g970(n2900 ,n2834 ,n2863);
    not g971(n1898 ,n1897);
    or g972(n301 ,n7[1] ,n7[0]);
    nor g973(n2077 ,n1885 ,n1866);
    nor g974(n1564 ,n1519 ,n1530);
    nor g975(n2858 ,n2813 ,n2830);
    nor g976(n618 ,n267 ,n524);
    xnor g977(n1223 ,n1030 ,n1163);
    not g978(n1380 ,n1379);
    xnor g979(n1759 ,n1709 ,n1646);
    nor g980(n1567 ,n1521 ,n1536);
    nor g981(n2192 ,n2020 ,n2084);
    nor g982(n1445 ,n1409 ,n1430);
    xor g983(n2236 ,n2114 ,n2045);
    or g984(n915 ,n897 ,n906);
    nor g985(n2525 ,n2334 ,n2392);
    xnor g986(n2821 ,n2763 ,n2775);
    or g987(n872 ,n753 ,n704);
    buf g988(n9[9], 1'b0);
    nor g989(n1275 ,n1234 ,n1208);
    buf g990(n11[15], 1'b0);
    xnor g991(n2451 ,n2265 ,n2097);
    nor g992(n1098 ,n1013 ,n1076);
    dff g993(.RN(n1), .SN(1'b1), .CK(n0), .D(n594), .Q(n10[9]));
    nor g994(n1501 ,n1500 ,n1482);
    not g995(n80 ,n25[4]);
    nor g996(n804 ,n201 ,n666);
    nor g997(n926 ,n97 ,n98);
    nor g998(n1110 ,n947 ,n1063);
    xnor g999(n3024 ,n3296 ,n3280);
    nor g1000(n2719 ,n2499 ,n2646);
    nor g1001(n2779 ,n2663 ,n2744);
    xnor g1002(n2916 ,n2867 ,n2898);
    nor g1003(n2300 ,n1938 ,n2219);
    nor g1004(n1573 ,n1521 ,n1535);
    nor g1005(n1801 ,n1581 ,n1787);
    nor g1006(n2324 ,n2173 ,n2279);
    xor g1007(n2545 ,n2432 ,n2422);
    dff g1008(.RN(n1), .SN(1'b1), .CK(n0), .D(n845), .Q(n20[3]));
    not g1009(n3094 ,n3258);
    not g1010(n2686 ,n2685);
    nor g1011(n695 ,n110 ,n661);
    xnor g1012(n2280 ,n2095 ,n1941);
    xnor g1013(n1367 ,n1293 ,n944);
    or g1014(n865 ,n614 ,n779);
    nor g1015(n1583 ,n1520 ,n1534);
    or g1016(n542 ,n389 ,n457);
    xnor g1017(n1185 ,n1016 ,n1094);
    xnor g1018(n3259 ,n3034 ,n3057);
    or g1019(n300 ,n26[6] ,n26[7]);
    not g1020(n195 ,n22[7]);
    or g1021(n856 ,n749 ,n702);
    not g1022(n273 ,n29[12]);
    nor g1023(n1268 ,n1173 ,n1205);
    nor g1024(n2933 ,n2905 ,n2918);
    xnor g1025(n2788 ,n2648 ,n2758);
    xnor g1026(n1250 ,n1187 ,n1140);
    nor g1027(n2996 ,n2975 ,n2995);
    nor g1028(n3215 ,n3102 ,n3155);
    nor g1029(n1766 ,n1679 ,n1730);
    not g1030(n244 ,n26[0]);
    nor g1031(n748 ,n116 ,n660);
    buf g1032(n11[3], 1'b0);
    nor g1033(n767 ,n221 ,n664);
    nor g1034(n1113 ,n960 ,n1063);
    not g1035(n194 ,n20[1]);
    not g1036(n256 ,n24[7]);
    nor g1037(n2188 ,n2054 ,n2034);
    not g1038(n2454 ,n2453);
    nor g1039(n1307 ,n944 ,n1272);
    not g1040(n2903 ,n2902);
    nor g1041(n1833 ,n1803 ,n1807);
    not g1042(n93 ,n92);
    nor g1043(n2531 ,n2462 ,n2458);
    nor g1044(n2809 ,n2754 ,n2770);
    xnor g1045(n1203 ,n1137 ,n1028);
    not g1046(n153 ,n31[7]);
    nor g1047(n722 ,n217 ,n651);
    xnor g1048(n1233 ,n1026 ,n1139);
    dff g1049(.RN(n1), .SN(1'b1), .CK(n0), .D(n586), .Q(n25[1]));
    dff g1050(.RN(n1), .SN(1'b1), .CK(n0), .D(n851), .Q(n19[5]));
    nor g1051(n1599 ,n1519 ,n1554);
    nor g1052(n769 ,n180 ,n652);
    nor g1053(n974 ,n20[6] ,n20[5]);
    nor g1054(n1435 ,n1378 ,n1412);
    nor g1055(n729 ,n209 ,n649);
    nor g1056(n1497 ,n1469 ,n1496);
    not g1057(n212 ,n28[0]);
    not g1058(n1990 ,n1989);
    not g1059(n991 ,n992);
    not g1060(n1865 ,n20[1]);
    or g1061(n567 ,n407 ,n464);
    nor g1062(n3213 ,n3101 ,n3155);
    not g1063(n169 ,n935);
    not g1064(n1353 ,n1352);
    nor g1065(n2622 ,n2582 ,n2505);
    nor g1066(n1475 ,n1470 ,n1459);
    not g1067(n2036 ,n2035);
    or g1068(n323 ,n118 ,n115);
    not g1069(n966 ,n20[2]);
    nor g1070(n364 ,n344 ,n345);
    xnor g1071(n2453 ,n2238 ,n2099);
    nor g1072(n105 ,n184 ,n319);
    nor g1073(n2053 ,n1865 ,n1881);
    not g1074(n2629 ,n2628);
    xnor g1075(n1221 ,n1029 ,n1160);
    nor g1076(n2164 ,n1893 ,n2045);
    xnor g1077(n1808 ,n1769 ,n1753);
    xnor g1078(n2273 ,n1979 ,n2128);
    not g1079(n3087 ,n3295);
    not g1080(n60 ,n30[2]);
    xnor g1081(n1374 ,n1325 ,n1330);
    nor g1082(n3208 ,n3081 ,n3155);
    buf g1083(n9[26], 1'b0);
    nor g1084(n3200 ,n3089 ,n3154);
    nor g1085(n1450 ,n1415 ,n1421);
    nor g1086(n717 ,n106 ,n668);
    nor g1087(n1162 ,n1048 ,n1131);
    xnor g1088(n2476 ,n2269 ,n2365);
    nor g1089(n747 ,n188 ,n660);
    not g1090(n963 ,n21[6]);
    buf g1091(n13[13], 1'b0);
    not g1092(n1794 ,n1793);
    buf g1093(n12[31], 1'b0);
    nor g1094(n465 ,n162 ,n102);
    xnor g1095(n3027 ,n3297 ,n3281);
    not g1096(n2429 ,n2428);
    xor g1097(n3265 ,n20[1] ,n21[1]);
    nor g1098(n1142 ,n1044 ,n1110);
    nor g1099(n2830 ,n2784 ,n2812);
    nor g1100(n1931 ,n1892 ,n1868);
    xnor g1101(n2240 ,n2035 ,n1947);
    buf g1102(n9[30], 1'b0);
    xnor g1103(n2704 ,n2586 ,n2635);
    nor g1104(n1684 ,n1636 ,n1644);
    or g1105(n900 ,n814 ,n889);
    not g1106(n137 ,n5[4]);
    nor g1107(n779 ,n129 ,n665);
    or g1108(n883 ,n761 ,n710);
    not g1109(n2344 ,n2343);
    nor g1110(n1276 ,n1236 ,n1210);
    nor g1111(n2517 ,n2338 ,n2412);
    not g1112(n1890 ,n21[4]);
    or g1113(n909 ,n865 ,n828);
    dff g1114(.RN(n1), .SN(1'b1), .CK(n0), .D(n842), .Q(n20[6]));
    nor g1115(n37 ,n35 ,n34);
    nor g1116(n1667 ,n1572 ,n1609);
    not g1117(n188 ,n19[5]);
    nor g1118(n3237 ,n3145 ,n3157);
    or g1119(n3154 ,n3099 ,n3067);
    nor g1120(n2155 ,n1923 ,n2057);
    nor g1121(n990 ,n963 ,n974);
    or g1122(n1985 ,n1884 ,n1862);
    xnor g1123(n1358 ,n1291 ,n1206);
    nor g1124(n1505 ,n1504 ,n1481);
    nor g1125(n1079 ,n948 ,n1032);
    not g1126(n2909 ,n2908);
    nor g1127(n3146 ,n3111 ,n3072);
    or g1128(n31[14] ,n3168 ,n3230);
    nor g1129(n721 ,n128 ,n651);
    not g1130(n949 ,n3306);
    buf g1131(n9[8], 1'b0);
    dff g1132(.RN(n1), .SN(1'b1), .CK(n0), .D(n873), .Q(n24[6]));
    nor g1133(n61 ,n30[1] ,n30[0]);
    not g1134(n2005 ,n2004);
    xnor g1135(n1296 ,n1224 ,n941);
    nor g1136(n2158 ,n2019 ,n2083);
    xnor g1137(n1028 ,n1006 ,n993);
    nor g1138(n3193 ,n3121 ,n3154);
    not g1139(n262 ,n28[13]);
    nor g1140(n2576 ,n2433 ,n2516);
    nor g1141(n1323 ,n1320 ,n1276);
    not g1142(n134 ,n31[15]);
    nor g1143(n2699 ,n2634 ,n2672);
    nor g1144(n1700 ,n1602 ,n1670);
    xnor g1145(n1555 ,n3269 ,n23[5]);
    nor g1146(n1133 ,n956 ,n1062);
    nor g1147(n704 ,n111 ,n657);
    or g1148(n3157 ,n3154 ,n3131);
    xnor g1149(n2840 ,n2806 ,n2481);
    not g1150(n2127 ,n2126);
    buf g1151(n11[30], n10[14]);
    or g1152(n574 ,n408 ,n481);
    not g1153(n1526 ,n3269);
    nor g1154(n731 ,n201 ,n649);
    nor g1155(n1967 ,n1887 ,n1877);
    nor g1156(n3207 ,n3068 ,n3155);
    not g1157(n962 ,n20[5]);
    nor g1158(n2902 ,n2873 ,n2897);
    not g1159(n1560 ,n1559);
    nor g1160(n1529 ,n3270 ,n23[6]);
    or g1161(n630 ,n339 ,n626);
    not g1162(n1515 ,n23[2]);
    not g1163(n180 ,n19[1]);
    nor g1164(n1430 ,n1369 ,n1410);
    xnor g1165(n2471 ,n2235 ,n2279);
    dff g1166(.RN(n1), .SN(1'b1), .CK(n0), .D(n538), .Q(n29[4]));
    nor g1167(n429 ,n247 ,n105);
    not g1168(n2052 ,n2051);
    or g1169(n840 ,n734 ,n672);
    or g1170(n583 ,n412 ,n517);
    not g1171(n1234 ,n1233);
    not g1172(n2627 ,n2626);
    not g1173(n235 ,n10[8]);
    not g1174(n280 ,n26[6]);
    nor g1175(n3198 ,n3117 ,n3141);
    nor g1176(n428 ,n141 ,n347);
    not g1177(n272 ,n26[12]);
    dff g1178(.RN(n1), .SN(1'b1), .CK(n0), .D(n570), .Q(n14));
    nor g1179(n2626 ,n2508 ,n2568);
    nor g1180(n1957 ,n1885 ,n1868);
    nor g1181(n2971 ,n2960 ,n2961);
    nor g1182(n2949 ,n2948 ,n2932);
    nor g1183(n442 ,n286 ,n103);
    nor g1184(n2293 ,n2105 ,n2166);
    not g1185(n1641 ,n1640);
    nor g1186(n1627 ,n1577 ,n1621);
    dff g1187(.RN(n1), .SN(1'b1), .CK(n0), .D(n576), .Q(n26[0]));
    nor g1188(n3134 ,n3321 ,n32[4]);
    not g1189(n2050 ,n2049);
    not g1190(n83 ,n25[5]);
    xnor g1191(n2260 ,n1913 ,n2029);
    or g1192(n540 ,n380 ,n353);
    xnor g1193(n1205 ,n1029 ,n1162);
    not g1194(n1214 ,n1213);
    xnor g1195(n2245 ,n2061 ,n2043);
    nor g1196(n1477 ,n1431 ,n1472);
    nor g1197(n389 ,n278 ,n105);
    nor g1198(n807 ,n218 ,n665);
    nor g1199(n2780 ,n2739 ,n2737);
    or g1200(n916 ,n900 ,n895);
    not g1201(n215 ,n21[1]);
    xnor g1202(n1717 ,n1647 ,n1623);
    or g1203(n554 ,n395 ,n358);
    dff g1204(.RN(n1), .SN(1'b1), .CK(n0), .D(n542), .Q(n29[13]));
    nor g1205(n1650 ,n1580 ,n1600);
    not g1206(n348 ,n349);
    nor g1207(n2835 ,n2735 ,n2794);
    xnor g1208(n1706 ,n1659 ,n1661);
    nor g1209(n1431 ,n1341 ,n1402);
    or g1210(n310 ,n5[13] ,n5[12]);
    xnor g1211(n2587 ,n2398 ,n2535);
    not g1212(n3092 ,n3288);
    nor g1213(n2678 ,n2399 ,n2595);
    nor g1214(n690 ,n113 ,n648);
    nor g1215(n1506 ,n1475 ,n1505);
    not g1216(n236 ,n26[7]);
    nor g1217(n1137 ,n1060 ,n1106);
    nor g1218(n2159 ,n2047 ,n2089);
    nor g1219(n435 ,n212 ,n103);
    nor g1220(n481 ,n148 ,n104);
    nor g1221(n353 ,n104 ,n328);
    not g1222(n2458 ,n2457);
    nor g1223(n1859 ,n1831 ,n1858);
    or g1224(n653 ,n523 ,n644);
    or g1225(n3223 ,n3180 ,n3177);
    not g1226(n2801 ,n2800);
    xnor g1227(n2824 ,n2773 ,n2683);
    dff g1228(.RN(n1), .SN(1'b1), .CK(n0), .D(n877), .Q(n24[3]));
    nor g1229(n2317 ,n2102 ,n2171);
    nor g1230(n2441 ,n2373 ,n2363);
    nor g1231(n1593 ,n1522 ,n1555);
    or g1232(n572 ,n406 ,n478);
    nor g1233(n3017 ,n2997 ,n2999);
    nor g1234(n2742 ,n2645 ,n2694);
    nor g1235(n2815 ,n2703 ,n2772);
    not g1236(n2116 ,n2115);
    not g1237(n2848 ,n2847);
    xnor g1238(n2592 ,n2472 ,n2396);
    xor g1239(n2433 ,n2241 ,n2135);
    buf g1240(n13[30], n10[6]);
    nor g1241(n2910 ,n2878 ,n2900);
    dff g1242(.RN(n1), .SN(1'b1), .CK(n0), .D(n841), .Q(n20[7]));
    nor g1243(n3195 ,n3088 ,n3141);
    nor g1244(n1744 ,n1695 ,n1716);
    xor g1245(n3261 ,n3037 ,n3062);
    dff g1246(.RN(n1), .SN(1'b1), .CK(n0), .D(n912), .Q(n9[6]));
    nor g1247(n2174 ,n2053 ,n2033);
    not g1248(n120 ,n21[0]);
    nor g1249(n1609 ,n1521 ,n1554);
    nor g1250(n1167 ,n1073 ,n1122);
    dff g1251(.RN(n1), .SN(1'b1), .CK(n0), .D(n554), .Q(n29[0]));
    xnor g1252(n1447 ,n1400 ,n1370);
    nor g1253(n423 ,n249 ,n347);
    not g1254(n189 ,n27[1]);
    not g1255(n1994 ,n1993);
    nor g1256(n2180 ,n2043 ,n2061);
    nor g1257(n2738 ,n2670 ,n2693);
    nor g1258(n1830 ,n1776 ,n1811);
    not g1259(n955 ,n20[0]);
    xnor g1260(n336 ,n212 ,n187);
    xnor g1261(n1287 ,n1207 ,n1233);
    nor g1262(n2665 ,n2584 ,n2616);
    or g1263(n571 ,n377 ,n477);
    or g1264(n631 ,n338 ,n624);
    or g1265(n311 ,n5[25] ,n5[24]);
    nor g1266(n1103 ,n948 ,n1063);
    not g1267(n187 ,n19[0]);
    nor g1268(n2017 ,n1886 ,n1881);
    buf g1269(n12[2], 1'b0);
    nor g1270(n1420 ,n1297 ,n1404);
    buf g1271(n13[3], 1'b0);
    nor g1272(n2087 ,n1890 ,n1889);
    xnor g1273(n526 ,n104 ,n30[0]);
    dff g1274(.RN(n1), .SN(1'b1), .CK(n0), .D(n625), .Q(n15));
    not g1275(n1970 ,n1969);
    nor g1276(n1465 ,n1427 ,n1443);
    nor g1277(n1272 ,n1211 ,n1214);
    buf g1278(n13[19], 1'b0);
    buf g1279(n9[31], 1'b0);
    or g1280(n49 ,n25[3] ,n25[2]);
    nor g1281(n2321 ,n2123 ,n2156);
    not g1282(n1426 ,n1425);
    xor g1283(n3263 ,n3023 ,n3066);
    not g1284(n2002 ,n2001);
    nor g1285(n2526 ,n2460 ,n2395);
    nor g1286(n2353 ,n2160 ,n2312);
    nor g1287(n1636 ,n1570 ,n1608);
    nor g1288(n1963 ,n1863 ,n1889);
    not g1289(n650 ,n651);
    not g1290(n2534 ,n2533);
    not g1291(n190 ,n24[2]);
    not g1292(n1877 ,n22[3]);
    nor g1293(n1092 ,n1014 ,n1085);
    nor g1294(n1410 ,n1379 ,n1357);
    nor g1295(n1630 ,n1540 ,n1614);
    nor g1296(n2133 ,n1885 ,n1891);
    not g1297(n1509 ,n3265);
    nor g1298(n2967 ,n22[7] ,n23[7]);
    not g1299(n128 ,n22[5]);
    nor g1300(n1159 ,n1058 ,n1118);
    or g1301(n1062 ,n1023 ,n1037);
    not g1302(n1444 ,n1443);
    nor g1303(n1743 ,n1691 ,n1718);
    nor g1304(n2968 ,n22[6] ,n23[6]);
    nor g1305(n1259 ,n1168 ,n1202);
    nor g1306(n2120 ,n1863 ,n1862);
    not g1307(n2330 ,n2329);
    not g1308(n251 ,n25[6]);
    nor g1309(n1685 ,n1661 ,n1659);
    nor g1310(n764 ,n214 ,n664);
    not g1311(n2028 ,n2027);
    xnor g1312(n2551 ,n2386 ,n2222);
    nor g1313(n2124 ,n1880 ,n1876);
    nor g1314(n2672 ,n2613 ,n2608);
    not g1315(n1302 ,n1301);
    nor g1316(n444 ,n156 ,n103);
    or g1317(n576 ,n399 ,n483);
    nor g1318(n2122 ,n1884 ,n1888);
    or g1319(n823 ,n722 ,n683);
    or g1320(n921 ,n50 ,n53);
    nor g1321(n1612 ,n1522 ,n1554);
    nor g1322(n679 ,n106 ,n663);
    nor g1323(n802 ,n116 ,n652);
    xnor g1324(n1557 ,n3265 ,n23[1]);
    nor g1325(n1691 ,n1637 ,n1645);
    nor g1326(n815 ,n220 ,n653);
    nor g1327(n1923 ,n1887 ,n1873);
    xnor g1328(n3032 ,n3293 ,n3277);
    not g1329(n266 ,n29[9]);
    or g1330(n317 ,n5[19] ,n5[18]);
    nor g1331(n1161 ,n1045 ,n1100);
    nor g1332(n2360 ,n2228 ,n2276);
    nor g1333(n1596 ,n1522 ,n1558);
    xnor g1334(n1790 ,n1751 ,n1725);
    buf g1335(n9[15], 1'b0);
    xnor g1336(n2242 ,n2027 ,n1895);
    nor g1337(n1503 ,n1491 ,n1502);
    xnor g1338(n2850 ,n2786 ,n2804);
    nor g1339(n496 ,n289 ,n105);
    xnor g1340(n1291 ,n1174 ,n1244);
    not g1341(n2413 ,n2412);
    nor g1342(n2376 ,n2207 ,n2287);
    nor g1343(n1132 ,n949 ,n1064);
    not g1344(n1403 ,n1402);
    not g1345(n269 ,n26[14]);
    not g1346(n206 ,n22[1]);
    nor g1347(n1681 ,n1626 ,n1669);
    nor g1348(n810 ,n127 ,n666);
    or g1349(n313 ,n5[31] ,n5[30]);
    or g1350(n827 ,n621 ,n772);
    nor g1351(n1407 ,n1388 ,n1384);
    not g1352(n231 ,n9[0]);
    or g1353(n561 ,n401 ,n470);
    or g1354(n581 ,n411 ,n514);
    xnor g1355(n32[5] ,n1835 ,n1840);
    or g1356(n580 ,n416 ,n516);
    nor g1357(n762 ,n197 ,n664);
    nor g1358(n2854 ,n2816 ,n2827);
    or g1359(n654 ,n323 ,n643);
    or g1360(n36 ,n30[6] ,n30[5]);
    not g1361(n1796 ,n1795);
    nor g1362(n38 ,n33 ,n37);
    xnor g1363(n2771 ,n2689 ,n2633);
    nor g1364(n1720 ,n1646 ,n1692);
    xnor g1365(n1175 ,n1017 ,n1097);
    xnor g1366(n1770 ,n1733 ,n1731);
    nor g1367(n2444 ,n2269 ,n2365);
    or g1368(n532 ,n387 ,n450);
    not g1369(n2123 ,n2122);
    or g1370(n1556 ,n1537 ,n1529);
    nor g1371(n814 ,n186 ,n652);
    nor g1372(n2507 ,n2353 ,n2442);
    xnor g1373(n2383 ,n2267 ,n2224);
    or g1374(n2003 ,n1882 ,n1878);
    not g1375(n3088 ,n3297);
    nor g1376(n2335 ,n2213 ,n2309);
    nor g1377(n808 ,n182 ,n652);
    xnor g1378(n3311 ,n2975 ,n2995);
    nor g1379(n445 ,n165 ,n103);
    or g1380(n854 ,n748 ,n701);
    nor g1381(n1694 ,n1629 ,n1643);
    not g1382(n240 ,n24[4]);
    buf g1383(n17[7], 1'b0);
    not g1384(n3080 ,n3302);
    nor g1385(n2316 ,n1992 ,n2150);
    xnor g1386(n1443 ,n1396 ,n1350);
    not g1387(n3128 ,n3299);
    xnor g1388(n1198 ,n1030 ,n1114);
    not g1389(n947 ,n3308);
    not g1390(n108 ,n18[2]);
    nor g1391(n2484 ,n2354 ,n2439);
    buf g1392(n10[25], 1'b0);
    xor g1393(n3269 ,n20[5] ,n21[5]);
    xnor g1394(n2406 ,n2247 ,n2006);
    not g1395(n3076 ,n3313);
    nor g1396(n2761 ,n2738 ,n2736);
    dff g1397(.RN(n1), .SN(1'b1), .CK(n0), .D(n600), .Q(n10[3]));
    or g1398(n537 ,n434 ,n354);
    not g1399(n131 ,n3);
    nor g1400(n735 ,n205 ,n662);
    not g1401(n1870 ,n23[3]);
    nor g1402(n1088 ,n946 ,n1040);
    buf g1403(n12[8], n10[0]);
    nor g1404(n479 ,n271 ,n102);
    nor g1405(n91 ,n25[3] ,n89);
    nor g1406(n2943 ,n2942 ,n2926);
    nor g1407(n1366 ,n1266 ,n1343);
    not g1408(n2336 ,n2335);
    buf g1409(n11[20], n10[4]);
    xnor g1410(n1350 ,n1288 ,n1320);
    nor g1411(n1304 ,n1167 ,n1284);
    nor g1412(n1344 ,n1261 ,n1315);
    or g1413(n831 ,n727 ,n686);
    xnor g1414(n2541 ,n2455 ,n2453);
    or g1415(n3256 ,n3202 ,n3232);
    dff g1416(.RN(n1), .SN(1'b1), .CK(n0), .D(n558), .Q(n17[3]));
    not g1417(n1664 ,n1663);
    nor g1418(n2190 ,n1972 ,n1958);
    dff g1419(.RN(n1), .SN(1'b1), .CK(n0), .D(n608), .Q(n30[3]));
    nor g1420(n1628 ,n1565 ,n1596);
    not g1421(n2774 ,n2773);
    nor g1422(n1394 ,n1339 ,n1368);
    nor g1423(n803 ,n211 ,n655);
    xnor g1424(n1478 ,n1438 ,n1395);
    xor g1425(n2255 ,n2103 ,n1951);
    nor g1426(n2350 ,n2187 ,n2321);
    not g1427(n2102 ,n2101);
    xnor g1428(n2479 ,n2355 ,n2343);
    not g1429(n260 ,n14);
    not g1430(n138 ,n31[3]);
    not g1431(n1873 ,n22[5]);
    nor g1432(n2365 ,n2183 ,n2295);
    nor g1433(n2606 ,n2527 ,n2548);
    not g1434(n1996 ,n1995);
    not g1435(n1863 ,n21[6]);
    nor g1436(n1411 ,n1303 ,n1381);
    not g1437(n1892 ,n21[7]);
    nor g1438(n2514 ,n2370 ,n2414);
    nor g1439(n2530 ,n2456 ,n2454);
    nor g1440(n2315 ,n1996 ,n2148);
    not g1441(n2022 ,n2021);
    nor g1442(n2179 ,n1918 ,n1926);
    not g1443(n277 ,n10[2]);
    buf g1444(n11[0], 1'b0);
    nor g1445(n1620 ,n1520 ,n1553);
    dff g1446(.RN(n1), .SN(1'b1), .CK(n0), .D(n855), .Q(n19[1]));
    xnor g1447(n2428 ,n2254 ,n1903);
    nor g1448(n2970 ,n2963 ,n2964);
    not g1449(n3120 ,n3259);
    not g1450(n1485 ,n1484);
    or g1451(n322 ,n5[3] ,n5[2]);
    not g1452(n3124 ,n3275);
    not g1453(n109 ,n6[2]);
    nor g1454(n1060 ,n956 ,n1034);
    nor g1455(n1340 ,n1258 ,n1307);
    nor g1456(n772 ,n194 ,n665);
    not g1457(n2409 ,n2408);
    nor g1458(n2492 ,n2461 ,n2457);
    nor g1459(n2674 ,n2599 ,n2600);
    not g1460(n164 ,n16);
    nor g1461(n493 ,n170 ,n104);
    nor g1462(n2568 ,n2471 ,n2489);
    xor g1463(n2642 ,n2554 ,n2468);
    nor g1464(n3312 ,n2967 ,n2996);
    or g1465(n2117 ,n1890 ,n1868);
    nor g1466(n2144 ,n1897 ,n1949);
    nor g1467(n518 ,n177 ,n348);
    nor g1468(n410 ,n250 ,n349);
    not g1469(n165 ,n30[3]);
    not g1470(n226 ,n26[5]);
    nor g1471(n2031 ,n1879 ,n1866);
    dff g1472(.RN(n1), .SN(1'b1), .CK(n0), .D(n532), .Q(n28[11]));
    nor g1473(n355 ,n104 ,n329);
    or g1474(n864 ,n617 ,n789);
    dff g1475(.RN(n1), .SN(1'b1), .CK(n0), .D(n529), .Q(n29[15]));
    nor g1476(n699 ,n114 ,n659);
    or g1477(n849 ,n706 ,n698);
    nor g1478(n2355 ,n2198 ,n2301);
    nor g1479(n1145 ,n1083 ,n1103);
    nor g1480(n1781 ,n1701 ,n1748);
    nor g1481(n2716 ,n2611 ,n2658);
    nor g1482(n441 ,n198 ,n105);
    nor g1483(n3153 ,n3077 ,n3068);
    nor g1484(n3201 ,n3078 ,n3142);
    xnor g1485(n2459 ,n2239 ,n1983);
    nor g1486(n1649 ,n1568 ,n1590);
    nor g1487(n1470 ,n1420 ,n1451);
    nor g1488(n1141 ,n1077 ,n1128);
    or g1489(n564 ,n393 ,n472);
    nor g1490(n1068 ,n947 ,n1032);
    nor g1491(n1590 ,n1520 ,n1555);
    nor g1492(n1725 ,n1650 ,n1681);
    buf g1493(n12[14], n10[6]);
    or g1494(n3142 ,n3067 ,n27[1]);
    not g1495(n175 ,n925);
    not g1496(n2559 ,n2558);
    nor g1497(n1780 ,n1726 ,n1751);
    nor g1498(n2173 ,n1935 ,n1945);
    xor g1499(n3268 ,n20[4] ,n21[4]);
    nor g1500(n3236 ,n3144 ,n3156);
    not g1501(n1510 ,n3271);
    buf g1502(n12[13], n10[5]);
    not g1503(n961 ,n21[4]);
    xnor g1504(n1207 ,n1158 ,n1028);
    nor g1505(n925 ,n100 ,n101);
    nor g1506(n2895 ,n2860 ,n2876);
    nor g1507(n2572 ,n2417 ,n2502);
    nor g1508(n1252 ,n1189 ,n1243);
    nor g1509(n3173 ,n3122 ,n3142);
    nor g1510(n511 ,n142 ,n346);
    nor g1511(n1607 ,n1520 ,n1558);
    nor g1512(n2745 ,n2649 ,n2705);
    not g1513(n270 ,n28[14]);
    nor g1514(n376 ,n273 ,n105);
    buf g1515(n13[2], 1'b0);
    not g1516(n2739 ,n2738);
    xnor g1517(n1461 ,n1417 ,n1425);
    nor g1518(n1597 ,n1519 ,n1556);
    not g1519(n1580 ,n1579);
    nor g1520(n1409 ,n1380 ,n1356);
    nor g1521(n811 ,n190 ,n653);
    dff g1522(.RN(n1), .SN(1'b1), .CK(n0), .D(n550), .Q(n30[5]));
    nor g1523(n1045 ,n946 ,n1038);
    nor g1524(n396 ,n225 ,n105);
    nor g1525(n1314 ,n1247 ,n1257);
    nor g1526(n524 ,n131 ,n346);
    nor g1527(n3257 ,n1519 ,n1553);
    xor g1528(n32[9] ,n1847 ,n1855);
    nor g1529(n701 ,n110 ,n659);
    or g1530(n31[13] ,n3184 ,n3222);
    or g1531(n655 ,n325 ,n643);
    not g1532(n2216 ,n2217);
    xnor g1533(n1791 ,n1755 ,n1698);
    nor g1534(n1702 ,n1606 ,n1671);
    nor g1535(n788 ,n197 ,n654);
    nor g1536(n384 ,n255 ,n103);
    nor g1537(n495 ,n117 ,n346);
    nor g1538(n3065 ,n3036 ,n3064);
    nor g1539(n2673 ,n2612 ,n2609);
    nor g1540(n2931 ,n2913 ,n2928);
    not g1541(n1736 ,n1735);
    not g1542(n1672 ,n1671);
    not g1543(n1372 ,n1371);
    nor g1544(n1742 ,n1655 ,n1714);
    nor g1545(n2012 ,n1867 ,n1874);
    not g1546(n1972 ,n1971);
    nor g1547(n1854 ,n1841 ,n1853);
    nor g1548(n2676 ,n2533 ,n2589);
    xnor g1549(n3314 ,n3027 ,n3053);
    not g1550(n1518 ,n23[0]);
    nor g1551(n3232 ,n3153 ,n3165);
    not g1552(n267 ,n9[5]);
    or g1553(n31[10] ,n3221 ,n3247);
    not g1554(n2613 ,n2612);
    nor g1555(n3181 ,n3124 ,n3142);
    nor g1556(n1392 ,n1328 ,n1355);
    dff g1557(.RN(n1), .SN(1'b1), .CK(n0), .D(n577), .Q(n30[7]));
    nor g1558(n1469 ,n1428 ,n1444);
    nor g1559(n2135 ,n1885 ,n1862);
    or g1560(n536 ,n373 ,n489);
    nor g1561(n2633 ,n2531 ,n2565);
    xnor g1562(n2804 ,n2729 ,n2606);
    dff g1563(.RN(n1), .SN(1'b1), .CK(n0), .D(n597), .Q(n10[6]));
    or g1564(n595 ,n424 ,n504);
    or g1565(n333 ,n18[2] ,n307);
    nor g1566(n3189 ,n3093 ,n3141);
    nor g1567(n2880 ,n2803 ,n2857);
    xnor g1568(n2938 ,n2918 ,n2904);
    not g1569(n1576 ,n1575);
    xnor g1570(n987 ,n961 ,n20[4]);
    nor g1571(n3057 ,n3010 ,n3056);
    buf g1572(n11[12], 1'b0);
    not g1573(n2326 ,n2325);
    nor g1574(n1376 ,n1327 ,n1354);
    nor g1575(n2210 ,n1896 ,n2028);
    not g1576(n2268 ,n2267);
    or g1577(n41 ,n30[4] ,n30[3]);
    buf g1578(n11[10], 1'b0);
    nor g1579(n2989 ,n2978 ,n2988);
    xor g1580(n2266 ,n1988 ,n1897);
    not g1581(n3095 ,n3289);
    nor g1582(n2207 ,n1922 ,n1952);
    nor g1583(n1453 ,n1302 ,n1426);
    xnor g1584(n2461 ,n2240 ,n2137);
    nor g1585(n1903 ,n1869 ,n1866);
    nor g1586(n2185 ,n1908 ,n2064);
    nor g1587(n2203 ,n1944 ,n2076);
    nor g1588(n497 ,n134 ,n346);
    nor g1589(n2147 ,n2015 ,n2139);
    not g1590(n232 ,n29[8]);
    nor g1591(n774 ,n199 ,n654);
    nor g1592(n2369 ,n2215 ,n2306);
    nor g1593(n2563 ,n2355 ,n2515);
    or g1594(n665 ,n322 ,n643);
    or g1595(n873 ,n754 ,n705);
    dff g1596(.RN(n1), .SN(1'b1), .CK(n0), .D(n858), .Q(n19[0]));
    nor g1597(n967 ,n20[3] ,n21[3]);
    nor g1598(n1008 ,n979 ,n998);
    not g1599(n1924 ,n1923);
    nor g1600(n1324 ,n1264 ,n1318);
    nor g1601(n1134 ,n1086 ,n1129);
    or g1602(n623 ,n409 ,n482);
    xnor g1603(n2885 ,n2850 ,n2792);
    nor g1604(n486 ,n166 ,n102);
    or g1605(n293 ,n18[1] ,n2);
    nor g1606(n1592 ,n1520 ,n1557);
    xnor g1607(n2920 ,n2884 ,n2860);
    nor g1608(n1427 ,n1389 ,n1401);
    xnor g1609(n1835 ,n1806 ,n1803);
    nor g1610(n2667 ,n2398 ,n2594);
    nor g1611(n1128 ,n959 ,n1063);
    xnor g1612(n1821 ,n1795 ,n1764);
    not g1613(n170 ,n934);
    nor g1614(n2985 ,n2980 ,n2984);
    nor g1615(n1644 ,n1547 ,n1615);
    xnor g1616(n2561 ,n2382 ,n2378);
    dff g1617(.RN(n1), .SN(1'b1), .CK(n0), .D(n596), .Q(n10[7]));
    xnor g1618(n1181 ,n1016 ,n1096);
    nor g1619(n2827 ,n2809 ,n2820);
    nor g1620(n1135 ,n1082 ,n1109);
    nor g1621(n2298 ,n2007 ,n2154);
    not g1622(n3075 ,n3319);
    not g1623(n2229 ,n2228);
    dff g1624(.RN(n1), .SN(1'b1), .CK(n0), .D(n546), .Q(n28[10]));
    nor g1625(n1332 ,n1254 ,n1313);
    nor g1626(n490 ,n171 ,n102);
    not g1627(n3005 ,n3285);
    xnor g1628(n2728 ,n2610 ,n2658);
    or g1629(n639 ,n632 ,n636);
    xnor g1630(n1297 ,n1239 ,n1172);
    xnor g1631(n1243 ,n1026 ,n1134);
    or g1632(n1535 ,n1510 ,n1517);
    not g1633(n2411 ,n2410);
    nor g1634(n975 ,n952 ,n962);
    nor g1635(n1778 ,n1742 ,n1761);
    nor g1636(n3009 ,n3289 ,n3273);
    nor g1637(n3175 ,n3126 ,n3142);
    nor g1638(n928 ,n91 ,n92);
    nor g1639(n417 ,n227 ,n347);
    not g1640(n2655 ,n2654);
    nor g1641(n1306 ,n1149 ,n1279);
    not g1642(n225 ,n29[14]);
    nor g1643(n711 ,n114 ,n663);
    nor g1644(n3050 ,n3025 ,n3049);
    nor g1645(n1468 ,n1383 ,n1453);
    or g1646(n613 ,n342 ,n365);
    nor g1647(n660 ,n525 ,n647);
    xnor g1648(n2838 ,n2798 ,n2730);
    nor g1649(n2817 ,n2696 ,n2776);
    nor g1650(n2319 ,n2032 ,n2223);
    not g1651(n2131 ,n2130);
    or g1652(n877 ,n757 ,n708);
    nor g1653(n65 ,n60 ,n63);
    not g1654(n2756 ,n2755);
    not g1655(n1527 ,n23[3]);
    nor g1656(n387 ,n290 ,n103);
    xnor g1657(n2463 ,n2280 ,n1901);
    buf g1658(n13[18], 1'b0);
    nor g1659(n2198 ,n2070 ,n2072);
    nor g1660(n673 ,n106 ,n661);
    nor g1661(n1663 ,n1566 ,n1593);
    nor g1662(n1260 ,n1180 ,n1237);
    nor g1663(n74 ,n59 ,n72);
    not g1664(n1524 ,n23[4]);
    nor g1665(n1653 ,n1573 ,n1619);
    nor g1666(n407 ,n121 ,n103);
    or g1667(n624 ,n302 ,n610);
    xnor g1668(n3301 ,n1488 ,n1504);
    nor g1669(n483 ,n242 ,n102);
    nor g1670(n2944 ,n2933 ,n2943);
    nor g1671(n2283 ,n1937 ,n2218);
    nor g1672(n2006 ,n1879 ,n1862);
    nor g1673(n3145 ,n3110 ,n3102);
    nor g1674(n2954 ,n2879 ,n2953);
    nor g1675(n3016 ,n3296 ,n3280);
    nor g1676(n88 ,n25[2] ,n86);
    nor g1677(n2339 ,n2178 ,n2307);
    xnor g1678(n2244 ,n2049 ,n1915);
    dff g1679(.RN(n1), .SN(1'b1), .CK(n0), .D(n604), .Q(n30[2]));
    not g1680(n1950 ,n1949);
    nor g1681(n2829 ,n2706 ,n2814);
    nor g1682(n1851 ,n1822 ,n1850);
    nor g1683(n2583 ,n2450 ,n2484);
    nor g1684(n2936 ,n2911 ,n2921);
    not g1685(n2842 ,n2841);
    or g1686(n303 ,n26[8] ,n26[9]);
    nor g1687(n1270 ,n1181 ,n1232);
    nor g1688(n2833 ,n2756 ,n2796);
    not g1689(n79 ,n25[0]);
    xnor g1690(n1746 ,n1713 ,n1655);
    nor g1691(n1441 ,n1411 ,n1432);
    or g1692(n914 ,n909 ,n903);
    not g1693(n1980 ,n1979);
    nor g1694(n499 ,n133 ,n346);
    not g1695(n979 ,n978);
    nor g1696(n3206 ,n3103 ,n3155);
    xnor g1697(n2726 ,n2652 ,n2626);
    xnor g1698(n1149 ,n1017 ,n1067);
    or g1699(n869 ,n798 ,n797);
    nor g1700(n2808 ,n2751 ,n2767);
    or g1701(n3217 ,n3167 ,n3204);
    nor g1702(n1070 ,n956 ,n1032);
    not g1703(n81 ,n25[3]);
    buf g1704(n12[17], n10[9]);
    xnor g1705(n1152 ,n1027 ,n1042);
    not g1706(n1726 ,n1725);
    xnor g1707(n1845 ,n1825 ,n1812);
    nor g1708(n1615 ,n1521 ,n1557);
    nor g1709(n2083 ,n1864 ,n1881);
    nor g1710(n2214 ,n1956 ,n1964);
    nor g1711(n1724 ,n1705 ,n1686);
    nor g1712(n3053 ,n3016 ,n3052);
    nor g1713(n397 ,n155 ,n103);
    or g1714(n34 ,n30[1] ,n30[0]);
    nor g1715(n1129 ,n959 ,n1062);
    xnor g1716(n1551 ,n3267 ,n23[3]);
    nor g1717(n2904 ,n2875 ,n2894);
    nor g1718(n691 ,n109 ,n648);
    dff g1719(.RN(n1), .SN(1'b1), .CK(n0), .D(n564), .Q(n26[10]));
    not g1720(n1658 ,n1657);
    not g1721(n2452 ,n2451);
    nor g1722(n1384 ,n1336 ,n1361);
    nor g1723(n789 ,n200 ,n665);
    not g1724(n2803 ,n2802);
    nor g1725(n2994 ,n2976 ,n2993);
    nor g1726(n1484 ,n1455 ,n1468);
    nor g1727(n2825 ,n2760 ,n2807);
    nor g1728(n2670 ,n2551 ,n2593);
    xnor g1729(n2823 ,n2732 ,n2765);
    nor g1730(n2781 ,n2716 ,n2743);
    nor g1731(n443 ,n222 ,n105);
    buf g1732(n12[0], 1'b0);
    not g1733(n1249 ,n1248);
    or g1734(n3159 ,n3154 ,n3133);
    nor g1735(n502 ,n152 ,n346);
    not g1736(n90 ,n89);
    nor g1737(n2624 ,n2520 ,n2563);
    not g1738(n1629 ,n1628);
    not g1739(n217 ,n22[4]);
    not g1740(n1147 ,n1146);
    or g1741(n3226 ,n3194 ,n3209);
    or g1742(n3249 ,n3192 ,n3242);
    xnor g1743(n1757 ,n1719 ,n1665);
    nor g1744(n517 ,n174 ,n348);
    buf g1745(n12[30], 1'b0);
    nor g1746(n786 ,n213 ,n666);
    xnor g1747(n1201 ,n1029 ,n1135);
    xnor g1748(n3296 ,n1457 ,n1494);
    nor g1749(n3190 ,n3118 ,n3142);
    not g1750(n124 ,n24[0]);
    not g1751(n237 ,n26[13]);
    not g1752(n1867 ,n20[7]);
    or g1753(n591 ,n403 ,n500);
    xnor g1754(n2688 ,n2628 ,n2579);
    nor g1755(n3197 ,n3096 ,n3142);
    nor g1756(n2635 ,n2528 ,n2573);
    nor g1757(n436 ,n318 ,n347);
    xnor g1758(n1345 ,n1318 ,n1264);
    xnor g1759(n32[4] ,n1821 ,n1816);
    not g1760(n2959 ,n22[2]);
    xnor g1761(n3291 ,n1346 ,n1329);
    nor g1762(n1574 ,n1522 ,n1532);
    nor g1763(n676 ,n107 ,n659);
    xnor g1764(n2238 ,n2051 ,n1961);
    not g1765(n3079 ,n3296);
    nor g1766(n780 ,n125 ,n666);
    not g1767(n1815 ,n1814);
    not g1768(n282 ,n10[6]);
    nor g1769(n2860 ,n2811 ,n2826);
    nor g1770(n2901 ,n2867 ,n2898);
    not g1771(n2040 ,n2039);
    not g1772(n952 ,n20[6]);
    not g1773(n2419 ,n2418);
    nor g1774(n689 ,n110 ,n648);
    or g1775(n880 ,n758 ,n709);
    nor g1776(n2057 ,n1864 ,n1874);
    nor g1777(n503 ,n143 ,n346);
    xnor g1778(n1177 ,n1016 ,n1092);
    not g1779(n59 ,n30[5]);
    nor g1780(n3136 ,n3314 ,n32[11]);
    nor g1781(n1603 ,n1519 ,n1558);
    buf g1782(n11[6], 1'b0);
    not g1783(n2107 ,n2106);
    nor g1784(n2450 ,n2327 ,n2325);
    dff g1785(.RN(n1), .SN(1'b1), .CK(n0), .D(n589), .Q(n10[13]));
    nor g1786(n1848 ,n1832 ,n1840);
    nor g1787(n1764 ,n1684 ,n1743);
    nor g1788(n101 ,n78 ,n99);
    nor g1789(n420 ,n263 ,n347);
    nor g1790(n1482 ,n1446 ,n1462);
    nor g1791(n3184 ,n3098 ,n3154);
    nor g1792(n1052 ,n957 ,n1038);
    not g1793(n308 ,n307);
    xnor g1794(n1290 ,n1028 ,n1243);
    nor g1795(n1774 ,n1698 ,n1755);
    nor g1796(n3178 ,n3091 ,n3142);
    or g1797(n533 ,n369 ,n447);
    nor g1798(n462 ,n138 ,n102);
    dff g1799(.RN(n1), .SN(1'b1), .CK(n0), .D(n553), .Q(n28[2]));
    nor g1800(n2281 ,n2031 ,n2222);
    not g1801(n115 ,n5[2]);
    dff g1802(.RN(n1), .SN(1'b1), .CK(n0), .D(n545), .Q(n28[12]));
    not g1803(n1888 ,n23[2]);
    not g1804(n221 ,n23[1]);
    nor g1805(n447 ,n246 ,n104);
    xnor g1806(n2408 ,n2243 ,n1993);
    xnor g1807(n2882 ,n2800 ,n2854);
    not g1808(n2818 ,n2817);
    nor g1809(n3243 ,n3143 ,n3162);
    nor g1810(n382 ,n248 ,n103);
    or g1811(n565 ,n383 ,n460);
    not g1812(n1908 ,n1907);
    or g1813(n3164 ,n3154 ,n3137);
    not g1814(n2889 ,n2888);
    nor g1815(n1899 ,n1887 ,n1872);
    or g1816(n906 ,n867 ,n866);
    buf g1817(n13[22], 1'b0);
    nor g1818(n2379 ,n2211 ,n2285);
    nor g1819(n2615 ,n2526 ,n2578);
    nor g1820(n1959 ,n1869 ,n1868);
    xor g1821(n3287 ,n2840 ,n2955);
    or g1822(n2132 ,n1879 ,n1888);
    not g1823(n1199 ,n1198);
    nor g1824(n2049 ,n1890 ,n1888);
    not g1825(n150 ,n24[5]);
    nor g1826(n1605 ,n1519 ,n1557);
    not g1827(n3098 ,n3261);
    not g1828(n119 ,n22[2]);
    not g1829(n2605 ,n2604);
    nor g1830(n3060 ,n3021 ,n3059);
    nor g1831(n1194 ,n1030 ,n1151);
    buf g1832(n11[14], 1'b0);
    nor g1833(n1271 ,n1219 ,n1204);
    or g1834(n822 ,n721 ,n682);
    nor g1835(n2619 ,n2557 ,n2569);
    nor g1836(n1834 ,n1794 ,n1809);
    nor g1837(n754 ,n224 ,n658);
    not g1838(n116 ,n19[4]);
    buf g1839(n11[24], n10[8]);
    not g1840(n1514 ,n3266);
    not g1841(n288 ,n15);
    nor g1842(n2045 ,n1892 ,n1891);
    xnor g1843(n985 ,n951 ,n20[2]);
    buf g1844(n12[18], n10[10]);
    not g1845(n1637 ,n1636);
    nor g1846(n377 ,n226 ,n105);
    buf g1847(n10[29], 1'b0);
    not g1848(n661 ,n662);
    nor g1849(n1282 ,n1198 ,n1229);
    or g1850(n640 ,n385 ,n638);
    nor g1851(n1855 ,n1842 ,n1854);
    xnor g1852(n32[8] ,n1846 ,n1853);
    not g1853(n2070 ,n2069);
    nor g1854(n796 ,n188 ,n652);
    nor g1855(n734 ,n120 ,n649);
    nor g1856(n506 ,n144 ,n346);
    xor g1857(n3274 ,n2637 ,n2584);
    xnor g1858(n3025 ,n3295 ,n3279);
    not g1859(n2651 ,n2650);
    xnor g1860(n2553 ,n2383 ,n2350);
    or g1861(n912 ,n896 ,n905);
    xnor g1862(n2922 ,n2892 ,n2869);
    nor g1863(n3135 ,n3313 ,n32[12]);
    xnor g1864(n1226 ,n1028 ,n1141);
    nor g1865(n3038 ,n3022 ,n3030);
    nor g1866(n1941 ,n1883 ,n1881);
    nor g1867(n1665 ,n1560 ,n1604);
    not g1868(n265 ,n26[8]);
    nor g1869(n2810 ,n2732 ,n2766);
    nor g1870(n1843 ,n1813 ,n1826);
    dff g1871(.RN(n1), .SN(1'b1), .CK(n0), .D(n913), .Q(n9[7]));
    nor g1872(n2212 ,n1942 ,n1902);
    nor g1873(n934 ,n70 ,n71);
    nor g1874(n1005 ,n975 ,n990);
    nor g1875(n2181 ,n1974 ,n2111);
    nor g1876(n1481 ,n1471 ,n1460);
    nor g1877(n714 ,n113 ,n663);
    nor g1878(n2807 ,n2702 ,n2771);
    or g1879(n837 ,n775 ,n781);
    nor g1880(n2749 ,n2614 ,n2713);
    xnor g1881(n1421 ,n1375 ,n1360);
    xnor g1882(n2975 ,n22[7] ,n23[7]);
    xnor g1883(n2976 ,n22[6] ,n23[6]);
    dff g1884(.RN(n1), .SN(1'b1), .CK(n0), .D(n598), .Q(n10[5]));
    xnor g1885(n1021 ,n1011 ,n995);
    nor g1886(n1146 ,n1079 ,n1121);
    not g1887(n3096 ,n3276);
    nor g1888(n1543 ,n1522 ,n1536);
    nor g1889(n671 ,n106 ,n648);
    not g1890(n1952 ,n1951);
    nor g1891(n675 ,n106 ,n659);
    not g1892(n2999 ,n3286);
    nor g1893(n1689 ,n1550 ,n1653);
    not g1894(n2770 ,n2769);
    xnor g1895(n1474 ,n1448 ,n1441);
    nor g1896(n2218 ,n2129 ,n1980);
    or g1897(n911 ,n902 ,n901);
    buf g1898(n9[10], 1'b0);
    or g1899(n559 ,n375 ,n467);
    nor g1900(n744 ,n185 ,n660);
    not g1901(n1355 ,n1354);
    xnor g1902(n3319 ,n3026 ,n3043);
    not g1903(n2328 ,n2327);
    not g1904(n2076 ,n2075);
    nor g1905(n2792 ,n2698 ,n2778);
    buf g1906(n12[1], 1'b0);
    nor g1907(n783 ,n205 ,n665);
    nor g1908(n1123 ,n958 ,n1089);
    xnor g1909(n1674 ,n1597 ,n1575);
    not g1910(n182 ,n19[3]);
    nor g1911(n2751 ,n2673 ,n2699);
    nor g1912(n3048 ,n3033 ,n3047);
    nor g1913(n92 ,n81 ,n90);
    not g1914(n253 ,n30[4]);
    or g1915(n3246 ,n3206 ,n3236);
    not g1916(n2346 ,n2345);
    not g1917(n173 ,n932);
    nor g1918(n2908 ,n2877 ,n2895);
    xnor g1919(n1373 ,n1017 ,n1344);
    not g1920(n129 ,n20[0]);
    or g1921(n570 ,n340 ,n360);
    not g1922(n1224 ,n1223);
    xnor g1923(n1710 ,n1583 ,n1634);
    nor g1924(n1762 ,n1731 ,n1733);
    nor g1925(n2302 ,n2005 ,n2163);
    buf g1926(n11[25], n10[9]);
    buf g1927(n11[28], n10[12]);
    nor g1928(n2314 ,n2014 ,n2172);
    nor g1929(n2347 ,n2179 ,n2296);
    not g1930(n2899 ,n2898);
    nor g1931(n1117 ,n956 ,n1064);
    nor g1932(n2708 ,n2636 ,n2643);
    not g1933(n919 ,n923);
    nor g1934(n2685 ,n2521 ,n2620);
    xnor g1935(n3289 ,n1185 ,n1065);
    buf g1936(n9[20], 1'b0);
    nor g1937(n1120 ,n947 ,n1062);
    nor g1938(n1153 ,n1046 ,n1112);
    not g1939(n3077 ,n3318);
    xnor g1940(n2790 ,n2727 ,n2661);
    not g1941(n3105 ,n3323);
    not g1942(n3097 ,n3301);
    nor g1943(n1571 ,n1521 ,n1532);
    xnor g1944(n2661 ,n2539 ,n2558);
    nor g1945(n3013 ,n3292 ,n3276);
    nor g1946(n2746 ,n2648 ,n2704);
    nor g1947(n2304 ,n2011 ,n2174);
    nor g1948(n1812 ,n1775 ,n1792);
    nor g1949(n3235 ,n3149 ,n3166);
    nor g1950(n1579 ,n1520 ,n1531);
    nor g1951(n2677 ,n2391 ,n2603);
    nor g1952(n3010 ,n3298 ,n3282);
    nor g1953(n2878 ,n2793 ,n2850);
    not g1954(n1904 ,n1903);
    dff g1955(.RN(n1), .SN(1'b1), .CK(n0), .D(n819), .Q(n22[7]));
    not g1956(n1809 ,n1808);
    not g1957(n160 ,n9[7]);
    nor g1958(n2481 ,n2186 ,n2437);
    not g1959(n1182 ,n1181);
    nor g1960(n494 ,n157 ,n104);
    nor g1961(n2575 ,n2427 ,n2496);
    not g1962(n2912 ,n2911);
    not g1963(n2960 ,n22[0]);
    nor g1964(n1728 ,n1651 ,n1677);
    not g1965(n2495 ,n2494);
    xnor g1966(n2785 ,n2734 ,n2742);
    nor g1967(n468 ,n134 ,n104);
    not g1968(n2227 ,n2226);
    not g1969(n104 ,n105);
    nor g1970(n1671 ,n1561 ,n1613);
    nor g1971(n2157 ,n2069 ,n2071);
    buf g1972(n13[23], 1'b0);
    nor g1973(n1588 ,n1522 ,n1556);
    xnor g1974(n331 ,n202 ,n116);
    nor g1975(n2434 ,n2335 ,n2331);
    not g1976(n2595 ,n2594);
    nor g1977(n988 ,n951 ,n970);
    nor g1978(n449 ,n230 ,n102);
    not g1979(n1442 ,n1441);
    nor g1980(n448 ,n152 ,n104);
    not g1981(n1382 ,n1381);
    nor g1982(n482 ,n248 ,n102);
    nor g1983(n2717 ,n2605 ,n2654);
    nor g1984(n406 ,n268 ,n105);
    not g1985(n1804 ,n1803);
    not g1986(n246 ,n28[8]);
    nor g1987(n2928 ,n2866 ,n2910);
    nor g1988(n2955 ,n2861 ,n2954);
    or g1989(n338 ,n295 ,n300);
    or g1990(n835 ,n730 ,n689);
    nor g1991(n1148 ,n1070 ,n1124);
    not g1992(n1635 ,n1634);
    not g1993(n1639 ,n1638);
    dff g1994(.RN(n1), .SN(1'b1), .CK(n0), .D(n835), .Q(n21[4]));
    not g1995(n2607 ,n2606);
    nor g1996(n2528 ,n2425 ,n2423);
    not g1997(n1328 ,n1327);
    nor g1998(n2950 ,n2949 ,n2925);
    dff g1999(.RN(n1), .SN(1'b1), .CK(n0), .D(n606), .Q(n30[1]));
    nor g2000(n3137 ,n3319 ,n32[6]);
    not g2001(n2074 ,n2073);
    not g2002(n2140 ,n2139);
    nor g2003(n1090 ,n958 ,n1032);
    xnor g2004(n1354 ,n1290 ,n1146);
    nor g2005(n1483 ,n1436 ,n1463);
    nor g2006(n706 ,n181 ,n660);
    not g2007(n285 ,n26[1]);
    not g2008(n2407 ,n2406);
    nor g2009(n359 ,n104 ,n326);
    nor g2010(n2698 ,n2626 ,n2652);
    nor g2011(n2812 ,n2684 ,n2773);
    buf g2012(n10[26], 1'b0);
    nor g2013(n1905 ,n1886 ,n1877);
    xnor g2014(n982 ,n963 ,n21[5]);
    nor g2015(n1929 ,n1863 ,n1866);
    nor g2016(n388 ,n230 ,n103);
    nor g2017(n739 ,n218 ,n662);
    nor g2018(n2202 ,n2026 ,n2078);
    buf g2019(n13[26], n10[2]);
    nor g2020(n1001 ,n949 ,n992);
    xnor g2021(n2465 ,n2261 ,n1923);
    nor g2022(n756 ,n240 ,n658);
    nor g2023(n2001 ,n1884 ,n1870);
    nor g2024(n3144 ,n3108 ,n3074);
    xnor g2025(n1379 ,n1200 ,n1331);
    xnor g2026(n1558 ,n3268 ,n23[4]);
    nor g2027(n3022 ,n3004 ,n3001);
    not g2028(n2609 ,n2608);
    nor g2029(n2598 ,n2511 ,n2546);
    not g2030(n2231 ,n2230);
    nor g2031(n794 ,n219 ,n654);
    nor g2032(n340 ,n260 ,n319);
    nor g2033(n1840 ,n1820 ,n1829);
    nor g2034(n2874 ,n2790 ,n2842);
    nor g2035(n1267 ,n1174 ,n1206);
    nor g2036(n352 ,n104 ,n331);
    not g2037(n264 ,n26[2]);
    nor g2038(n3066 ,n3017 ,n3065);
    xnor g2039(n2841 ,n2787 ,n2767);
    nor g2040(n612 ,n348 ,n437);
    not g2041(n233 ,n26[9]);
    nor g2042(n2170 ,n1917 ,n1925);
    or g2043(n3231 ,n3208 ,n3179);
    or g2044(n3251 ,n3188 ,n3241);
    not g2045(n54 ,n30[6]);
    nor g2046(n2004 ,n1882 ,n1889);
    or g2047(n896 ,n790 ,n864);
    nor g2048(n662 ,n322 ,n646);
    not g2049(n2007 ,n2006);
    or g2050(n1530 ,n1509 ,n1525);
    nor g2051(n1897 ,n1883 ,n1877);
    xnor g2052(n2430 ,n2255 ,n1921);
    nor g2053(n3241 ,n3152 ,n3160);
    nor g2054(n3054 ,n3027 ,n3053);
    xnor g2055(n3034 ,n3299 ,n3283);
    or g2056(n601 ,n431 ,n510);
    nor g2057(n2200 ,n2048 ,n2090);
    nor g2058(n2442 ,n2270 ,n2366);
    nor g2059(n2354 ,n2194 ,n2297);
    nor g2060(n2023 ,n1883 ,n1861);
    or g2061(n1285 ,n1029 ,n1226);
    nor g2062(n1389 ,n1325 ,n1349);
    nor g2063(n1913 ,n1892 ,n1878);
    nor g2064(n3216 ,n3084 ,n3142);
    xnor g2065(n1356 ,n1289 ,n1215);
    not g2066(n1029 ,n1030);
    nor g2067(n451 ,n225 ,n104);
    not g2068(n1807 ,n1806);
    or g2069(n592 ,n421 ,n501);
    xnor g2070(n2650 ,n2545 ,n2424);
    or g2071(n546 ,n368 ,n448);
    not g2072(n1000 ,n21[0]);
    not g2073(n2088 ,n2087);
    not g2074(n2018 ,n2017);
    nor g2075(n453 ,n136 ,n104);
    nor g2076(n718 ,n107 ,n668);
    nor g2077(n2496 ,n2362 ,n2438);
    not g2078(n186 ,n19[2]);
    nor g2079(n2872 ,n2763 ,n2848);
    nor g2080(n816 ,n221 ,n654);
    xor g2081(n3271 ,n20[7] ,n21[7]);
    not g2082(n2754 ,n2753);
    nor g2083(n1124 ,n949 ,n1089);
    xnor g2084(n3306 ,n2980 ,n2983);
    nor g2085(n461 ,n144 ,n102);
    not g2086(n1528 ,n3268);
    or g2087(n829 ,n725 ,n669);
    nor g2088(n1059 ,n946 ,n1036);
    not g2089(n229 ,n25[5]);
    nor g2090(n1895 ,n1883 ,n1872);
    not g2091(n1598 ,n1597);
    nor g2092(n1559 ,n1520 ,n1536);
    nor g2093(n1065 ,n1016 ,n1039);
    not g2094(n2129 ,n2128);
    nor g2095(n432 ,n259 ,n347);
    nor g2096(n1489 ,n1484 ,n1478);
    not g2097(n202 ,n28[4]);
    nor g2098(n71 ,n56 ,n69);
    nor g2099(n1634 ,n1544 ,n1587);
    nor g2100(n422 ,n139 ,n347);
    nor g2101(n1775 ,n1737 ,n1753);
    nor g2102(n1731 ,n1678 ,n1720);
    nor g2103(n760 ,n124 ,n658);
    nor g2104(n2564 ,n2348 ,n2517);
    nor g2105(n2489 ,n2463 ,n2451);
    nor g2106(n2721 ,n2632 ,n2681);
    nor g2107(n2167 ,n1921 ,n1951);
    not g2108(n205 ,n20[7]);
    nor g2109(n52 ,n47 ,n51);
    not g2110(n1978 ,n1977);
    xnor g2111(n1184 ,n1016 ,n1093);
    nor g2112(n1144 ,n1052 ,n1120);
    or g2113(n855 ,n751 ,n675);
    nor g2114(n1949 ,n1884 ,n1866);
    nor g2115(n2318 ,n2086 ,n2216);
    or g2116(n588 ,n418 ,n498);
    xnor g2117(n1708 ,n1644 ,n1636);
    not g2118(n263 ,n10[13]);
    or g2119(n913 ,n910 ,n904);
    nor g2120(n1043 ,n958 ,n1036);
    not g2121(n1818 ,n1817);
    not g2122(n228 ,n10[7]);
    nor g2123(n2176 ,n1941 ,n1901);
    not g2124(n3099 ,n27[1]);
    not g2125(n1284 ,n1283);
    nor g2126(n67 ,n30[3] ,n65);
    nor g2127(n1454 ,n1414 ,n1423);
    nor g2128(n2329 ,n2208 ,n2286);
    nor g2129(n3196 ,n3083 ,n3154);
    nor g2130(n1917 ,n1880 ,n1873);
    nor g2131(n1784 ,n1736 ,n1750);
    not g2132(n1998 ,n1997);
    xnor g2133(n2277 ,n2012 ,n2106);
    nor g2134(n521 ,n292 ,n347);
    xnor g2135(n2692 ,n2588 ,n2533);
    nor g2136(n403 ,n276 ,n347);
    or g2137(n857 ,n750 ,n703);
    nor g2138(n2759 ,n2677 ,n2708);
    nor g2139(n2915 ,n2868 ,n2899);
    or g2140(n891 ,n766 ,n715);
    or g2141(n335 ,n5[1] ,n297);
    nor g2142(n2073 ,n1865 ,n1875);
    xnor g2143(n3293 ,n1397 ,n1437);
    xnor g2144(n2542 ,n2404 ,n2420);
    not g2145(n3072 ,n32[5]);
    nor g2146(n3191 ,n3082 ,n3141);
    not g2147(n1300 ,n1299);
    dff g2148(.RN(n1), .SN(1'b1), .CK(n0), .D(n916), .Q(n9[2]));
    dff g2149(.RN(n1), .SN(1'b1), .CK(n0), .D(n579), .Q(n29[7]));
    nor g2150(n3205 ,n3071 ,n3155);
    nor g2151(n512 ,n162 ,n346);
    or g2152(n584 ,n413 ,n518);
    not g2153(n2111 ,n2110);
    or g2154(n3222 ,n3175 ,n3169);
    xnor g2155(n1030 ,n1007 ,n995);
    nor g2156(n2449 ,n2336 ,n2332);
    nor g2157(n1798 ,n1767 ,n1784);
    not g2158(n1940 ,n1939);
    buf g2159(n9[11], 1'b0);
    nor g2160(n2618 ,n2581 ,n2504);
    nor g2161(n1704 ,n1624 ,n1647);
    nor g2162(n702 ,n113 ,n659);
    not g2163(n3004 ,n3288);
    or g2164(n562 ,n496 ,n471);
    xnor g2165(n2387 ,n2271 ,n1953);
    nor g2166(n667 ,n525 ,n645);
    or g2167(n885 ,n762 ,n711);
    not g2168(n1881 ,n22[4]);
    xnor g2169(n2798 ,n2725 ,n2700);
    xnor g2170(n1289 ,n1242 ,n1222);
    nor g2171(n1280 ,n1195 ,n1227);
    not g2172(n1936 ,n1935);
    or g2173(n832 ,n728 ,n687);
    or g2174(n828 ,n777 ,n776);
    not g2175(n96 ,n95);
    xnor g2176(n1438 ,n1404 ,n1297);
    nor g2177(n818 ,n256 ,n653);
    nor g2178(n705 ,n114 ,n657);
    nor g2179(n716 ,n111 ,n650);
    not g2180(n523 ,n524);
    nor g2181(n2836 ,n2734 ,n2795);
    xor g2182(n32[3] ,n1788 ,n1778);
    nor g2183(n703 ,n109 ,n659);
    nor g2184(n427 ,n241 ,n347);
    nor g2185(n2104 ,n1892 ,n1889);
    nor g2186(n2438 ,n2350 ,n2361);
    nor g2187(n2934 ,n2912 ,n2920);
    nor g2188(n1099 ,n1015 ,n1071);
    nor g2189(n2206 ,n2082 ,n2088);
    xnor g2190(n2540 ,n2461 ,n2457);
    nor g2191(n2620 ,n2514 ,n2559);
    nor g2192(n400 ,n269 ,n105);
    dff g2193(.RN(n1), .SN(1'b1), .CK(n0), .D(n882), .Q(n24[0]));
    nor g2194(n1961 ,n1865 ,n1874);
    nor g2195(n2211 ,n1898 ,n1950);
    nor g2196(n1721 ,n1667 ,n1688);
    or g2197(n902 ,n827 ,n824);
    not g2198(n2030 ,n2029);
    dff g2199(.RN(n1), .SN(1'b1), .CK(n0), .D(n602), .Q(n10[1]));
    nor g2200(n2574 ,n2426 ,n2497);
    not g2201(n72 ,n71);
    nor g2202(n2864 ,n2802 ,n2856);
    nor g2203(n1779 ,n1725 ,n1752);
    nor g2204(n682 ,n112 ,n650);
    nor g2205(n776 ,n196 ,n655);
    xor g2206(n3309 ,n2979 ,n2990);
    xor g2207(n944 ,n1196 ,n1184);
    nor g2208(n2027 ,n1869 ,n1889);
    not g2209(n3081 ,n3257);
    nor g2210(n1786 ,n1689 ,n1760);
    nor g2211(n2226 ,n2125 ,n2131);
    nor g2212(n1907 ,n1883 ,n1873);
    nor g2213(n1696 ,n1664 ,n1631);
    not g2214(n176 ,n937);
    xnor g2215(n1553 ,n3264 ,n23[0]);
    nor g2216(n2286 ,n2100 ,n2142);
    nor g2217(n1257 ,n1182 ,n942);
    or g2218(n897 ,n796 ,n868);
    not g2219(n241 ,n10[5]);
    or g2220(n3227 ,n3185 ,n3210);
    nor g2221(n1852 ,n1843 ,n1851);
    not g2222(n1351 ,n1350);
    nor g2223(n758 ,n190 ,n658);
    not g2224(n1550 ,n1549);
    xnor g2225(n3036 ,n3302 ,n3286);
    nor g2226(n1577 ,n1520 ,n1530);
    xnor g2227(n2845 ,n2785 ,n2794);
    nor g2228(n2171 ,n1971 ,n1957);
    or g2229(n824 ,n771 ,n770);
    xor g2230(n942 ,n1030 ,n1151);
    nor g2231(n457 ,n262 ,n104);
    nor g2232(n2509 ,n2339 ,n2407);
    nor g2233(n3015 ,n3294 ,n3278);
    nor g2234(n2311 ,n2003 ,n2168);
    not g2235(n2225 ,n2224);
    xnor g2236(n2600 ,n2479 ,n2418);
    nor g2237(n1816 ,n1781 ,n1797);
    nor g2238(n2671 ,n2598 ,n2601);
    nor g2239(n2041 ,n1863 ,n1891);
    not g2240(n2844 ,n2843);
    dff g2241(.RN(n1), .SN(1'b1), .CK(n0), .D(n918), .Q(n9[4]));
    or g2242(n2014 ,n1882 ,n1888);
    xnor g2243(n3282 ,n2939 ,n2945);
    nor g2244(n1254 ,n1233 ,n1207);
    nor g2245(n2333 ,n2206 ,n2288);
    nor g2246(n2570 ,n2416 ,n2503);
    or g2247(n878 ,n805 ,n806);
    not g2248(n1932 ,n1931);
    not g2249(n219 ,n23[5]);
    dff g2250(.RN(n1), .SN(1'b1), .CK(n0), .D(n854), .Q(n19[4]));
    not g2251(n3073 ,n32[2]);
    xnor g2252(n3031 ,n3298 ,n3282);
    not g2253(n1206 ,n1205);
    nor g2254(n2706 ,n2575 ,n2682);
    not g2255(n238 ,n25[3]);
    nor g2256(n3239 ,n3150 ,n3159);
    nor g2257(n516 ,n175 ,n348);
    xor g2258(n2536 ,n2470 ,n2394);
    xnor g2259(n2767 ,n2688 ,n2632);
    nor g2260(n1566 ,n1519 ,n1534);
    not g2261(n1982 ,n1981);
    nor g2262(n1107 ,n957 ,n1064);
    not g2263(n168 ,n930);
    not g2264(n1171 ,n1170);
    nor g2265(n492 ,n153 ,n102);
    nor g2266(n1395 ,n1334 ,n1364);
    nor g2267(n1334 ,n1017 ,n1316);
    not g2268(n2026 ,n2025);
    not g2269(n2505 ,n2504);
    not g2270(n197 ,n23[6]);
    nor g2271(n2744 ,n2625 ,n2701);
    nor g2272(n1589 ,n1521 ,n1551);
    not g2273(n2094 ,n2093);
    nor g2274(n3011 ,n3297 ,n3281);
    xnor g2275(n2794 ,n2728 ,n2660);
    nor g2276(n2695 ,n2468 ,n2644);
    not g2277(n3102 ,n32[9]);
    not g2278(n1666 ,n1665);
    or g2279(n31[6] ,n3220 ,n3246);
    not g2280(n3085 ,n3277);
    xnor g2281(n2544 ,n2463 ,n2451);
    buf g2282(n12[9], n10[1]);
    nor g2283(n1562 ,n1519 ,n1535);
    dff g2284(.RN(n1), .SN(1'b1), .CK(n0), .D(n823), .Q(n22[4]));
    nor g2285(n2865 ,n2832 ,n2859);
    or g2286(n3233 ,n3199 ,n3215);
    xnor g2287(n1039 ,n1017 ,n999);
    not g2288(n252 ,n9[6]);
    nor g2289(n390 ,n126 ,n105);
    nor g2290(n730 ,n203 ,n649);
    nor g2291(n1047 ,n948 ,n1036);
    not g2292(n2274 ,n2273);
    nor g2293(n1042 ,n958 ,n1034);
    not g2294(n2038 ,n2037);
    or g2295(n39 ,n30[7] ,n38);
    xnor g2296(n1402 ,n1286 ,n1371);
    nor g2297(n2991 ,n2979 ,n2990);
    not g2298(n1464 ,n1463);
    nor g2299(n2777 ,n2758 ,n2746);
    nor g2300(n2051 ,n1885 ,n1878);
    or g2301(n666 ,n324 ,n643);
    or g2302(n626 ,n314 ,n609);
    not g2303(n2223 ,n2222);
    nor g2304(n430 ,n161 ,n347);
    nor g2305(n3051 ,n3007 ,n3050);
    xnor g2306(n2478 ,n1931 ,n2345);
    nor g2307(n2308 ,n2117 ,n2143);
    buf g2308(n13[14], 1'b0);
    nor g2309(n2047 ,n1886 ,n1873);
    nor g2310(n1997 ,n1863 ,n1888);
    xnor g2311(n2390 ,n2252 ,n2120);
    nor g2312(n2142 ,n1961 ,n2051);
    not g2313(n1984 ,n1983);
    buf g2314(n9[19], 1'b0);
    nor g2315(n2527 ,n2411 ,n2401);
    not g2316(n2703 ,n2702);
    not g2317(n1339 ,n1338);
    dff g2318(.RN(n1), .SN(1'b1), .CK(n0), .D(n836), .Q(n21[3]));
    not g2319(n1987 ,n1986);
    nor g2320(n487 ,n151 ,n102);
    nor g2321(n761 ,n193 ,n664);
    nor g2322(n2357 ,n2229 ,n2275);
    or g2323(n560 ,n400 ,n451);
    nor g2324(n2168 ,n2073 ,n1903);
    not g2325(n222 ,n29[10]);
    nor g2326(n2197 ,n1916 ,n2050);
    nor g2327(n2617 ,n2506 ,n2570);
    not g2328(n1460 ,n1459);
    buf g2329(n9[17], 1'b0);
    not g2330(n155 ,n30[1]);
    nor g2331(n1014 ,n960 ,n992);
    nor g2332(n1053 ,n956 ,n1036);
    or g2333(n3220 ,n3173 ,n3171);
    nor g2334(n1112 ,n958 ,n1063);
    nor g2335(n2730 ,n2671 ,n2710);
    not g2336(n2066 ,n2065);
    or g2337(n309 ,n5[11] ,n5[10]);
    nor g2338(n1595 ,n1521 ,n1553);
    dff g2339(.RN(n1), .SN(1'b1), .CK(n0), .D(n840), .Q(n21[0]));
    nor g2340(n2361 ,n2224 ,n2268);
    not g2341(n1521 ,n24[2]);
    nor g2342(n3171 ,n3119 ,n3141);
    buf g2343(n12[11], n10[3]);
    nor g2344(n1979 ,n1867 ,n1876);
    nor g2345(n2162 ,n2079 ,n2055);
    nor g2346(n51 ,n49 ,n48);
    nor g2347(n1616 ,n1522 ,n1551);
    nor g2348(n3202 ,n3116 ,n3141);
    xor g2349(n2263 ,n2117 ,n1909);
    nor g2350(n2065 ,n1865 ,n1877);
    dff g2351(.RN(n1), .SN(1'b1), .CK(n0), .D(n822), .Q(n22[5]));
    nor g2352(n2375 ,n2212 ,n2289);
    xnor g2353(n2641 ,n2494 ,n2583);
    or g2354(n598 ,n427 ,n507);
    not g2355(n1027 ,n1028);
    nor g2356(n2112 ,n1871 ,n1861);
    or g2357(n882 ,n760 ,n678);
    buf g2358(n10[30], 1'b0);
    nor g2359(n2307 ,n2114 ,n2164);
    dff g2360(.RN(n1), .SN(1'b1), .CK(n0), .D(n856), .Q(n19[3]));
    not g2361(n1886 ,n20[3]);
    nor g2362(n1108 ,n947 ,n1064);
    or g2363(n908 ,n878 ,n875);
    nor g2364(n2969 ,n22[0] ,n23[0]);
    nor g2365(n2149 ,n2023 ,n1965);
    not g2366(n1317 ,n1316);
    nor g2367(n1480 ,n1435 ,n1464);
    nor g2368(n1056 ,n947 ,n1034);
    nor g2369(n1269 ,n1199 ,n1228);
    not g2370(n2334 ,n2333);
    nor g2371(n89 ,n84 ,n87);
    or g2372(n575 ,n390 ,n461);
    nor g2373(n438 ,n223 ,n347);
    xnor g2374(n1031 ,n969 ,n1019);
    nor g2375(n3151 ,n3075 ,n3103);
    xnor g2376(n1325 ,n1251 ,n1225);
    nor g2377(n3020 ,n3000 ,n3006);
    dff g2378(.RN(n1), .SN(1'b1), .CK(n0), .D(n880), .Q(n24[2]));
    not g2379(n2733 ,n2732);
    not g2380(n1738 ,n1737);
    nor g2381(n3132 ,n3323 ,n32[2]);
    dff g2382(.RN(n1), .SN(1'b1), .CK(n0), .D(n539), .Q(n26[13]));
    nor g2383(n1140 ,n1084 ,n1126);
    not g2384(n2034 ,n2033);
    nor g2385(n473 ,n920 ,n102);
    not g2386(n2466 ,n2465);
    not g2387(n1216 ,n1215);
    nor g2388(n2512 ,n2367 ,n2397);
    not g2389(n3106 ,n3322);
    not g2390(n284 ,n29[7]);
    nor g2391(n2974 ,n2958 ,n2962);
    xnor g2392(n1397 ,n1368 ,n1338);
    or g2393(n585 ,n414 ,n519);
    xnor g2394(n3273 ,n2217 ,n2537);
    buf g2395(n13[5], 1'b0);
    nor g2396(n488 ,n176 ,n102);
    xnor g2397(n1240 ,n1026 ,n1144);
    xnor g2398(n2558 ,n2385 ,n2351);
    nor g2399(n1491 ,n1485 ,n1479);
    nor g2400(n3167 ,n3085 ,n3142);
    xnor g2401(n1755 ,n1710 ,n1667);
    or g2402(n339 ,n298 ,n312);
    xnor g2403(n2640 ,n2504 ,n2581);
    nor g2404(n1697 ,n1584 ,n1634);
    xnor g2405(n2612 ,n2476 ,n2353);
    or g2406(n304 ,n5[23] ,n5[22]);
    nor g2407(n2312 ,n2134 ,n2141);
    nor g2408(n2351 ,n2184 ,n2291);
    nor g2409(n1451 ,n1395 ,n1433);
    nor g2410(n1196 ,n1028 ,n1152);
    nor g2411(n413 ,n238 ,n349);
    nor g2412(n2061 ,n1892 ,n1862);
    not g2413(n2366 ,n2365);
    nor g2414(n2707 ,n2627 ,n2653);
    nor g2415(n1601 ,n1519 ,n1552);
    nor g2416(n2630 ,n2519 ,n2576);
    dff g2417(.RN(n1), .SN(1'b1), .CK(n0), .D(n572), .Q(n26[4]));
    not g2418(n1229 ,n1228);
    not g2419(n1976 ,n1975);
    or g2420(n525 ,n146 ,n337);
    not g2421(n224 ,n24[6]);
    nor g2422(n2230 ,n1990 ,n1987);
    xnor g2423(n1805 ,n1786 ,n1581);
    nor g2424(n3052 ,n3024 ,n3051);
    xnor g2425(n2418 ,n2250 ,n2112);
    buf g2426(n13[4], 1'b0);
    nor g2427(n1915 ,n1887 ,n1881);
    nor g2428(n1002 ,n946 ,n992);
    or g2429(n3250 ,n3183 ,n3239);
    nor g2430(n1581 ,n1520 ,n1535);
    nor g2431(n619 ,n257 ,n524);
    nor g2432(n1283 ,n1183 ,n1241);
    not g2433(n2737 ,n2736);
    or g2434(n365 ,n313 ,n341);
    or g2435(n31[0] ,n3231 ,n3248);
    nor g2436(n1995 ,n1882 ,n1868);
    nor g2437(n1493 ,n1449 ,n1490);
    nor g2438(n2222 ,n2000 ,n2127);
    nor g2439(n768 ,n199 ,n664);
    nor g2440(n1075 ,n949 ,n1040);
    nor g2441(n1933 ,n1863 ,n1868);
    xnor g2442(n329 ,n121 ,n180);
    not g2443(n1281 ,n1280);
    nor g2444(n1841 ,n1818 ,n1827);
    xnor g2445(n2237 ,n2063 ,n1907);
    nor g2446(n777 ,n120 ,n666);
    or g2447(n3166 ,n3154 ,n3135);
    not g2448(n437 ,n436);
    or g2449(n31[11] ,n3227 ,n3223);
    nor g2450(n1413 ,n1365 ,n1386);
    not g2451(n204 ,n28[3]);
    nor g2452(n2937 ,n2909 ,n2923);
    buf g2453(n10[31], 1'b0);
    not g2454(n1034 ,n1033);
    xnor g2455(n1712 ,n1630 ,n1663);
    not g2456(n2705 ,n2704);
    nor g2457(n1313 ,n1249 ,n1275);
    not g2458(n2221 ,n2220);
    xnor g2459(n2787 ,n2751 ,n2706);
    dff g2460(.RN(n1), .SN(1'b1), .CK(n0), .D(n857), .Q(n19[2]));
    nor g2461(n2713 ,n2607 ,n2650);
    nor g2462(n1378 ,n1352 ,n1350);
    nor g2463(n1761 ,n1703 ,n1741);
    not g2464(n1752 ,n1751);
    nor g2465(n1338 ,n1267 ,n1310);
    nor g2466(n2664 ,n2494 ,n2630);
    xnor g2467(n1219 ,n1029 ,n1143);
    not g2468(n2044 ,n2043);
    dff g2469(.RN(n1), .SN(1'b1), .CK(n0), .D(n567), .Q(n28[1]));
    xnor g2470(n3298 ,n1486 ,n1498);
    nor g2471(n100 ,n25[6] ,n98);
    xnor g2472(n1183 ,n1027 ,n1113);
    or g2473(n547 ,n388 ,n458);
    not g2474(n1926 ,n1925);
    not g2475(n1930 ,n1929);
    or g2476(n918 ,n898 ,n907);
    nor g2477(n2966 ,n22[1] ,n23[1]);
    or g2478(n860 ,n782 ,n818);
    nor g2479(n1086 ,n960 ,n1038);
    not g2480(n1446 ,n1445);
    xnor g2481(n1458 ,n1398 ,n1429);
    not g2482(n166 ,n933);
    nor g2483(n1074 ,n949 ,n1032);
    or g2484(n826 ,n724 ,n685);
    not g2485(n2064 ,n2063);
    not g2486(n114 ,n6[6]);
    not g2487(n1754 ,n1753);
    nor g2488(n466 ,n255 ,n102);
    not g2489(n346 ,n347);
    xnor g2490(n3303 ,n1458 ,n1508);
    not g2491(n198 ,n28[7]);
    nor g2492(n3204 ,n3072 ,n3155);
    xnor g2493(n3276 ,n2824 ,n2784);
    not g2494(n953 ,n21[7]);
    or g2495(n342 ,n316 ,n317);
    xnor g2496(n2472 ,n2367 ,n2375);
    nor g2497(n637 ,n305 ,n635);
    or g2498(n887 ,n763 ,n712);
    nor g2499(n2566 ,n2347 ,n2513);
    not g2500(n1517 ,n23[7]);
    xnor g2501(n1473 ,n1444 ,n1427);
    nor g2502(n1549 ,n1520 ,n1538);
    not g2503(n2556 ,n2555);
    nor g2504(n1082 ,n959 ,n1036);
    nor g2505(n1999 ,n1886 ,n1876);
    not g2506(n994 ,n993);
    not g2507(n3101 ,n32[3]);
    nor g2508(n1561 ,n1519 ,n1536);
    nor g2509(n1730 ,n1693 ,n1728);
    nor g2510(n2436 ,n2177 ,n2381);
    nor g2511(n2126 ,n1871 ,n1875);
    xnor g2512(n3321 ,n3028 ,n3039);
    not g2513(n254 ,n10[11]);
    xnor g2514(n2652 ,n2543 ,n2469);
    xnor g2515(n2396 ,n2237 ,n2004);
    not g2516(n207 ,n22[6]);
    not g2517(n1032 ,n1031);
    not g2518(n1826 ,n1825);
    dff g2519(.RN(n1), .SN(1'b1), .CK(n0), .D(n585), .Q(n25[2]));
    nor g2520(n2146 ,n2029 ,n1913);
    buf g2521(n12[29], 1'b0);
    nor g2522(n1993 ,n1884 ,n1868);
    xnor g2523(n2494 ,n2322 ,n2352);
    nor g2524(n1155 ,n1061 ,n1111);
    or g2525(n3219 ,n3200 ,n3182);
    not g2526(n1813 ,n1812);
    dff g2527(.RN(n1), .SN(1'b1), .CK(n0), .D(n574), .Q(n26[2]));
    xnor g2528(n1737 ,n1674 ,n1668);
    xnor g2529(n1186 ,n1016 ,n1099);
    nor g2530(n1261 ,n1222 ,n1215);
    xnor g2531(n2648 ,n2542 ,n2430);
    xnor g2532(n327 ,n204 ,n182);
    or g2533(n836 ,n731 ,n690);
    xnor g2534(n1318 ,n1030 ,n1226);
    nor g2535(n1363 ,n1282 ,n1324);
    buf g2536(n11[2], 1'b0);
    nor g2537(n405 ,n280 ,n103);
    nor g2538(n2986 ,n2973 ,n2985);
    not g2539(n2653 ,n2652);
    nor g2540(n2440 ,n2284 ,n2352);
    dff g2541(.RN(n1), .SN(1'b1), .CK(n0), .D(n605), .Q(n29[3]));
    not g2542(n2276 ,n2275);
    buf g2543(n12[15], n10[7]);
    buf g2544(n13[9], 1'b0);
    not g2545(n958 ,n3304);
    not g2546(n2046 ,n2045);
    not g2547(n2857 ,n2856);
    not g2548(n3086 ,n3274);
    nor g2549(n2205 ,n2092 ,n1910);
    nor g2550(n680 ,n107 ,n663);
    not g2551(n3121 ,n3260);
    not g2552(n2997 ,n3302);
    or g2553(n3165 ,n3154 ,n3139);
    xnor g2554(n2883 ,n2802 ,n2856);
    not g2555(n1584 ,n1583);
    not g2556(n3108 ,n3317);
    nor g2557(n1839 ,n1814 ,n1823);
    nor g2558(n2446 ,n1932 ,n2345);
    nor g2559(n1975 ,n1882 ,n1862);
    not g2560(n111 ,n6[7]);
    nor g2561(n2373 ,n2209 ,n2311);
    not g2562(n3089 ,n3263);
    nor g2563(n2859 ,n2815 ,n2825);
    nor g2564(n2043 ,n1867 ,n1861);
    not g2565(n1218 ,n1217);
    nor g2566(n3174 ,n3123 ,n3142);
    nor g2567(n2696 ,n2685 ,n2656);
    or g2568(n553 ,n394 ,n463);
    not g2569(n3070 ,n32[4]);
    nor g2570(n3043 ,n3008 ,n3042);
    nor g2571(n1626 ,n1579 ,n1599);
    or g2572(n296 ,n26[10] ,n26[11]);
    not g2573(n2499 ,n2498);
    nor g2574(n3039 ,n3009 ,n3038);
    not g2575(n2096 ,n2095);
    or g2576(n603 ,n433 ,n512);
    not g2577(n2011 ,n2010);
    or g2578(n1534 ,n1526 ,n1511);
    nor g2579(n1248 ,n1186 ,n1193);
    not g2580(n281 ,n30[7]);
    nor g2581(n446 ,n234 ,n105);
    or g2582(n907 ,n870 ,n869);
    buf g2583(n11[4], 1'b0);
    xnor g2584(n2426 ,n2248 ,n2230);
    nor g2585(n2925 ,n2887 ,n2907);
    dff g2586(.RN(n1), .SN(1'b1), .CK(n0), .D(n881), .Q(n24[1]));
    buf g2587(n9[14], 1'b0);
    nor g2588(n1012 ,n948 ,n992);
    nor g2589(n1165 ,n1081 ,n1101);
    nor g2590(n2029 ,n1871 ,n1881);
    nor g2591(n2521 ,n2369 ,n2415);
    nor g2592(n366 ,n236 ,n105);
    not g2593(n1880 ,n20[6]);
    nor g2594(n2299 ,n2116 ,n2175);
    buf g2595(n9[13], 1'b0);
    xnor g2596(n2658 ,n2540 ,n2467);
    nor g2597(n2523 ,n2342 ,n2465);
    not g2598(n951 ,n21[2]);
    not g2599(n1513 ,n3267);
    not g2600(n950 ,n20[1]);
    not g2601(n2105 ,n2104);
    or g2602(n642 ,n137 ,n639);
    buf g2603(n10[18], 1'b0);
    nor g2604(n798 ,n203 ,n666);
    dff g2605(.RN(n1), .SN(1'b1), .CK(n0), .D(n911), .Q(n9[1]));
    not g2606(n178 ,n926);
    buf g2607(n11[16], n10[0]);
    nor g2608(n439 ,n279 ,n103);
    buf g2609(n9[16], 1'b0);
    nor g2610(n781 ,n117 ,n656);
    not g2611(n2905 ,n2904);
    nor g2612(n1646 ,n1546 ,n1616);
    nor g2613(n2926 ,n2902 ,n2891);
    not g2614(n1416 ,n1415);
    nor g2615(n3059 ,n3034 ,n3058);
    xnor g2616(n1022 ,n1000 ,n997);
    nor g2617(n3211 ,n3074 ,n3155);
    buf g2618(n10[21], 1'b0);
    nor g2619(n765 ,n216 ,n664);
    xnor g2620(n2248 ,n1919 ,n1959);
    xnor g2621(n1729 ,n1686 ,n1704);
    not g2622(n2032 ,n2031);
    xnor g2623(n2822 ,n2769 ,n2753);
    nor g2624(n724 ,n119 ,n651);
    or g2625(n904 ,n860 ,n859);
    nor g2626(n1792 ,n1739 ,n1782);
    xnor g2627(n2404 ,n2253 ,n1975);
    nor g2628(n723 ,n211 ,n651);
    not g2629(n247 ,n30[5]);
    or g2630(n48 ,n25[1] ,n25[0]);
    or g2631(n31[3] ,n3224 ,n3249);
    nor g2632(n3140 ,n3320 ,n32[5]);
    nor g2633(n3323 ,n3022 ,n3014);
    not g2634(n3067 ,n27[0]);
    xnor g2635(n1417 ,n1383 ,n1301);
    not g2636(n1520 ,n24[3]);
    nor g2637(n1844 ,n1815 ,n1824);
    or g2638(n627 ,n311 ,n613);
    dff g2639(.RN(n1), .SN(1'b1), .CK(n0), .D(n541), .Q(n29[1]));
    not g2640(n179 ,n931);
    nor g2641(n409 ,n285 ,n105);
    nor g2642(n2091 ,n1886 ,n1861);
    nor g2643(n1659 ,n1545 ,n1591);
    nor g2644(n1434 ,n1340 ,n1403);
    nor g2645(n742 ,n129 ,n662);
    not g2646(n130 ,n20[5]);
    or g2647(n298 ,n5[17] ,n5[16]);
    nor g2648(n2519 ,n2371 ,n2403);
    not g2649(n2497 ,n2496);
    xnor g2650(n2980 ,n22[2] ,n23[2]);
    nor g2651(n2485 ,n2424 ,n2422);
    nor g2652(n2753 ,n2678 ,n2711);
    not g2653(n3117 ,n3292);
    xnor g2654(n1418 ,n1385 ,n1303);
    nor g2655(n354 ,n104 ,n332);
    nor g2656(n500 ,n163 ,n346);
    nor g2657(n688 ,n112 ,n648);
    nor g2658(n1611 ,n1522 ,n1557);
    nor g2659(n2195 ,n1900 ,n2022);
    xnor g2660(n1554 ,n3271 ,n23[7]);
    nor g2661(n2115 ,n1884 ,n1889);
    not g2662(n960 ,n3312);
    nor g2663(n1849 ,n1833 ,n1848);
    not g2664(n250 ,n25[7]);
    buf g2665(n11[31], n10[15]);
    nor g2666(n3021 ,n3003 ,n3002);
    dff g2667(.RN(n1), .SN(1'b1), .CK(n0), .D(n568), .Q(n26[7]));
    not g2668(n1882 ,n21[0]);
    nor g2669(n2059 ,n1892 ,n1866);
    nor g2670(n1004 ,n956 ,n992);
    nor g2671(n452 ,n149 ,n102);
    nor g2672(n2694 ,n2615 ,n2666);
    nor g2673(n414 ,n140 ,n349);
    not g2674(n1016 ,n1017);
    xnor g2675(n2322 ,n2220 ,n2041);
    not g2676(n1038 ,n1037);
    xnor g2677(n983 ,n953 ,n20[7]);
    xor g2678(n32[2] ,n1746 ,n1702);
    not g2679(n292 ,n17[3]);
    nor g2680(n1131 ,n946 ,n1064);
    nor g2681(n1104 ,n956 ,n1063);
    nor g2682(n2349 ,n2203 ,n2305);
    or g2683(n3161 ,n3154 ,n3140);
    nor g2684(n2285 ,n1988 ,n2144);
    xnor g2685(n3278 ,n2885 ,n2900);
    not g2686(n1326 ,n1325);
    nor g2687(n3182 ,n3114 ,n3142);
    xnor g2688(n2386 ,n2278 ,n2031);
    xor g2689(n938 ,n973 ,n985);
    nor g2690(n2813 ,n2683 ,n2774);
    nor g2691(n2224 ,n1982 ,n2109);
    not g2692(n1705 ,n1704);
    xnor g2693(n2890 ,n2837 ,n2841);
    nor g2694(n367 ,n266 ,n105);
    nor g2695(n2947 ,n2936 ,n2946);
    nor g2696(n1901 ,n1887 ,n1874);
    xnor g2697(n2800 ,n2640 ,n2759);
    nor g2698(n472 ,n222 ,n102);
    xnor g2699(n2416 ,n2236 ,n1893);
    nor g2700(n2522 ,n2282 ,n2429);
    not g2701(n2963 ,n22[3]);
    not g2702(n3110 ,n3316);
    not g2703(n3113 ,n3283);
    nor g2704(n94 ,n25[4] ,n92);
    or g2705(n362 ,n5[9] ,n335);
    nor g2706(n930 ,n86 ,n85);
    not g2707(n1178 ,n1177);
    nor g2708(n347 ,n108 ,n321);
    not g2709(n2701 ,n2700);
    not g2710(n1956 ,n1955);
    or g2711(n324 ,n115 ,n5[3]);
    nor g2712(n1188 ,n1027 ,n1146);
    dff g2713(.RN(n1), .SN(1'b1), .CK(n0), .D(n601), .Q(n10[2]));
    nor g2714(n1857 ,n1839 ,n1856);
    not g2715(n2984 ,n2983);
    nor g2716(n2743 ,n2660 ,n2715);
    nor g2717(n799 ,n240 ,n653);
    not g2718(n213 ,n21[6]);
    xnor g2719(n2729 ,n2650 ,n2614);
    or g2720(n848 ,n742 ,n674);
    nor g2721(n1951 ,n1890 ,n1870);
    not g2722(n2599 ,n2598);
    or g2723(n917 ,n899 ,n908);
    not g2724(n3083 ,n3262);
    nor g2725(n1945 ,n1890 ,n1866);
    xnor g2726(n2610 ,n2473 ,n2392);
    xnor g2727(n2773 ,n2692 ,n2662);
    not g2728(n274 ,n29[15]);
    not g2729(n140 ,n25[2]);
    nor g2730(n1010 ,n987 ,n980);
    nor g2731(n1330 ,n1256 ,n1312);
    xnor g2732(n332 ,n126 ,n185);
    nor g2733(n381 ,n274 ,n103);
    buf g2734(n10[28], 1'b0);
    nor g2735(n683 ,n110 ,n650);
    not g2736(n2456 ,n2455);
    or g2737(n858 ,n752 ,n676);
    nor g2738(n393 ,n275 ,n105);
    not g2739(n3000 ,n3300);
    or g2740(n910 ,n784 ,n861);
    buf g2741(n12[10], n10[2]);
    nor g2742(n809 ,n119 ,n655);
    nor g2743(n3185 ,n3120 ,n3154);
    or g2744(n3245 ,n3187 ,n3198);
    or g2745(n859 ,n780 ,n778);
    nor g2746(n2035 ,n1867 ,n1877);
    nor g2747(n2683 ,n2530 ,n2621);
    not g2748(n177 ,n928);
    nor g2749(n696 ,n113 ,n661);
    nor g2750(n318 ,n183 ,n18[2]);
    nor g2751(n745 ,n189 ,n667);
    xnor g2752(n1245 ,n1026 ,n1161);
    buf g2753(n10[22], 1'b0);
    nor g2754(n1312 ,n1245 ,n1271);
    not g2755(n192 ,n20[2]);
    nor g2756(n617 ,n252 ,n524);
    nor g2757(n1311 ,n941 ,n1274);
    nor g2758(n3014 ,n3288 ,n3272);
    nor g2759(n1118 ,n946 ,n1063);
    xnor g2760(n2847 ,n2788 ,n2704);
    nor g2761(n2145 ,n2065 ,n1911);
    xnor g2762(n2539 ,n2414 ,n2369);
    nor g2763(n2097 ,n1869 ,n1870);
    dff g2764(.RN(n1), .SN(1'b1), .CK(n0), .D(n533), .Q(n29[8]));
    nor g2765(n1546 ,n1519 ,n1531);
    nor g2766(n1617 ,n1520 ,n1552);
    dff g2767(.RN(n1), .SN(1'b1), .CK(n0), .D(n843), .Q(n20[5]));
    or g2768(n31[9] ,n3233 ,n3254);
    nor g2769(n1013 ,n947 ,n992);
    buf g2770(n9[12], 1'b0);
    nor g2771(n458 ,n143 ,n102);
    or g2772(n898 ,n802 ,n871);
    xnor g2773(n2736 ,n2642 ,n2596);
    or g2774(n529 ,n381 ,n466);
    not g2775(n133 ,n31[13]);
    nor g2776(n970 ,n20[2] ,n20[1]);
    not g2777(n110 ,n6[4]);
    nor g2778(n411 ,n229 ,n349);
    nor g2779(n2863 ,n2833 ,n2858);
    or g2780(n558 ,n521 ,n495);
    nor g2781(n1508 ,n1466 ,n1507);
    xnor g2782(n2264 ,n2021 ,n1899);
    not g2783(n1758 ,n1757);
    not g2784(n1197 ,n1196);
    not g2785(n2554 ,n2553);
    xnor g2786(n1711 ,n1638 ,n1640);
    or g2787(n862 ,n786 ,n785);
    xnor g2788(n1715 ,n1585 ,n1649);
    nor g2789(n750 ,n186 ,n660);
    not g2790(n3125 ,n3281);
    nor g2791(n2380 ,n2199 ,n2298);
    nor g2792(n1623 ,n1519 ,n1551);
    nor g2793(n2621 ,n2532 ,n2562);
    not g2794(n2056 ,n2055);
    buf g2795(n12[3], 1'b0);
    nor g2796(n418 ,n287 ,n347);
    nor g2797(n670 ,n107 ,n650);
    buf g2798(n12[26], 1'b0);
    nor g2799(n2160 ,n1928 ,n2040);
    not g2800(n2042 ,n2041);
    nor g2801(n1504 ,n1503 ,n1489);
    nor g2802(n2215 ,n1960 ,n1920);
    or g2803(n3162 ,n3154 ,n3136);
    nor g2804(n2946 ,n2945 ,n2934);
    not g2805(n984 ,n983);
    nor g2806(n45 ,n40 ,n44);
    buf g2807(n13[17], 1'b0);
    not g2808(n214 ,n23[4]);
    not g2809(n1974 ,n1973);
    not g2810(n2793 ,n2792);
    nor g2811(n1320 ,n1231 ,n1253);
    nor g2812(n2614 ,n2512 ,n2547);
    nor g2813(n509 ,n138 ,n346);
    or g2814(n541 ,n382 ,n355);
    not g2815(n1765 ,n1764);
    nor g2816(n697 ,n109 ,n661);
    nor g2817(n469 ,n278 ,n104);
    not g2818(n1948 ,n1947);
    xor g2819(n2432 ,n2242 ,n1995);
    dff g2820(.RN(n1), .SN(1'b1), .CK(n0), .D(n849), .Q(n19[7]));
    nor g2821(n378 ,n158 ,n105);
    nor g2822(n2709 ,n2675 ,n2662);
    nor g2823(n2356 ,n1954 ,n2271);
    nor g2824(n2294 ,n2136 ,n2158);
    not g2825(n1828 ,n1827);
    nor g2826(n2506 ,n2320 ,n2440);
    nor g2827(n1668 ,n1569 ,n1618);
    nor g2828(n1390 ,n1260 ,n1372);
    or g2829(n884 ,n810 ,n809);
    or g2830(n600 ,n430 ,n509);
    nor g2831(n2019 ,n1887 ,n1861);
    nor g2832(n2015 ,n1883 ,n1875);
    or g2833(n31[5] ,n3217 ,n3256);
    nor g2834(n2579 ,n2444 ,n2507);
    nor g2835(n1083 ,n959 ,n1034);
    nor g2836(n491 ,n169 ,n102);
    nor g2837(n416 ,n251 ,n349);
    xnor g2838(n2588 ,n2477 ,n2329);
    not g2839(n1424 ,n1423);
    or g2840(n551 ,n391 ,n452);
    nor g2841(n2911 ,n2864 ,n2893);
    xnor g2842(n1398 ,n1347 ,n1304);
    not g2843(n1368 ,n1367);
    nor g2844(n97 ,n25[5] ,n95);
    not g2845(n2923 ,n2922);
    nor g2846(n1935 ,n1884 ,n1878);
    xor g2847(n941 ,n1025 ,n1150);
    xnor g2848(n2870 ,n2823 ,n2783);
    nor g2849(n2377 ,n2210 ,n2315);
    nor g2850(n1172 ,n1068 ,n1125);
    not g2851(n2084 ,n2083);
    nor g2852(n2896 ,n2869 ,n2881);
    xnor g2853(n2246 ,n1969 ,n1967);
    nor g2854(n1619 ,n1520 ,n1554);
    nor g2855(n2337 ,n2188 ,n2304);
    xnor g2856(n3299 ,n1487 ,n1500);
    nor g2857(n2747 ,n2624 ,n2700);
    nor g2858(n1122 ,n947 ,n1089);
    nor g2859(n2130 ,n1867 ,n1875);
    not g2860(n1204 ,n1203);
    nor g2861(n3041 ,n3012 ,n3040);
    not g2862(n2957 ,n22[4]);
    not g2863(n2891 ,n2890);
    nor g2864(n3169 ,n3097 ,n3141);
    xnor g2865(n2474 ,n2337 ,n2348);
    nor g2866(n1362 ,n1190 ,n1331);
    nor g2867(n1415 ,n1278 ,n1390);
    xnor g2868(n3023 ,n3303 ,n3287);
    xnor g2869(n2979 ,n22[5] ,n23[5]);
    xnor g2870(n2608 ,n2475 ,n2465);
    nor g2871(n2287 ,n2103 ,n2167);
    nor g2872(n307 ,n18[0] ,n18[1]);
    not g2873(n157 ,n28[10]);
    xnor g2874(n2691 ,n2390 ,n2602);
    nor g2875(n2345 ,n2189 ,n2293);
    nor g2876(n1544 ,n1521 ,n1538);
    nor g2877(n1432 ,n1385 ,n1408);
    nor g2878(n2715 ,n2610 ,n2659);
    not g2879(n2768 ,n2767);
    buf g2880(n10[16], 1'b0);
    not g2881(n2068 ,n2067);
    or g2882(n901 ,n821 ,n893);
    nor g2883(n2161 ,n2081 ,n2087);
    not g2884(n1992 ,n1991);
    not g2885(n47 ,n25[4]);
    nor g2886(n380 ,n148 ,n103);
    not g2887(n126 ,n28[6]);
    not g2888(n2086 ,n2085);
    xnor g2889(n1352 ,n1292 ,n1168);
    or g2890(n656 ,n523 ,n645);
    not g2891(n3119 ,n3294);
    not g2892(n2138 ,n2137);
    not g2893(n3129 ,n3291);
    not g2894(n2597 ,n2596);
    buf g2895(n11[13], 1'b0);
    xnor g2896(n2596 ,n2474 ,n2412);
    nor g2897(n1055 ,n957 ,n1036);
    dff g2898(.RN(n1), .SN(1'b1), .CK(n0), .D(n535), .Q(n29[12]));
    nor g2899(n368 ,n157 ,n105);
    nor g2900(n3192 ,n3129 ,n3141);
    nor g2901(n1322 ,n1175 ,n1299);
    not g2902(n1660 ,n1659);
    not g2903(n2113 ,n2112);
    not g2904(n144 ,n31[6]);
    not g2905(n2393 ,n2392);
    dff g2906(.RN(n1), .SN(1'b1), .CK(n0), .D(n885), .Q(n23[6]));
    dff g2907(.RN(n1), .SN(1'b1), .CK(n0), .D(n536), .Q(n29[11]));
    not g2908(n87 ,n86);
    not g2909(n2962 ,n23[5]);
    or g2910(n3141 ,n27[1] ,n27[0]);
    dff g2911(.RN(n1), .SN(1'b1), .CK(n0), .D(n599), .Q(n10[4]));
    nor g2912(n1693 ,n1641 ,n1639);
    xnor g2913(n1024 ,n1010 ,n993);
    dff g2914(.RN(n1), .SN(1'b1), .CK(n0), .D(n831), .Q(n21[7]));
    buf g2915(n12[4], 1'b0);
    not g2916(n148 ,n29[2]);
    nor g2917(n1041 ,n958 ,n1038);
    nor g2918(n2927 ,n2903 ,n2890);
    not g2919(n2098 ,n2097);
    nor g2920(n2106 ,n1880 ,n1877);
    xnor g2921(n2271 ,n2008 ,n1977);
    nor g2922(n2720 ,n2686 ,n2657);
    buf g2923(n13[1], 1'b0);
    not g2924(n1964 ,n1963);
    xnor g2925(n1200 ,n1017 ,n1170);
    not g2926(n196 ,n22[0]);
    nor g2927(n358 ,n104 ,n336);
    buf g2928(n9[27], 1'b0);
    nor g2929(n787 ,n224 ,n653);
    not g2930(n3091 ,n3272);
    nor g2931(n801 ,n191 ,n665);
    not g2932(n2764 ,n2763);
    nor g2933(n2362 ,n2225 ,n2267);
    not g2934(n2684 ,n2683);
    not g2935(n3090 ,n3303);
    nor g2936(n1989 ,n1864 ,n1876);
    nor g2937(n412 ,n245 ,n349);
    xnor g2938(n2662 ,n2544 ,n2471);
    nor g2939(n3179 ,n3092 ,n3141);
    not g2940(n2399 ,n2398);
    xnor g2941(n2727 ,n2604 ,n2654);
    or g2942(n629 ,n361 ,n628);
    buf g2943(n17[6], 1'b0);
    not g2944(n218 ,n20[3]);
    xnor g2945(n2267 ,n1986 ,n1989);
    or g2946(n833 ,n729 ,n688);
    nor g2947(n1020 ,n994 ,n1006);
    xor g2948(n32[7] ,n1845 ,n1851);
    nor g2949(n773 ,n124 ,n653);
    nor g2950(n401 ,n272 ,n103);
    xnor g2951(n2402 ,n2249 ,n2093);
    not g2952(n2080 ,n2079);
    or g2953(n881 ,n759 ,n677);
    dff g2954(.RN(n1), .SN(1'b1), .CK(n0), .D(n556), .Q(n29[14]));
    dff g2955(.RN(n1), .SN(1'b1), .CK(n0), .D(n888), .Q(n23[4]));
    nor g2956(n1548 ,n1522 ,n1531);
    nor g2957(n1541 ,n1521 ,n1533);
    not g2958(n2961 ,n23[0]);
    xnor g2959(n993 ,n20[5] ,n21[5]);
    xor g2960(n3307 ,n2981 ,n2986);
    not g2961(n1875 ,n22[0]);
    nor g2962(n3177 ,n3128 ,n3141);
    nor g2963(n2632 ,n2529 ,n2577);
    not g2964(n2503 ,n2502);
    xnor g2965(n3035 ,n3300 ,n3284);
    nor g2966(n2488 ,n2380 ,n2448);
    nor g2967(n2199 ,n2068 ,n1934);
    nor g2968(n1054 ,n947 ,n1036);
    not g2969(n158 ,n26[3]);
    xnor g2970(n1288 ,n1209 ,n1235);
    not g2971(n2766 ,n2765);
    or g2972(n42 ,n30[2] ,n30[0]);
    not g2973(n1519 ,n24[0]);
    or g2974(n863 ,n788 ,n787);
    nor g2975(n3130 ,n3317 ,n32[8]);
    not g2976(n248 ,n29[1]);
    nor g2977(n425 ,n228 ,n347);
    or g2978(n577 ,n440 ,n485);
    nor g2979(n2152 ,n1947 ,n2035);
    nor g2980(n638 ,n346 ,n637);
    xnor g2981(n2763 ,n2690 ,n2608);
    not g2982(n1876 ,n22[1]);
    nor g2983(n399 ,n244 ,n105);
    xnor g2984(n2796 ,n2726 ,n2740);
    nor g2985(n1106 ,n949 ,n1063);
    nor g2986(n972 ,n20[0] ,n21[0]);
    nor g2987(n1111 ,n957 ,n1062);
    nor g2988(n2644 ,n2553 ,n2596);
    xnor g2989(n3322 ,n3030 ,n3022);
    xnor g2990(n1749 ,n1711 ,n1728);
    or g2991(n876 ,n756 ,n707);
    nor g2992(n1680 ,n1628 ,n1642);
    not g2993(n2016 ,n2015);
    xnor g2994(n3302 ,n1474 ,n1506);
    not g2995(n1462 ,n1461);
    or g2996(n644 ,n322 ,n642);
    nor g2997(n1143 ,n1055 ,n1108);
    nor g2998(n1647 ,n1567 ,n1620);
    nor g2999(n1018 ,n996 ,n1007);
    nor g3000(n1433 ,n1298 ,n1405);
    xnor g3001(n2241 ,n2083 ,n2019);
    nor g3002(n736 ,n200 ,n662);
    nor g3003(n793 ,n150 ,n653);
    not g3004(n2603 ,n2602);
    nor g3005(n1893 ,n1864 ,n1872);
    not g3006(n2338 ,n2337);
    nor g3007(n1820 ,n1764 ,n1796);
    not g3008(n1944 ,n1943);
    xnor g3009(n2789 ,n2702 ,n2760);
    nor g3010(n86 ,n82 ,n79);
    nor g3011(n2816 ,n2753 ,n2769);
    not g3012(n171 ,n936);
    or g3013(n861 ,n616 ,n783);
    not g3014(n199 ,n23[0]);
    nor g3015(n1575 ,n1520 ,n1532);
    xnor g3016(n3290 ,n1294 ,n1246);
    xnor g3017(n1209 ,n1142 ,n1028);
    or g3018(n643 ,n523 ,n641);
    xnor g3019(n1348 ,n1287 ,n1248);
    nor g3020(n1500 ,n1480 ,n1499);
    not g3021(n3104 ,n3314);
    not g3022(n1195 ,n1194);
    not g3023(n2647 ,n2646);
    not g3024(n659 ,n660);
    not g3025(n291 ,n29[11]);
    nor g3026(n616 ,n160 ,n524);
    nor g3027(n1246 ,n1066 ,n1185);
    or g3028(n645 ,n324 ,n642);
    not g3029(n1298 ,n1297);
    nor g3030(n1044 ,n957 ,n1034);
    or g3031(n539 ,n370 ,n469);
    nor g3032(n2873 ,n2764 ,n2847);
    nor g3033(n1279 ,n1169 ,n1201);
    nor g3034(n2303 ,n1984 ,n2159);
    nor g3035(n1127 ,n946 ,n1089);
    not g3036(n2340 ,n2339);
    not g3037(n210 ,n28[5]);
    nor g3038(n3242 ,n3146 ,n3161);
    not g3039(n1263 ,n1262);
    xnor g3040(n1385 ,n1321 ,n1262);
    or g3041(n544 ,n386 ,n455);
    or g3042(n582 ,n392 ,n462);
    buf g3043(n11[27], n10[11]);
    nor g3044(n2973 ,n2959 ,n2956);
    not g3045(n3069 ,n32[11]);
    not g3046(n2631 ,n2630);
    dff g3047(.RN(n1), .SN(1'b1), .CK(n0), .D(n830), .Q(n22[0]));
    xnor g3048(n1404 ,n1345 ,n1282);
    xnor g3049(n1286 ,n1180 ,n1237);
    nor g3050(n505 ,n153 ,n346);
    nor g3051(n2435 ,n2351 ,n2358);
    nor g3052(n2560 ,n2445 ,n2493);
    xnor g3053(n2412 ,n2257 ,n2118);
    not g3054(n1701 ,n1700);
    nor g3055(n2663 ,n2572 ,n2617);
    not g3056(n149 ,n31[5]);
    nor g3057(n1305 ,n1188 ,n1252);
    xnor g3058(n1463 ,n1419 ,n1369);
    dff g3059(.RN(n1), .SN(1'b1), .CK(n0), .D(n876), .Q(n24[4]));
    not g3060(n2993 ,n2992);
    xnor g3061(n1327 ,n1167 ,n1283);
    xnor g3062(n981 ,n951 ,n21[1]);
    or g3063(n636 ,n309 ,n634);
    nor g3064(n927 ,n94 ,n95);
    not g3065(n663 ,n664);
    nor g3066(n2169 ,n1959 ,n1919);
    xnor g3067(n1371 ,n1296 ,n1217);
    or g3068(n3253 ,n3176 ,n3237);
    not g3069(n2611 ,n2610);
    nor g3070(n356 ,n104 ,n327);
    xnor g3071(n2420 ,n2251 ,n1991);
    nor g3072(n2305 ,n2121 ,n2151);
    nor g3073(n508 ,n151 ,n346);
    nor g3074(n1335 ,n1016 ,n1317);
    xnor g3075(n3033 ,n3294 ,n3278);
    xnor g3076(n2239 ,n2089 ,n2047);
    not g3077(n3118 ,n3280);
    xnor g3078(n1215 ,n1164 ,n1028);
    nor g3079(n2875 ,n2791 ,n2841);
    dff g3080(.RN(n1), .SN(1'b1), .CK(n0), .D(n914), .Q(n9[0]));
    not g3081(n3107 ,n3321);
    not g3082(n2601 ,n2600);
    not g3083(n2735 ,n2734);
    nor g3084(n2775 ,n2714 ,n2749);
    nor g3085(n434 ,n147 ,n105);
    not g3086(n102 ,n105);
    dff g3087(.RN(n1), .SN(1'b1), .CK(n0), .D(n575), .Q(n28[6]));
    nor g3088(n485 ,n179 ,n104);
    not g3089(n1787 ,n1786);
    not g3090(n1928 ,n1927);
    xnor g3091(n1827 ,n1790 ,n1766);
    nor g3092(n1563 ,n1521 ,n1530);
    xnor g3093(n2502 ,n2233 ,n2381);
    not g3094(n2649 ,n2648);
    not g3095(n33 ,n30[4]);
    or g3096(n839 ,n733 ,n671);
    buf g3097(n13[16], 1'b0);
    xnor g3098(n1675 ,n1621 ,n1577);
    not g3099(n3103 ,n32[6]);
    xnor g3100(n986 ,n963 ,n20[6]);
    or g3101(n888 ,n764 ,n713);
    nor g3102(n386 ,n262 ,n103);
    nor g3103(n726 ,n196 ,n651);
    nor g3104(n2151 ,n1943 ,n2075);
    xnor g3105(n2537 ,n2428 ,n2085);
    not g3106(n276 ,n10[12]);
    xnor g3107(n1396 ,n1352 ,n1332);
    not g3108(n56 ,n30[4]);
    nor g3109(n1727 ,n1652 ,n1683);
    xnor g3110(n2732 ,n2638 ,n2500);
    not g3111(n2958 ,n22[5]);
    or g3112(n548 ,n402 ,n459);
    nor g3113(n3056 ,n3031 ,n3055);
    not g3114(n3112 ,n3279);
    not g3115(n201 ,n21[3]);
    nor g3116(n778 ,n195 ,n655);
    not g3117(n163 ,n31[12]);
    nor g3118(n2178 ,n1894 ,n2046);
    nor g3119(n1370 ,n1308 ,n1337);
    xnor g3120(n2388 ,n2256 ,n2025);
    nor g3121(n622 ,n283 ,n524);
    nor g3122(n372 ,n270 ,n105);
    dff g3123(.RN(n1), .SN(1'b1), .CK(n0), .D(n580), .Q(n25[6]));
    nor g3124(n775 ,n187 ,n652);
    not g3125(n1864 ,n20[5]);
    nor g3126(n1722 ,n1666 ,n1694);
    buf g3127(n9[22], 1'b0);
    nor g3128(n1490 ,n1434 ,n1477);
    buf g3129(n12[19], n10[11]);
    dff g3130(.RN(n1), .SN(1'b1), .CK(n0), .D(n583), .Q(n25[4]));
    nor g3131(n2290 ,n2098 ,n2145);
    nor g3132(n2828 ,n2730 ,n2798);
    nor g3133(n1377 ,n1338 ,n1367);
    xnor g3134(n2400 ,n2246 ,n2122);
    nor g3135(n1158 ,n1056 ,n1104);
    not g3136(n1604 ,n1603);
    not g3137(n156 ,n29[5]);
    xnor g3138(n997 ,n20[1] ,n21[1]);
    not g3139(n208 ,n28[2]);
    nor g3140(n504 ,n145 ,n346);
    not g3141(n2403 ,n2402);
    nor g3142(n3152 ,n3107 ,n3070);
    not g3143(n184 ,n18[0]);
    nor g3144(n369 ,n232 ,n103);
    or g3145(n538 ,n439 ,n352);
    xnor g3146(n1673 ,n1599 ,n1579);
    or g3147(n834 ,n774 ,n773);
    dff g3148(.RN(n1), .SN(1'b1), .CK(n0), .D(n874), .Q(n24[5]));
    xnor g3149(n32[11] ,n1805 ,n1859);
    nor g3150(n2079 ,n1871 ,n1873);
    or g3151(n632 ,n304 ,n627);
    dff g3152(.RN(n1), .SN(1'b1), .CK(n0), .D(n551), .Q(n28[5]));
    nor g3153(n1814 ,n1779 ,n1802);
    nor g3154(n615 ,n288 ,n436);
    nor g3155(n1947 ,n1880 ,n1881);
    not g3156(n1920 ,n1919);
    or g3157(n875 ,n804 ,n803);
    nor g3158(n385 ,n164 ,n347);
    nor g3159(n2898 ,n2828 ,n2865);
    nor g3160(n2175 ,n1899 ,n2021);
    xnor g3161(n1187 ,n1026 ,n1115);
    not g3162(n2370 ,n2369);
    nor g3163(n2194 ,n2030 ,n1914);
    not g3164(n257 ,n9[4]);
    xnor g3165(n3295 ,n1456 ,n1490);
    or g3166(n555 ,n435 ,n465);
    not g3167(n123 ,n24[3]);
    nor g3168(n3138 ,n3315 ,n32[10]);
    not g3169(n2427 ,n2426);
    nor g3170(n2209 ,n2074 ,n1904);
    or g3171(n841 ,n735 ,n692);
    xnor g3172(n2392 ,n2263 ,n2091);
    nor g3173(n2291 ,n1976 ,n2149);
    not g3174(n954 ,n21[0]);
    not g3175(n2082 ,n2081);
    not g3176(n1934 ,n1933);
    xnor g3177(n2482 ,n2339 ,n2347);
    xnor g3178(n3026 ,n3292 ,n3276);
    dff g3179(.RN(n1), .SN(1'b1), .CK(n0), .D(n526), .Q(n30[0]));
    nor g3180(n1440 ,n1394 ,n1437);
    not g3181(n2782 ,n2781);
    buf g3182(n13[20], 1'b0);
    not g3183(n1512 ,n23[6]);
    not g3184(n242 ,n29[0]);
    or g3185(n566 ,n371 ,n474);
    not g3186(n1748 ,n1747);
    nor g3187(n2660 ,n2571 ,n2619);
    or g3188(n3155 ,n3099 ,n27[0]);
    nor g3189(n2341 ,n2197 ,n2310);
    not g3190(n2024 ,n2023);
    xnor g3191(n2725 ,n2663 ,n2624);
    nor g3192(n2520 ,n2343 ,n2419);
    not g3193(n261 ,n26[15]);
    dff g3194(.RN(n1), .SN(1'b1), .CK(n0), .D(n872), .Q(n24[7]));
    or g3195(n3247 ,n3205 ,n3235);
    dff g3196(.RN(n1), .SN(1'b1), .CK(n0), .D(n587), .Q(n10[15]));
    or g3197(n590 ,n446 ,n480);
    nor g3198(n3194 ,n3127 ,n3142);
    nor g3199(n792 ,n209 ,n666);
    nor g3200(n2722 ,n2623 ,n2665);
    nor g3201(n1156 ,n1059 ,n1116);
    nor g3202(n1858 ,n1830 ,n1857);
    nor g3203(n2201 ,n1948 ,n2036);
    nor g3204(n1965 ,n1871 ,n1877);
    not g3205(n1303 ,n943);
    not g3206(n1522 ,n24[1]);
    or g3207(n899 ,n808 ,n879);
    nor g3208(n2165 ,n1915 ,n2049);
    buf g3209(n13[0], 1'b0);
    dff g3210(.RN(n1), .SN(1'b1), .CK(n0), .D(n561), .Q(n26[12]));
    nor g3211(n1831 ,n1777 ,n1810);
    dff g3212(.RN(n1), .SN(1'b1), .CK(n0), .D(n825), .Q(n22[3]));
    not g3213(n1357 ,n1356);
    nor g3214(n408 ,n264 ,n103);
    xnor g3215(n1751 ,n1706 ,n1715);
    or g3216(n1533 ,n1528 ,n1524);
    nor g3217(n782 ,n193 ,n654);
    xnor g3218(n2455 ,n2266 ,n1949);
    nor g3219(n2309 ,n2132 ,n2155);
    nor g3220(n2616 ,n2388 ,n2549);
    not g3221(n2562 ,n2561);
    not g3222(n1902 ,n1901);
    nor g3223(n1467 ,n1442 ,n1448);
    nor g3224(n2217 ,n2016 ,n2140);
    nor g3225(n2297 ,n1998 ,n2146);
    or g3226(n1988 ,n1882 ,n1870);
    nor g3227(n1138 ,n1047 ,n1107);
    nor g3228(n973 ,n20[1] ,n21[1]);
    xnor g3229(n2504 ,n2245 ,n2349);
    xnor g3230(n2590 ,n2480 ,n2354);
    not g3231(n185 ,n19[6]);
    xnor g3232(n1747 ,n1708 ,n1717);
    or g3233(n610 ,n26[15] ,n363);
    nor g3234(n1799 ,n1582 ,n1786);
    nor g3235(n2141 ,n1927 ,n2039);
    xnor g3236(n2258 ,n1939 ,n2037);
    nor g3237(n2877 ,n2817 ,n2846);
    xnor g3238(n2646 ,n2541 ,n2561);
    xnor g3239(n2977 ,n22[1] ,n23[1]);
    nor g3240(n3064 ,n3018 ,n3063);
    nor g3241(n672 ,n107 ,n648);
    xnor g3242(n3030 ,n3273 ,n3289);
    dff g3243(.RN(n1), .SN(1'b1), .CK(n0), .D(n894), .Q(n23[0]));
    not g3244(n3006 ,n3284);
    not g3245(n132 ,n31[14]);
    not g3246(n2907 ,n2906);
    or g3247(n879 ,n620 ,n807);
    buf g3248(n13[25], n10[1]);
    nor g3249(n1587 ,n1520 ,n1556);
    not g3250(n1887 ,n20[2]);
    not g3251(n112 ,n6[5]);
    nor g3252(n1472 ,n1377 ,n1440);
    xnor g3253(n1346 ,n1176 ,n1299);
    or g3254(n2114 ,n1890 ,n1862);
    or g3255(n31[8] ,n3229 ,n3252);
    nor g3256(n1943 ,n1880 ,n1861);
    nor g3257(n2529 ,n2405 ,n2421);
    nor g3258(n2137 ,n1871 ,n1872);
    or g3259(n634 ,n310 ,n630);
    buf g3260(n13[24], n10[0]);
    nor g3261(n2935 ,n2904 ,n2919);
    or g3262(n573 ,n378 ,n479);
    nor g3263(n1594 ,n1521 ,n1555);
    nor g3264(n1939 ,n1867 ,n1873);
    nor g3265(n2183 ,n1906 ,n1930);
    nor g3266(n1986 ,n1880 ,n1875);
    not g3267(n1238 ,n1237);
    not g3268(n162 ,n31[0]);
    not g3269(n1868 ,n23[6]);
    nor g3270(n459 ,n145 ,n102);
    xnor g3271(n2279 ,n2126 ,n1999);
    xor g3272(n32[6] ,n1836 ,n1849);
    nor g3273(n1072 ,n947 ,n1040);
    not g3274(n1879 ,n21[5]);
    buf g3275(n12[16], n10[8]);
    xor g3276(n1769 ,n1738 ,n1739);
    not g3277(n1910 ,n1909);
    nor g3278(n2374 ,n2192 ,n2294);
    nor g3279(n515 ,n172 ,n348);
    not g3280(n1824 ,n1823);
    or g3281(n866 ,n792 ,n791);
    xnor g3282(n2235 ,n1945 ,n1935);
    or g3283(n867 ,n794 ,n793);
    xor g3284(n939 ,n968 ,n986);
    nor g3285(n2343 ,n2205 ,n2308);
    nor g3286(n2992 ,n2974 ,n2991);
    nor g3287(n2189 ,n2038 ,n1940);
    nor g3288(n2491 ,n2459 ,n2394);
    nor g3289(n3240 ,n3148 ,n3163);
    dff g3290(.RN(n1), .SN(1'b1), .CK(n0), .D(n591), .Q(n10[12]));
    nor g3291(n395 ,n242 ,n105);
    or g3292(n3218 ,n3201 ,n3214);
    nor g3293(n433 ,n239 ,n347);
    not g3294(n3109 ,n3315);
    not g3295(n1687 ,n1686);
    nor g3296(n978 ,n955 ,n954);
    not g3297(n279 ,n29[4]);
    or g3298(n3158 ,n3154 ,n3132);
    dff g3299(.RN(n1), .SN(1'b1), .CK(n0), .D(n578), .Q(n25[7]));
    nor g3300(n3049 ,n3015 ,n3048);
    not g3301(n1889 ,n23[5]);
    dff g3302(.RN(n1), .SN(1'b1), .CK(n0), .D(n629), .Q(n18[2]));
    xnor g3303(n1847 ,n1823 ,n1814);
    nor g3304(n932 ,n76 ,n77);
    nor g3305(n3018 ,n2998 ,n3005);
    dff g3306(.RN(n1), .SN(1'b1), .CK(n0), .D(n829), .Q(n22[1]));
    nor g3307(n1412 ,n1332 ,n1391);
    not g3308(n1878 ,n23[1]);
    nor g3309(n2987 ,n2981 ,n2986);
    nor g3310(n1315 ,n1242 ,n1273);
    or g3311(n31[12] ,n3218 ,n3234);
    or g3312(n893 ,n816 ,n815);
    not g3313(n289 ,n26[11]);
    nor g3314(n806 ,n123 ,n653);
    or g3315(n31[15] ,n3203 ,n3219);
    nor g3316(n2762 ,n2622 ,n2759);
    not g3317(n1871 ,n20[4]);
    not g3318(n200 ,n20[6]);
    xnor g3319(n2480 ,n2325 ,n2327);
    not g3320(n1523 ,n3270);
    xnor g3321(n2839 ,n2796 ,n2755);
    xnor g3322(n2702 ,n2585 ,n2506);
    nor g3323(n1921 ,n1865 ,n1872);
    dff g3324(.RN(n1), .SN(1'b1), .CK(n0), .D(n552), .Q(n28[4]));
    nor g3325(n1955 ,n1879 ,n1868);
    xor g3326(n3285 ,n2916 ,n2951);
    or g3327(n550 ,n429 ,n486);
    nor g3328(n1638 ,n1542 ,n1594);
    nor g3329(n3172 ,n3112 ,n3142);
    nor g3330(n1983 ,n1890 ,n1891);
    nor g3331(n1496 ,n1495 ,n1452);
    nor g3332(n1782 ,n1738 ,n1754);
    or g3333(n3225 ,n3172 ,n3207);
    nor g3334(n1192 ,n1026 ,n1150);
    not g3335(n3100 ,n32[12]);
    nor g3336(n522 ,n919 ,n337);
    nor g3337(n2693 ,n2560 ,n2669);
    not g3338(n1210 ,n1209);
    nor g3339(n1073 ,n957 ,n1032);
    xnor g3340(n1239 ,n1026 ,n1155);
    xnor g3341(n1037 ,n939 ,n1020);
    xnor g3342(n3280 ,n2929 ,n2941);
    xnor g3343(n2604 ,n2483 ,n2376);
    nor g3344(n1819 ,n1765 ,n1795);
    xnor g3345(n2802 ,n2724 ,n2757);
    nor g3346(n2834 ,n2755 ,n2797);
    or g3347(n563 ,n522 ,n364);
    nor g3348(n2861 ,n2800 ,n2854);
    xnor g3349(n2384 ,n2277 ,n1937);
    not g3350(n2580 ,n2579);
    xor g3351(n3310 ,n2976 ,n2992);
    nor g3352(n3147 ,n3105 ,n3073);
    buf g3353(n12[28], 1'b0);
    xnor g3354(n2251 ,n2059 ,n2017);
    nor g3355(n1793 ,n1762 ,n1785);
    xnor g3356(n1837 ,n1776 ,n1810);
    xnor g3357(n3300 ,n1492 ,n1502);
    xor g3358(n2262 ,n1985 ,n2069);
    nor g3359(n2468 ,n2319 ,n2323);
    not g3360(n57 ,n30[3]);
    xnor g3361(n2929 ,n2890 ,n2902);
    or g3362(n31[1] ,n3226 ,n3250);
    nor g3363(n1909 ,n1879 ,n1889);
    nor g3364(n743 ,n112 ,n657);
    nor g3365(n1677 ,n1625 ,n1668);
    nor g3366(n3139 ,n3318 ,n32[7]);
    nor g3367(n1570 ,n1519 ,n1532);
    nor g3368(n3062 ,n3020 ,n3061);
    not g3369(n1236 ,n1235);
    not g3370(n1516 ,n3264);
    nor g3371(n2623 ,n2389 ,n2550);
    nor g3372(n2085 ,n1883 ,n1876);
    nor g3373(n1337 ,n1285 ,n1309);
    nor g3374(n2819 ,n2745 ,n2777);
    not g3375(n1193 ,n1192);
    not g3376(n1600 ,n1599);
    nor g3377(n498 ,n132 ,n346);
    nor g3378(n2071 ,n1892 ,n1870);
    not g3379(n181 ,n19[7]);
    xnor g3380(n2557 ,n2384 ,n2218);
    not g3381(n118 ,n5[3]);
    nor g3382(n1336 ,n1176 ,n1300);
    xor g3383(n3266 ,n20[2] ,n21[2]);
    nor g3384(n1278 ,n1179 ,n1238);
    nor g3385(n746 ,n117 ,n667);
    nor g3386(n454 ,n132 ,n102);
    nor g3387(n2995 ,n2968 ,n2994);
    or g3388(n350 ,n17[2] ,n347);
    or g3389(n579 ,n419 ,n357);
    or g3390(n351 ,n18[2] ,n330);
    xnor g3391(n2930 ,n2906 ,n2886);
    dff g3392(.RN(n1), .SN(1'b1), .CK(n0), .D(n559), .Q(n26[15]));
    buf g3393(n13[28], n10[4]);
    xnor g3394(n2843 ,n2789 ,n2771);
    nor g3395(n2184 ,n2024 ,n1966);
    nor g3396(n1723 ,n1704 ,n1687);
    nor g3397(n1015 ,n959 ,n992);
    or g3398(n609 ,n5[6] ,n362);
    nor g3399(n1154 ,n1053 ,n1132);
    or g3400(n3234 ,n3193 ,n3191);
    nor g3401(n2306 ,n2169 ,n2231);
    xnor g3402(n2939 ,n2920 ,n2911);
    or g3403(n825 ,n723 ,n684);
    nor g3404(n1071 ,n948 ,n1040);
    nor g3405(n936 ,n64 ,n65);
    nor g3406(n1688 ,n1583 ,n1635);
    nor g3407(n1067 ,n960 ,n1040);
    dff g3408(.RN(n1), .SN(1'b1), .CK(n0), .D(n853), .Q(n27[0]));
    dff g3409(.RN(n1), .SN(1'b1), .CK(n0), .D(n592), .Q(n10[11]));
    nor g3410(n2852 ,n2761 ,n2831);
    nor g3411(n76 ,n30[6] ,n74);
    not g3412(n78 ,n25[6]);
    not g3413(n1885 ,n21[2]);
    not g3414(n959 ,n3311);
    nor g3415(n1009 ,n986 ,n982);
    nor g3416(n1760 ,n1690 ,n1745);
    not g3417(n1918 ,n1917);
    not g3418(n84 ,n25[2]);
    nor g3419(n2313 ,n2138 ,n2152);
    nor g3420(n1829 ,n1819 ,n1816);
    not g3421(n1622 ,n1621);
    xnor g3422(n1753 ,n1712 ,n1727);
    not g3423(n2342 ,n2341);
    xnor g3424(n2549 ,n2387 ,n2373);
    nor g3425(n2467 ,n2300 ,n2364);
    nor g3426(n1803 ,n1724 ,n1773);
    nor g3427(n1085 ,n959 ,n1040);
    nor g3428(n2177 ,n1955 ,n1963);
    nor g3429(n2331 ,n2191 ,n2316);
    buf g3430(n13[21], 1'b0);
    nor g3431(n2075 ,n1867 ,n1872);
    nor g3432(n2093 ,n1879 ,n1891);
    not g3433(n3078 ,n3284);
    xnor g3434(n1241 ,n1026 ,n1165);
    not g3435(n1202 ,n1201);
    nor g3436(n738 ,n191 ,n662);
    not g3437(n2389 ,n2388);
    xnor g3438(n1846 ,n1827 ,n1817);
    nor g3439(n1690 ,n1549 ,n1654);
    nor g3440(n2988 ,n2970 ,n2987);
    nor g3441(n752 ,n187 ,n660);
    xnor g3442(n334 ,n198 ,n181);
    not g3443(n1922 ,n1921);
    dff g3444(.RN(n1), .SN(1'b1), .CK(n0), .D(n846), .Q(n20[2]));
    nor g3445(n1661 ,n1562 ,n1612);
    or g3446(n589 ,n420 ,n499);
    nor g3447(n1856 ,n1844 ,n1855);
    not g3448(n1174 ,n1173);
    or g3449(n3255 ,n3197 ,n3244);
    not g3450(n151 ,n31[4]);
    or g3451(n871 ,n619 ,n801);
    or g3452(n850 ,n744 ,n699);
    nor g3453(n1498 ,n1465 ,n1497);
    nor g3454(n2055 ,n1863 ,n1870);
    or g3455(n874 ,n755 ,n743);
    nor g3456(n1651 ,n1576 ,n1598);
    buf g3457(n10[23], 1'b0);
    dff g3458(.RN(n1), .SN(1'b1), .CK(n0), .D(n850), .Q(n19[6]));
    nor g3459(n374 ,n136 ,n105);
    nor g3460(n1046 ,n946 ,n1034);
    nor g3461(n2101 ,n1869 ,n1862);
    nor g3462(n2196 ,n2080 ,n2056);
    nor g3463(n2289 ,n2096 ,n2176);
    or g3464(n625 ,n615 ,n612);
    not g3465(n2092 ,n2091);
    nor g3466(n2914 ,n2852 ,n2889);
    xnor g3467(n2724 ,n2656 ,n2685);
    nor g3468(n361 ,n921 ,n348);
    or g3469(n892 ,n767 ,n679);
    not g3470(n2368 ,n2367);
    nor g3471(n1191 ,n1016 ,n1170);
    or g3472(n635 ,n306 ,n631);
    not g3473(n40 ,n30[5]);
    nor g3474(n467 ,n274 ,n102);
    nor g3475(n1657 ,n1574 ,n1610);
    not g3476(n2372 ,n2371);
    nor g3477(n2913 ,n2853 ,n2888);
    or g3478(n3230 ,n3196 ,n3216);
    nor g3479(n3019 ,n3293 ,n3277);
    nor g3480(n999 ,n958 ,n992);
    or g3481(n607 ,n444 ,n359);
    not g3482(n1212 ,n1211);
    xnor g3483(n1713 ,n1670 ,n1601);
    nor g3484(n2682 ,n2574 ,n2635);
    nor g3485(n95 ,n80 ,n93);
    or g3486(n819 ,n719 ,n716);
    xnor g3487(n1439 ,n1402 ,n1340);
    nor g3488(n2513 ,n2340 ,n2406);
    nor g3489(n1019 ,n983 ,n1005);
    not g3490(n1343 ,n1342);
    xnor g3491(n2424 ,n2232 ,n2133);
    nor g3492(n2645 ,n2555 ,n2590);
    nor g3493(n2371 ,n2200 ,n2303);
    nor g3494(n2063 ,n1886 ,n1874);
    not g3495(n203 ,n21[4]);
    or g3496(n35 ,n30[3] ,n30[2]);
    dff g3497(.RN(n1), .SN(1'b1), .CK(n0), .D(n595), .Q(n10[8]));
    or g3498(n586 ,n415 ,n520);
    not g3499(n2550 ,n2549);
    nor g3500(n1542 ,n1522 ,n1534);
    xnor g3501(n2253 ,n1965 ,n2023);
    nor g3502(n1767 ,n1682 ,n1740);
    not g3503(n3114 ,n3287);
    dff g3504(.RN(n1), .SN(1'b1), .CK(n0), .D(n852), .Q(n27[1]));
    nor g3505(n763 ,n219 ,n664);
    nor g3506(n1069 ,n957 ,n1040);
    nor g3507(n2894 ,n2819 ,n2874);
    not g3508(n146 ,n2);
    nor g3509(n460 ,n266 ,n102);
    buf g3510(n9[23], 1'b0);
    or g3511(n3254 ,n3195 ,n3243);
    not g3512(n1220 ,n1219);
    nor g3513(n2089 ,n1879 ,n1870);
    nor g3514(n633 ,n333 ,n628);
    nor g3515(n2945 ,n2944 ,n2935);
    dff g3516(.RN(n1), .SN(1'b1), .CK(n0), .D(n537), .Q(n29[6]));
    not g3517(n2501 ,n2500);
    nor g3518(n513 ,n189 ,n346);
    nor g3519(n1625 ,n1575 ,n1597);
    buf g3520(n11[5], 1'b0);
    xnor g3521(n1294 ,n1182 ,n942);
    nor g3522(n1585 ,n1520 ,n1533);
    not g3523(n2799 ,n2798);
    xnor g3524(n2475 ,n2341 ,n2377);
    nor g3525(n935 ,n67 ,n68);
    xnor g3526(n1425 ,n1373 ,n1316);
    not g3527(n2855 ,n2854);
    or g3528(n593 ,n422 ,n502);
    not g3529(n1606 ,n1605);
    nor g3530(n2832 ,n2731 ,n2799);
    not g3531(n2182 ,n2181);
    nor g3532(n1393 ,n1281 ,n1358);
    dff g3533(.RN(n1), .SN(1'b1), .CK(n0), .D(n530), .Q(n30[4]));
    not g3534(n2415 ,n2414);
    xnor g3535(n2483 ,n2331 ,n2335);
    or g3536(n602 ,n432 ,n511);
    nor g3537(n3007 ,n3295 ,n3279);
    nor g3538(n2447 ,n2181 ,n2330);
    not g3539(n1405 ,n1404);
    nor g3540(n1572 ,n1522 ,n1535);
    or g3541(n53 ,n25[7] ,n52);
    nor g3542(n687 ,n114 ,n648);
    nor g3543(n1170 ,n1074 ,n1127);
    nor g3544(n1802 ,n1766 ,n1780);
    not g3545(n1861 ,n22[7]);
    buf g3546(n11[21], n10[5]);
    nor g3547(n475 ,n284 ,n104);
    nor g3548(n976 ,n966 ,n950);
    xnor g3549(n1242 ,n1026 ,n1157);
    nor g3550(n2826 ,n2783 ,n2810);
    not g3551(n2460 ,n2459);
    not g3552(n3068 ,n32[7]);
    or g3553(n821 ,n769 ,n817);
    nor g3554(n1695 ,n1662 ,n1660);
    nor g3555(n2364 ,n2283 ,n2277);
    nor g3556(n677 ,n106 ,n657);
    nor g3557(n2301 ,n1985 ,n2157);
    xnor g3558(n2884 ,n2845 ,n2817);
    buf g3559(n13[11], 1'b0);
    nor g3560(n345 ,n315 ,n301);
    xnor g3561(n1227 ,n1030 ,n1156);
    nor g3562(n2679 ,n2554 ,n2597);
    not g3563(n2868 ,n2867);
    xnor g3564(n2940 ,n2922 ,n2908);
    not g3565(n159 ,n31[2]);
    not g3566(n1414 ,n1413);
    nor g3567(n3272 ,n2147 ,n2217);
    nor g3568(n1640 ,n1539 ,n1588);
    or g3569(n568 ,n366 ,n475);
    nor g3570(n2849 ,n2742 ,n2835);
    not g3571(n1662 ,n1661);
    not g3572(n147 ,n29[6]);
    or g3573(n316 ,n5[21] ,n5[20]);
    nor g3574(n2069 ,n1864 ,n1873);
    dff g3575(.RN(n1), .SN(1'b1), .CK(n0), .D(n915), .Q(n9[5]));
    not g3576(n1732 ,n1731);
    buf g3577(n12[5], 1'b0);
    nor g3578(n2567 ,n2377 ,n2523);
    xnor g3579(n1179 ,n1016 ,n1095);
    buf g3580(n11[17], n10[1]);
    xnor g3581(n3317 ,n3033 ,n3047);
    nor g3582(n1365 ,n945 ,n1342);
    nor g3583(n463 ,n159 ,n102);
    nor g3584(n2643 ,n2390 ,n2602);
    nor g3585(n1494 ,n1450 ,n1493);
    nor g3586(n1230 ,n1090 ,n1178);
    nor g3587(n1076 ,n956 ,n1040);
    or g3588(n305 ,n26[2] ,n26[3]);
    or g3589(n587 ,n417 ,n497);
    or g3590(n534 ,n384 ,n468);
    nor g3591(n685 ,n109 ,n650);
    nor g3592(n933 ,n73 ,n74);
    nor g3593(n3012 ,n3290 ,n3274);
    nor g3594(n969 ,n20[7] ,n21[7]);
    nor g3595(n1977 ,n1865 ,n1876);
    nor g3596(n3042 ,n3029 ,n3041);
    dff g3597(.RN(n1), .SN(1'b1), .CK(n0), .D(n531), .Q(n29[10]));
    nor g3598(n2569 ,n2408 ,n2501);
    xnor g3599(n3279 ,n2917 ,n2928);
    not g3600(n948 ,n3310);
    xnor g3601(n3318 ,n3032 ,n3045);
    not g3602(n258 ,n25[1]);
    nor g3603(n766 ,n122 ,n664);
    not g3604(n2109 ,n2108);
    nor g3605(n2490 ,n2376 ,n2449);
endmodule
