module top(n0, n1, n2, n3, n4, n5, n6, n7);
    input n0, n1, n2, n3;
    input [15:0] n4;
    output [15:0] n5;
    output n6, n7;
    wire n0, n1, n2, n3;
    wire [15:0] n4;
    wire [15:0] n5;
    wire n6, n7;
    wire [15:0] n8;
    wire [15:0] n9;
    wire [15:0] n10;
    wire [15:0] n11;
    wire [15:0] n12;
    wire [15:0] n13;
    wire [15:0] n14;
    wire [15:0] n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [15:0] n18;
    wire [15:0] n19;
    wire [15:0] n20;
    wire [15:0] n21;
    wire [15:0] n22;
    wire [15:0] n23;
    wire [15:0] n24;
    wire [15:0] n25;
    wire [15:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire n31, n32, n33, n34, n35, n36, n37, n38;
    wire n39, n40, n41, n42, n43, n44, n45, n46;
    wire n47, n48, n49, n50, n51, n52, n53, n54;
    wire n55, n56, n57, n58, n59, n60, n61, n62;
    wire n63, n64, n65, n66, n67, n68, n69, n70;
    wire n71, n72, n73, n74, n75, n76, n77, n78;
    wire n79, n80, n81, n82, n83, n84, n85, n86;
    wire n87, n88, n89, n90, n91, n92, n93, n94;
    wire n95, n96, n97, n98, n99, n100, n101, n102;
    wire n103, n104, n105, n106, n107, n108, n109, n110;
    wire n111, n112, n113, n114, n115, n116, n117, n118;
    wire n119, n120, n121, n122, n123, n124, n125, n126;
    wire n127, n128, n129, n130, n131, n132, n133, n134;
    wire n135, n136, n137, n138, n139, n140, n141, n142;
    wire n143, n144, n145, n146, n147, n148, n149, n150;
    wire n151, n152, n153, n154, n155, n156, n157, n158;
    wire n159, n160, n161, n162, n163, n164, n165, n166;
    wire n167, n168, n169, n170, n171, n172, n173, n174;
    wire n175, n176, n177, n178, n179, n180, n181, n182;
    wire n183, n184, n185, n186, n187, n188, n189, n190;
    wire n191, n192, n193, n194, n195, n196, n197, n198;
    wire n199, n200, n201, n202, n203, n204, n205, n206;
    wire n207, n208, n209, n210, n211, n212, n213, n214;
    wire n215, n216, n217, n218, n219, n220, n221, n222;
    wire n223, n224, n225, n226, n227, n228, n229, n230;
    wire n231, n232, n233, n234, n235, n236, n237, n238;
    wire n239, n240, n241, n242, n243, n244, n245, n246;
    wire n247, n248, n249, n250, n251, n252, n253, n254;
    wire n255, n256, n257, n258, n259, n260, n261, n262;
    wire n263, n264, n265, n266, n267, n268, n269, n270;
    wire n271, n272, n273, n274, n275, n276, n277, n278;
    wire n279, n280, n281, n282, n283, n284, n285, n286;
    wire n287, n288, n289, n290, n291, n292, n293, n294;
    wire n295, n296, n297, n298, n299, n300, n301, n302;
    wire n303, n304, n305, n306, n307, n308, n309, n310;
    wire n311, n312, n313, n314, n315, n316, n317, n318;
    wire n319, n320, n321, n322, n323, n324, n325, n326;
    wire n327, n328, n329, n330, n331, n332, n333, n334;
    wire n335, n336, n337, n338, n339, n340, n341, n342;
    wire n343, n344, n345, n346, n347, n348, n349, n350;
    wire n351, n352, n353, n354, n355, n356, n357, n358;
    wire n359, n360, n361, n362, n363, n364, n365, n366;
    wire n367, n368, n369, n370, n371, n372, n373, n374;
    wire n375, n376, n377, n378, n379, n380, n381, n382;
    wire n383, n384, n385, n386, n387, n388, n389, n390;
    wire n391, n392, n393, n394, n395, n396, n397, n398;
    wire n399, n400, n401, n402, n403, n404, n405, n406;
    wire n407, n408, n409, n410, n411, n412, n413, n414;
    wire n415, n416, n417, n418, n419, n420, n421, n422;
    wire n423, n424, n425, n426, n427, n428, n429, n430;
    wire n431, n432, n433, n434, n435, n436, n437, n438;
    wire n439, n440, n441, n442, n443, n444, n445, n446;
    wire n447, n448, n449, n450, n451, n452, n453, n454;
    wire n455, n456, n457, n458, n459, n460, n461, n462;
    wire n463, n464, n465, n466, n467, n468, n469, n470;
    wire n471, n472, n473, n474, n475, n476, n477, n478;
    wire n479, n480, n481, n482, n483, n484, n485, n486;
    wire n487, n488, n489, n490, n491, n492, n493, n494;
    wire n495, n496, n497, n498, n499, n500, n501, n502;
    wire n503, n504, n505, n506, n507, n508, n509, n510;
    wire n511, n512, n513, n514, n515, n516, n517, n518;
    wire n519, n520, n521, n522, n523, n524, n525, n526;
    wire n527, n528, n529, n530, n531, n532, n533, n534;
    wire n535, n536, n537, n538, n539, n540, n541, n542;
    wire n543, n544, n545, n546, n547, n548, n549, n550;
    wire n551, n552, n553, n554, n555, n556, n557, n558;
    wire n559, n560, n561, n562, n563, n564, n565, n566;
    wire n567, n568, n569, n570, n571, n572, n573, n574;
    wire n575, n576, n577, n578, n579, n580, n581, n582;
    wire n583, n584, n585, n586, n587, n588, n589, n590;
    wire n591, n592, n593, n594, n595, n596, n597, n598;
    wire n599, n600, n601, n602, n603, n604, n605, n606;
    wire n607, n608, n609, n610, n611, n612, n613, n614;
    wire n615, n616, n617, n618, n619, n620, n621, n622;
    wire n623, n624, n625, n626, n627, n628, n629, n630;
    wire n631, n632, n633, n634, n635, n636, n637, n638;
    wire n639, n640, n641, n642, n643, n644, n645, n646;
    wire n647, n648, n649, n650, n651, n652, n653, n654;
    wire n655, n656, n657, n658, n659, n660, n661, n662;
    wire n663, n664, n665, n666, n667, n668, n669, n670;
    wire n671, n672, n673, n674, n675, n676, n677, n678;
    wire n679, n680, n681, n682, n683, n684, n685, n686;
    wire n687, n688, n689, n690, n691, n692, n693, n694;
    wire n695, n696, n697, n698, n699, n700, n701, n702;
    wire n703, n704, n705, n706, n707, n708, n709, n710;
    wire n711, n712, n713, n714, n715, n716, n717, n718;
    wire n719, n720, n721, n722, n723, n724, n725, n726;
    wire n727, n728, n729, n730, n731, n732, n733, n734;
    wire n735, n736, n737, n738, n739, n740, n741, n742;
    wire n743, n744, n745, n746, n747, n748, n749, n750;
    wire n751, n752, n753, n754, n755, n756, n757, n758;
    wire n759, n760, n761, n762, n763, n764, n765, n766;
    wire n767, n768, n769, n770, n771, n772, n773, n774;
    wire n775, n776, n777, n778, n779, n780, n781, n782;
    wire n783, n784, n785, n786, n787, n788, n789, n790;
    wire n791, n792, n793, n794, n795, n796, n797, n798;
    wire n799, n800, n801, n802, n803, n804, n805, n806;
    wire n807, n808, n809, n810, n811, n812, n813, n814;
    wire n815, n816, n817, n818, n819, n820, n821, n822;
    wire n823, n824, n825, n826, n827, n828, n829, n830;
    wire n831, n832, n833, n834, n835, n836, n837, n838;
    wire n839, n840, n841, n842, n843, n844, n845, n846;
    wire n847, n848, n849, n850, n851, n852, n853, n854;
    wire n855, n856, n857, n858, n859, n860, n861, n862;
    wire n863, n864, n865, n866, n867, n868, n869, n870;
    wire n871, n872, n873, n874, n875, n876, n877, n878;
    wire n879, n880, n881, n882, n883, n884, n885, n886;
    wire n887, n888, n889, n890, n891, n892, n893, n894;
    wire n895, n896, n897, n898, n899, n900, n901, n902;
    wire n903, n904, n905, n906, n907, n908, n909, n910;
    wire n911, n912, n913, n914, n915, n916, n917, n918;
    wire n919, n920, n921, n922, n923, n924, n925, n926;
    wire n927, n928, n929, n930, n931, n932, n933, n934;
    wire n935, n936, n937, n938, n939, n940, n941, n942;
    wire n943, n944, n945, n946, n947, n948, n949, n950;
    wire n951, n952, n953, n954, n955, n956, n957, n958;
    wire n959, n960, n961, n962, n963, n964, n965, n966;
    wire n967, n968, n969, n970, n971, n972, n973, n974;
    wire n975, n976, n977, n978, n979, n980, n981, n982;
    wire n983, n984, n985, n986, n987, n988, n989, n990;
    wire n991, n992, n993, n994, n995, n996, n997, n998;
    wire n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006;
    wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
    wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
    wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
    wire n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
    wire n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046;
    wire n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
    wire n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062;
    wire n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070;
    wire n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078;
    wire n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086;
    wire n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094;
    wire n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102;
    wire n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110;
    wire n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118;
    wire n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126;
    wire n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134;
    wire n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142;
    wire n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150;
    wire n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158;
    wire n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166;
    wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
    wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
    wire n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190;
    wire n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198;
    wire n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206;
    wire n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214;
    wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
    wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
    wire n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238;
    wire n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246;
    wire n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254;
    wire n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262;
    wire n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270;
    wire n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278;
    wire n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286;
    wire n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294;
    wire n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302;
    wire n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310;
    wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
    wire n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326;
    wire n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334;
    wire n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342;
    wire n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350;
    wire n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358;
    wire n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366;
    wire n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374;
    wire n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
    wire n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390;
    wire n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398;
    wire n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406;
    wire n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414;
    wire n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422;
    wire n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430;
    wire n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438;
    wire n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446;
    wire n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454;
    wire n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462;
    wire n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470;
    wire n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478;
    wire n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486;
    wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
    wire n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502;
    wire n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510;
    wire n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518;
    wire n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526;
    wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
    wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
    wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
    wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
    wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
    wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
    wire n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582;
    wire n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590;
    wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
    wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
    wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
    wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
    wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
    wire n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638;
    wire n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646;
    wire n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654;
    wire n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;
    wire n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670;
    wire n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678;
    wire n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686;
    wire n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694;
    wire n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702;
    wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
    wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
    wire n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726;
    wire n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734;
    wire n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742;
    wire n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750;
    wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758;
    wire n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766;
    wire n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774;
    wire n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782;
    wire n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790;
    wire n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798;
    wire n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806;
    wire n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814;
    wire n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822;
    wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    wire n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838;
    wire n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846;
    wire n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854;
    wire n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
    wire n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870;
    wire n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878;
    wire n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886;
    wire n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894;
    wire n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902;
    wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
    wire n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918;
    wire n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926;
    wire n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934;
    wire n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942;
    wire n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950;
    wire n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958;
    wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
    wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974;
    wire n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982;
    wire n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990;
    wire n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998;
    wire n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
    wire n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014;
    wire n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022;
    wire n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;
    wire n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038;
    wire n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046;
    wire n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
    wire n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062;
    wire n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070;
    wire n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078;
    wire n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086;
    wire n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094;
    wire n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
    wire n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110;
    wire n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118;
    wire n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126;
    wire n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134;
    wire n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142;
    wire n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150;
    wire n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158;
    wire n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166;
    wire n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174;
    wire n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182;
    wire n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190;
    wire n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198;
    wire n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
    wire n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214;
    wire n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222;
    wire n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230;
    wire n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238;
    wire n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246;
    wire n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
    wire n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262;
    wire n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270;
    wire n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278;
    wire n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286;
    wire n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294;
    wire n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
    wire n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310;
    wire n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318;
    wire n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326;
    wire n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334;
    wire n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342;
    wire n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
    wire n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358;
    wire n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366;
    wire n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374;
    wire n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382;
    wire n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390;
    wire n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398;
    wire n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
    wire n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414;
    wire n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422;
    wire n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430;
    wire n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
    wire n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446;
    wire n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
    wire n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462;
    wire n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470;
    wire n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478;
    wire n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486;
    wire n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494;
    wire n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
    wire n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510;
    wire n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;
    wire n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526;
    wire n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534;
    wire n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542;
    wire n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
    wire n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558;
    wire n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566;
    wire n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574;
    wire n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582;
    wire n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590;
    wire n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598;
    wire n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606;
    wire n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614;
    wire n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622;
    wire n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630;
    wire n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;
    wire n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646;
    wire n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
    wire n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662;
    wire n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670;
    wire n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678;
    wire n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686;
    wire n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694;
    wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
    wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
    wire n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718;
    wire n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726;
    wire n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734;
    wire n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742;
    wire n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
    wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
    wire n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766;
    wire n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774;
    wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
    wire n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790;
    wire n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
    wire n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806;
    wire n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814;
    wire n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822;
    wire n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830;
    wire n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838;
    wire n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846;
    wire n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854;
    wire n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862;
    wire n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870;
    wire n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878;
    wire n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886;
    wire n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894;
    wire n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
    wire n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910;
    wire n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918;
    wire n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926;
    wire n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934;
    wire n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942;
    wire n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950;
    wire n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958;
    wire n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966;
    wire n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974;
    wire n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982;
    wire n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990;
    wire n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
    wire n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006;
    wire n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014;
    wire n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022;
    wire n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030;
    wire n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038;
    wire n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046;
    wire n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054;
    wire n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062;
    wire n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070;
    wire n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078;
    wire n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
    wire n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
    wire n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102;
    wire n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110;
    wire n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118;
    wire n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126;
    wire n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134;
    wire n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142;
    wire n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150;
    wire n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158;
    wire n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166;
    wire n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174;
    wire n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182;
    wire n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190;
    wire n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198;
    wire n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206;
    wire n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214;
    wire n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222;
    wire n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230;
    wire n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238;
    wire n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246;
    wire n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254;
    wire n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262;
    wire n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270;
    wire n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278;
    wire n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286;
    wire n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294;
    wire n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302;
    wire n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310;
    wire n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318;
    wire n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326;
    wire n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334;
    wire n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342;
    wire n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350;
    wire n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358;
    wire n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366;
    wire n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374;
    wire n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382;
    wire n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390;
    wire n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398;
    wire n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406;
    wire n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414;
    wire n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422;
    wire n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430;
    wire n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438;
    wire n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446;
    wire n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454;
    wire n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462;
    wire n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470;
    wire n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478;
    wire n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486;
    wire n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494;
    wire n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502;
    wire n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510;
    wire n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518;
    wire n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526;
    wire n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534;
    wire n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542;
    wire n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550;
    wire n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558;
    wire n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566;
    wire n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574;
    wire n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582;
    wire n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590;
    wire n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598;
    wire n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606;
    wire n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614;
    wire n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622;
    wire n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630;
    wire n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638;
    wire n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646;
    wire n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654;
    wire n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662;
    wire n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670;
    wire n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678;
    wire n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686;
    wire n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694;
    wire n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702;
    wire n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710;
    wire n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718;
    wire n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726;
    wire n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734;
    wire n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742;
    wire n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750;
    wire n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758;
    wire n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766;
    wire n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774;
    wire n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782;
    wire n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790;
    wire n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798;
    wire n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806;
    wire n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814;
    wire n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822;
    wire n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830;
    wire n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838;
    wire n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846;
    wire n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854;
    wire n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862;
    wire n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870;
    wire n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878;
    wire n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886;
    wire n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894;
    wire n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902;
    wire n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910;
    wire n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918;
    wire n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926;
    wire n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934;
    wire n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942;
    wire n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950;
    wire n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958;
    wire n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966;
    wire n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974;
    wire n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982;
    wire n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990;
    wire n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998;
    wire n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006;
    wire n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014;
    wire n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022;
    wire n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030;
    wire n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038;
    wire n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046;
    wire n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054;
    wire n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062;
    wire n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070;
    wire n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078;
    wire n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086;
    wire n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094;
    wire n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102;
    wire n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110;
    wire n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118;
    wire n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126;
    wire n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134;
    wire n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142;
    wire n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150;
    wire n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158;
    wire n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166;
    wire n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174;
    wire n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182;
    wire n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190;
    wire n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198;
    wire n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206;
    wire n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214;
    wire n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222;
    wire n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230;
    wire n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238;
    wire n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246;
    wire n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254;
    wire n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262;
    wire n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270;
    wire n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278;
    wire n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286;
    wire n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294;
    wire n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302;
    wire n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310;
    wire n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318;
    wire n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326;
    wire n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334;
    wire n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342;
    wire n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350;
    wire n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358;
    wire n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366;
    wire n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374;
    wire n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382;
    wire n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390;
    wire n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398;
    wire n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406;
    wire n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414;
    wire n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422;
    wire n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430;
    wire n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438;
    wire n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446;
    wire n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454;
    wire n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462;
    wire n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470;
    wire n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478;
    wire n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486;
    wire n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494;
    wire n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502;
    wire n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510;
    wire n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518;
    wire n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526;
    wire n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534;
    wire n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542;
    wire n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550;
    wire n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558;
    wire n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566;
    wire n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574;
    wire n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582;
    wire n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590;
    wire n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598;
    wire n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606;
    wire n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614;
    wire n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622;
    wire n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630;
    wire n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638;
    wire n4639;
    dff g0(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2065), .Q(n6));
    dff g1(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2082), .Q(n7));
    dff g2(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n8[0]));
    dff g3(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n8[1]));
    dff g4(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1809), .Q(n8[2]));
    dff g5(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n8[3]));
    dff g6(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1761), .Q(n8[4]));
    dff g7(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1745), .Q(n8[5]));
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1742), .Q(n8[6]));
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n8[7]));
    dff g10(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n8[8]));
    dff g11(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1713), .Q(n8[9]));
    dff g12(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1670), .Q(n8[10]));
    dff g13(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n8[11]));
    dff g14(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n8[12]));
    dff g15(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n8[13]));
    dff g16(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n8[14]));
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n8[15]));
    dff g18(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n9[0]));
    dff g19(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n9[1]));
    dff g20(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n9[2]));
    dff g21(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n9[3]));
    dff g22(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1864), .Q(n9[4]));
    dff g23(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n9[5]));
    dff g24(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n9[6]));
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n9[7]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n9[8]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n9[9]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n9[10]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n9[11]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1801), .Q(n9[12]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n9[13]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n9[14]));
    dff g33(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n9[15]));
    dff g34(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n10[0]));
    dff g35(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n10[1]));
    dff g36(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1760), .Q(n10[2]));
    dff g37(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n10[3]));
    dff g38(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n10[4]));
    dff g39(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n10[5]));
    dff g40(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n10[6]));
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1744), .Q(n10[7]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1740), .Q(n10[8]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1734), .Q(n10[9]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1733), .Q(n10[10]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1730), .Q(n10[11]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1727), .Q(n10[12]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1724), .Q(n10[13]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1722), .Q(n10[14]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1716), .Q(n10[15]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1712), .Q(n11[0]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1703), .Q(n11[1]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1695), .Q(n11[2]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1692), .Q(n11[3]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1681), .Q(n11[4]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n11[5]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1667), .Q(n11[6]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1656), .Q(n11[7]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1650), .Q(n11[8]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n11[9]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n11[10]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n11[11]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n11[12]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n11[13]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n11[14]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n11[15]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n12[0]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n12[1]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n12[2]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n12[3]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1941), .Q(n12[4]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n12[5]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n12[6]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n12[7]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n12[8]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n12[9]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n12[10]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n12[11]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n12[12]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n12[13]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n12[14]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n12[15]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n13[0]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n13[1]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n13[2]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1852), .Q(n13[3]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n13[4]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n13[5]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n13[6]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1837), .Q(n13[7]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1834), .Q(n13[8]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n13[9]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n13[10]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1823), .Q(n13[11]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n13[12]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n13[13]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1811), .Q(n13[14]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1807), .Q(n13[15]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n14[0]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n14[1]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n14[2]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n14[3]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n14[4]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n14[5]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n14[6]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n14[7]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n14[8]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n14[9]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n14[10]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n14[11]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1762), .Q(n14[12]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1759), .Q(n14[13]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1758), .Q(n14[14]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n14[15]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n15[0]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n15[1]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1752), .Q(n15[2]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n15[3]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n15[4]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1747), .Q(n15[5]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1746), .Q(n15[6]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1743), .Q(n15[7]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1741), .Q(n15[8]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1739), .Q(n15[9]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1738), .Q(n15[10]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1737), .Q(n15[11]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1735), .Q(n15[12]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1732), .Q(n15[13]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1731), .Q(n15[14]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1729), .Q(n15[15]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1728), .Q(n16[0]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1726), .Q(n16[1]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1725), .Q(n16[2]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1723), .Q(n16[3]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1721), .Q(n16[4]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1720), .Q(n16[5]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n16[6]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1714), .Q(n16[7]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1710), .Q(n16[8]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1708), .Q(n16[9]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1705), .Q(n16[10]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1702), .Q(n16[11]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1699), .Q(n16[12]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1694), .Q(n16[13]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1691), .Q(n16[14]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1687), .Q(n16[15]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1684), .Q(n17[0]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1679), .Q(n17[1]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n17[2]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1671), .Q(n17[3]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1666), .Q(n17[4]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1663), .Q(n17[5]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n17[6]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1655), .Q(n17[7]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n17[8]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n17[9]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1644), .Q(n17[10]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n17[11]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1637), .Q(n17[12]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n17[13]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n17[14]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1626), .Q(n17[15]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1685), .Q(n18[0]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n18[1]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n18[2]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n18[3]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n18[4]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n18[5]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n18[6]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n18[7]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n18[8]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n18[9]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n18[10]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n18[11]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n18[12]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n18[13]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n18[14]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n18[15]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n19[0]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1940), .Q(n19[1]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1937), .Q(n19[2]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n19[3]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1928), .Q(n19[4]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n19[5]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1921), .Q(n19[6]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n19[7]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n19[8]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n19[9]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n19[10]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n19[11]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n19[12]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n19[13]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n19[14]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n19[15]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n20[0]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n20[1]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n20[2]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n20[3]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n20[4]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n20[5]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n20[6]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n20[7]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n20[8]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n20[9]));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n20[10]));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n20[11]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n20[12]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n20[13]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n20[14]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1851), .Q(n20[15]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n21[0]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n21[1]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n21[2]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n21[3]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n21[4]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n21[5]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n21[6]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n21[7]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1835), .Q(n21[8]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n21[9]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n21[10]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n21[11]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n21[12]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1825), .Q(n21[13]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n21[14]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n21[15]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n22[0]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n22[1]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n22[2]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n22[3]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1717), .Q(n22[4]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n22[5]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1808), .Q(n22[6]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n22[7]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n22[8]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n22[9]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n22[10]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n22[11]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n22[12]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n22[13]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n22[14]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n22[15]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n23[0]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n23[1]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n23[2]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n23[3]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n23[4]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n23[5]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n23[6]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n23[7]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n23[8]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n23[9]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n23[10]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n23[11]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n23[12]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1767), .Q(n23[13]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n23[14]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n23[15]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n738), .Q(n24[0]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n755), .Q(n24[1]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n739), .Q(n24[2]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n737), .Q(n24[3]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n676), .Q(n24[4]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n675), .Q(n24[5]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n674), .Q(n24[6]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n679), .Q(n24[7]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n736), .Q(n25[0]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n735), .Q(n25[1]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n734), .Q(n25[2]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n733), .Q(n25[3]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n669), .Q(n25[4]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n668), .Q(n25[5]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n667), .Q(n25[6]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n666), .Q(n25[7]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n770), .Q(n26[0]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n763), .Q(n26[1]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n852), .Q(n26[2]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n851), .Q(n26[3]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n796), .Q(n26[4]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n797), .Q(n26[5]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n799), .Q(n26[6]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n798), .Q(n26[7]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n761), .Q(n26[8]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n771), .Q(n26[9]));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n760), .Q(n26[10]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n754), .Q(n26[11]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n762), .Q(n26[12]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n764), .Q(n26[13]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n765), .Q(n26[14]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n759), .Q(n26[15]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2218), .Q(n5[0]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2205), .Q(n5[1]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2200), .Q(n5[2]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2213), .Q(n5[3]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2203), .Q(n5[4]));
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2214), .Q(n5[5]));
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2217), .Q(n5[6]));
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2208), .Q(n5[7]));
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2211), .Q(n5[8]));
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2210), .Q(n5[9]));
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2216), .Q(n5[10]));
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2209), .Q(n5[11]));
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2215), .Q(n5[12]));
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2212), .Q(n5[13]));
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2206), .Q(n5[14]));
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2207), .Q(n5[15]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n613), .Q(n27[0]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n614), .Q(n27[1]));
    dff g308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n603), .Q(n27[2]));
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n601), .Q(n27[3]));
    dff g310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n608), .Q(n27[4]));
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n612), .Q(n27[5]));
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n609), .Q(n27[6]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n611), .Q(n27[7]));
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n600), .Q(n28[0]));
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n595), .Q(n28[1]));
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n593), .Q(n28[2]));
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n596), .Q(n28[3]));
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n617), .Q(n28[4]));
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n621), .Q(n28[5]));
    dff g320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n615), .Q(n28[6]));
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n618), .Q(n28[7]));
    or g322(n2218 ,n2145 ,n2199);
    or g323(n2217 ,n2154 ,n2202);
    or g324(n2216 ,n2150 ,n2201);
    or g325(n2215 ,n2148 ,n2204);
    or g326(n2214 ,n2140 ,n2197);
    or g327(n2213 ,n2142 ,n2198);
    or g328(n2212 ,n2181 ,n2176);
    or g329(n2211 ,n2183 ,n2179);
    or g330(n2210 ,n2182 ,n2178);
    or g331(n2209 ,n2192 ,n2177);
    or g332(n2208 ,n2188 ,n2180);
    or g333(n2207 ,n2194 ,n2174);
    or g334(n2206 ,n2195 ,n2175);
    or g335(n2205 ,n2184 ,n2173);
    or g336(n2204 ,n778 ,n2196);
    or g337(n2203 ,n2186 ,n2171);
    or g338(n2202 ,n782 ,n2189);
    or g339(n2201 ,n787 ,n2193);
    or g340(n2200 ,n2191 ,n2172);
    or g341(n2199 ,n790 ,n2187);
    or g342(n2198 ,n793 ,n2190);
    or g343(n2197 ,n792 ,n2185);
    nor g344(n2196 ,n144 ,n2161);
    nor g345(n2195 ,n146 ,n2159);
    nor g346(n2194 ,n143 ,n2158);
    nor g347(n2193 ,n142 ,n2163);
    nor g348(n2192 ,n139 ,n2162);
    nor g349(n2191 ,n137 ,n2170);
    nor g350(n2190 ,n138 ,n2139);
    nor g351(n2189 ,n134 ,n2167);
    nor g352(n2188 ,n136 ,n2166);
    nor g353(n2187 ,n132 ,n2157);
    nor g354(n2186 ,n135 ,n2153);
    nor g355(n2185 ,n133 ,n2152);
    nor g356(n2184 ,n131 ,n2156);
    nor g357(n2183 ,n29[8] ,n2165);
    nor g358(n2182 ,n29[9] ,n2164);
    nor g359(n2181 ,n29[13] ,n2160);
    or g360(n2180 ,n786 ,n2151);
    or g361(n2179 ,n783 ,n2169);
    or g362(n2178 ,n788 ,n2168);
    or g363(n2177 ,n780 ,n2149);
    or g364(n2176 ,n784 ,n2155);
    or g365(n2175 ,n789 ,n2147);
    or g366(n2174 ,n781 ,n2146);
    or g367(n2173 ,n791 ,n2144);
    or g368(n2172 ,n779 ,n2143);
    or g369(n2171 ,n785 ,n2141);
    or g370(n2170 ,n746 ,n2116);
    nor g371(n2169 ,n141 ,n2135);
    nor g372(n2168 ,n140 ,n2133);
    or g373(n2167 ,n746 ,n2108);
    or g374(n2166 ,n746 ,n2130);
    or g375(n2165 ,n746 ,n2136);
    or g376(n2164 ,n746 ,n2134);
    or g377(n2163 ,n746 ,n2132);
    or g378(n2162 ,n746 ,n2138);
    or g379(n2161 ,n746 ,n2128);
    or g380(n2160 ,n746 ,n2126);
    or g381(n2159 ,n746 ,n2124);
    or g382(n2158 ,n746 ,n2114);
    or g383(n2157 ,n746 ,n2120);
    or g384(n2156 ,n746 ,n2118);
    nor g385(n2155 ,n145 ,n2125);
    nor g386(n2154 ,n29[6] ,n2107);
    or g387(n2153 ,n746 ,n2112);
    or g388(n2152 ,n746 ,n2110);
    nor g389(n2151 ,n29[7] ,n2129);
    nor g390(n2150 ,n29[10] ,n2131);
    nor g391(n2149 ,n29[11] ,n2137);
    nor g392(n2148 ,n29[12] ,n2127);
    nor g393(n2147 ,n29[14] ,n2123);
    nor g394(n2146 ,n29[15] ,n2113);
    nor g395(n2145 ,n29[0] ,n2119);
    nor g396(n2144 ,n29[1] ,n2117);
    nor g397(n2143 ,n29[2] ,n2115);
    nor g398(n2142 ,n29[3] ,n2121);
    nor g399(n2141 ,n29[4] ,n2111);
    nor g400(n2140 ,n29[5] ,n2109);
    or g401(n2139 ,n746 ,n2122);
    not g402(n2138 ,n2137);
    not g403(n2136 ,n2135);
    not g404(n2134 ,n2133);
    not g405(n2132 ,n2131);
    not g406(n2130 ,n2129);
    not g407(n2128 ,n2127);
    not g408(n2126 ,n2125);
    not g409(n2124 ,n2123);
    nor g410(n2137 ,n2042 ,n2101);
    nor g411(n2135 ,n2051 ,n2104);
    nor g412(n2133 ,n2048 ,n2103);
    nor g413(n2131 ,n2045 ,n2106);
    nor g414(n2129 ,n2054 ,n2105);
    nor g415(n2127 ,n2039 ,n2100);
    nor g416(n2125 ,n2036 ,n2102);
    nor g417(n2123 ,n2033 ,n2091);
    not g418(n2122 ,n2121);
    not g419(n2120 ,n2119);
    not g420(n2118 ,n2117);
    not g421(n2116 ,n2115);
    not g422(n2114 ,n2113);
    not g423(n2112 ,n2111);
    not g424(n2110 ,n2109);
    not g425(n2108 ,n2107);
    nor g426(n2121 ,n2018 ,n2094);
    nor g427(n2119 ,n2027 ,n2097);
    nor g428(n2117 ,n2024 ,n2096);
    nor g429(n2115 ,n2021 ,n2095);
    nor g430(n2113 ,n2030 ,n2098);
    nor g431(n2111 ,n2015 ,n2093);
    nor g432(n2109 ,n2012 ,n2092);
    nor g433(n2107 ,n2009 ,n2099);
    or g434(n2106 ,n1950 ,n2086);
    or g435(n2105 ,n1992 ,n2089);
    or g436(n2104 ,n1978 ,n2088);
    or g437(n2103 ,n1964 ,n2087);
    or g438(n2102 ,n1906 ,n2083);
    or g439(n2101 ,n1936 ,n2085);
    or g440(n2100 ,n1922 ,n2084);
    or g441(n2099 ,n1623 ,n2075);
    or g442(n2098 ,n1700 ,n2074);
    or g443(n2097 ,n1711 ,n2081);
    or g444(n2096 ,n1842 ,n2080);
    or g445(n2095 ,n1680 ,n2079);
    or g446(n2094 ,n1665 ,n2078);
    or g447(n2093 ,n1651 ,n2077);
    or g448(n2092 ,n1638 ,n2076);
    or g449(n2091 ,n1893 ,n2090);
    or g450(n2090 ,n1891 ,n2066);
    or g451(n2089 ,n1990 ,n2069);
    or g452(n2088 ,n1977 ,n2072);
    or g453(n2087 ,n1962 ,n2071);
    or g454(n2086 ,n1948 ,n2070);
    or g455(n2085 ,n1935 ,n2073);
    or g456(n2084 ,n1919 ,n2068);
    or g457(n2083 ,n1904 ,n2067);
    xnor g458(n2082 ,n131 ,n2008);
    or g459(n2081 ,n1709 ,n2064);
    or g460(n2080 ,n1693 ,n2063);
    or g461(n2079 ,n1678 ,n2062);
    or g462(n2078 ,n1664 ,n2061);
    or g463(n2077 ,n1649 ,n2060);
    or g464(n2076 ,n1636 ,n2059);
    or g465(n2075 ,n1622 ,n2058);
    or g466(n2074 ,n1877 ,n2057);
    or g467(n2073 ,n2041 ,n2040);
    or g468(n2072 ,n2050 ,n2049);
    or g469(n2071 ,n2047 ,n2046);
    or g470(n2070 ,n2044 ,n2043);
    or g471(n2069 ,n2053 ,n2052);
    or g472(n2068 ,n2038 ,n2037);
    or g473(n2067 ,n2035 ,n2034);
    or g474(n2066 ,n2032 ,n2031);
    xnor g475(n2065 ,n29[0] ,n1815);
    or g476(n2064 ,n2026 ,n2025);
    or g477(n2063 ,n2023 ,n2022);
    or g478(n2062 ,n2020 ,n2019);
    or g479(n2061 ,n2017 ,n2016);
    or g480(n2060 ,n2014 ,n2013);
    or g481(n2059 ,n2011 ,n2010);
    or g482(n2058 ,n2055 ,n2056);
    or g483(n2057 ,n2029 ,n2028);
    or g484(n2056 ,n2001 ,n2000);
    or g485(n2055 ,n2004 ,n2002);
    or g486(n2054 ,n1995 ,n1994);
    or g487(n2053 ,n1988 ,n1987);
    or g488(n2052 ,n1986 ,n1985);
    or g489(n2051 ,n1981 ,n1980);
    or g490(n2050 ,n1975 ,n1974);
    or g491(n2049 ,n1972 ,n1970);
    or g492(n2048 ,n1967 ,n1966);
    or g493(n2047 ,n1960 ,n1959);
    or g494(n2046 ,n1958 ,n1957);
    or g495(n2045 ,n1953 ,n1952);
    or g496(n2044 ,n1946 ,n1945);
    or g497(n2043 ,n1942 ,n1943);
    or g498(n2042 ,n1939 ,n1938);
    or g499(n2041 ,n1931 ,n1932);
    or g500(n2040 ,n1930 ,n1929);
    or g501(n2039 ,n1924 ,n1923);
    or g502(n2038 ,n1917 ,n1915);
    or g503(n2037 ,n1914 ,n1913);
    or g504(n2036 ,n1909 ,n1908);
    or g505(n2035 ,n1902 ,n1901);
    or g506(n2034 ,n1900 ,n1899);
    or g507(n2033 ,n1883 ,n1895);
    or g508(n2032 ,n1890 ,n1888);
    or g509(n2031 ,n1886 ,n1885);
    or g510(n2030 ,n1881 ,n1880);
    or g511(n2029 ,n1876 ,n1875);
    or g512(n2028 ,n1696 ,n1873);
    or g513(n2027 ,n1718 ,n1715);
    or g514(n2026 ,n1707 ,n1706);
    or g515(n2025 ,n1704 ,n1701);
    or g516(n2024 ,n1698 ,n1697);
    or g517(n2023 ,n1690 ,n1689);
    or g518(n2022 ,n1688 ,n1686);
    or g519(n2021 ,n1683 ,n1682);
    or g520(n2020 ,n1677 ,n1676);
    or g521(n2019 ,n1673 ,n1672);
    or g522(n2018 ,n1669 ,n1668);
    or g523(n2017 ,n1662 ,n1661);
    or g524(n2016 ,n1659 ,n1657);
    or g525(n2015 ,n1654 ,n1653);
    or g526(n2014 ,n1647 ,n1646);
    or g527(n2013 ,n1645 ,n1643);
    or g528(n2012 ,n1640 ,n1639);
    or g529(n2011 ,n1635 ,n2005);
    or g530(n2010 ,n1631 ,n1630);
    or g531(n2009 ,n1625 ,n1624);
    nor g532(n2008 ,n850 ,n1816);
    or g533(n2007 ,n1370 ,n1098);
    or g534(n2006 ,n1284 ,n988);
    or g535(n2005 ,n1501 ,n1420);
    or g536(n2004 ,n1617 ,n1616);
    or g537(n2003 ,n1174 ,n959);
    or g538(n2002 ,n1615 ,n1614);
    or g539(n2001 ,n1613 ,n1612);
    or g540(n2000 ,n1610 ,n1611);
    or g541(n1999 ,n1406 ,n1095);
    or g542(n1998 ,n1408 ,n1088);
    or g543(n1997 ,n1159 ,n1104);
    or g544(n1996 ,n1402 ,n1061);
    or g545(n1995 ,n1606 ,n1605);
    or g546(n1994 ,n1604 ,n1433);
    or g547(n1993 ,n1162 ,n1105);
    or g548(n1992 ,n1602 ,n1603);
    or g549(n1991 ,n1357 ,n876);
    or g550(n1990 ,n1601 ,n1435);
    or g551(n1989 ,n1169 ,n886);
    or g552(n1988 ,n1600 ,n1599);
    or g553(n1987 ,n1596 ,n1597);
    or g554(n1986 ,n1594 ,n1595);
    or g555(n1985 ,n1470 ,n1593);
    or g556(n1984 ,n1401 ,n877);
    or g557(n1983 ,n1398 ,n895);
    or g558(n1982 ,n1399 ,n1101);
    or g559(n1981 ,n1155 ,n1154);
    or g560(n1980 ,n1153 ,n1109);
    or g561(n1979 ,n1397 ,n1100);
    or g562(n1978 ,n1123 ,n1118);
    or g563(n1977 ,n1152 ,n1110);
    or g564(n1976 ,n1396 ,n905);
    or g565(n1975 ,n1112 ,n1151);
    or g566(n1974 ,n1150 ,n1111);
    or g567(n1973 ,n1395 ,n937);
    or g568(n1972 ,n1149 ,n1115);
    or g569(n1971 ,n1394 ,n1097);
    or g570(n1970 ,n1113 ,n1148);
    or g571(n1969 ,n1388 ,n983);
    or g572(n1968 ,n1393 ,n1094);
    or g573(n1967 ,n1114 ,n1117);
    or g574(n1966 ,n1147 ,n1127);
    or g575(n1965 ,n1239 ,n947);
    or g576(n1964 ,n1146 ,n1119);
    or g577(n1963 ,n1225 ,n1092);
    or g578(n1962 ,n1144 ,n1145);
    or g579(n1961 ,n1618 ,n874);
    or g580(n1960 ,n1120 ,n1121);
    or g581(n1959 ,n1142 ,n1122);
    or g582(n1958 ,n1141 ,n1125);
    or g583(n1957 ,n1124 ,n1140);
    or g584(n1956 ,n1382 ,n1036);
    or g585(n1955 ,n1387 ,n1089);
    or g586(n1954 ,n1257 ,n971);
    or g587(n1953 ,n1584 ,n1503);
    or g588(n1952 ,n1583 ,n1582);
    or g589(n1951 ,n1386 ,n853);
    or g590(n1950 ,n1580 ,n1579);
    or g591(n1949 ,n1280 ,n990);
    or g592(n1948 ,n1578 ,n1504);
    or g593(n1947 ,n1270 ,n1090);
    or g594(n1946 ,n1577 ,n1576);
    or g595(n1945 ,n1575 ,n1505);
    or g596(n1944 ,n1383 ,n1084);
    or g597(n1943 ,n1570 ,n1571);
    or g598(n1942 ,n1573 ,n1572);
    or g599(n1941 ,n1296 ,n1004);
    or g600(n1940 ,n1381 ,n1001);
    or g601(n1939 ,n1568 ,n1567);
    or g602(n1938 ,n1566 ,n1508);
    or g603(n1937 ,n1310 ,n1083);
    or g604(n1936 ,n1564 ,n1565);
    or g605(n1935 ,n1563 ,n1507);
    or g606(n1934 ,n1323 ,n1027);
    or g607(n1933 ,n1380 ,n1035);
    or g608(n1932 ,n1559 ,n1560);
    or g609(n1931 ,n1562 ,n1561);
    or g610(n1930 ,n1557 ,n1558);
    or g611(n1929 ,n1509 ,n1556);
    or g612(n1928 ,n1328 ,n1038);
    or g613(n1927 ,n1378 ,n1078);
    or g614(n1926 ,n1346 ,n1058);
    or g615(n1925 ,n1373 ,n865);
    or g616(n1924 ,n1554 ,n1512);
    or g617(n1923 ,n1553 ,n1552);
    or g618(n1922 ,n1551 ,n1527);
    or g619(n1921 ,n1355 ,n1059);
    or g620(n1920 ,n1371 ,n1076);
    or g621(n1919 ,n1549 ,n1548);
    or g622(n1918 ,n1403 ,n1075);
    or g623(n1917 ,n1533 ,n1531);
    or g624(n1916 ,n1374 ,n1018);
    or g625(n1915 ,n1547 ,n1546);
    or g626(n1914 ,n1545 ,n1555);
    or g627(n1913 ,n1543 ,n1544);
    or g628(n1912 ,n1372 ,n1074);
    or g629(n1911 ,n1285 ,n987);
    or g630(n1910 ,n1317 ,n1086);
    or g631(n1909 ,n1126 ,n1139);
    or g632(n1908 ,n1136 ,n1137);
    or g633(n1907 ,n1367 ,n1068);
    or g634(n1906 ,n1135 ,n1143);
    or g635(n1905 ,n1390 ,n1071);
    or g636(n1904 ,n1133 ,n1134);
    or g637(n1903 ,n1368 ,n1069);
    or g638(n1902 ,n1132 ,n1156);
    or g639(n1901 ,n1130 ,n1131);
    or g640(n1900 ,n1129 ,n1128);
    or g641(n1899 ,n1116 ,n1138);
    or g642(n1898 ,n1160 ,n854);
    or g643(n1897 ,n1379 ,n1070);
    or g644(n1896 ,n1263 ,n864);
    or g645(n1895 ,n1538 ,n1607);
    or g646(n1894 ,n1404 ,n927);
    or g647(n1893 ,n1536 ,n1430);
    or g648(n1892 ,n1180 ,n1065);
    or g649(n1891 ,n1535 ,n1591);
    or g650(n1890 ,n1526 ,n1569);
    or g651(n1889 ,n1358 ,n1063);
    or g652(n1888 ,n1540 ,n1585);
    or g653(n1887 ,n1334 ,n1080);
    or g654(n1886 ,n1530 ,n1438);
    or g655(n1885 ,n1529 ,n1528);
    or g656(n1884 ,n1360 ,n967);
    or g657(n1883 ,n1608 ,n1539);
    or g658(n1882 ,n1391 ,n1020);
    or g659(n1881 ,n1525 ,n1485);
    or g660(n1880 ,n1523 ,n1422);
    or g661(n1879 ,n1361 ,n1005);
    or g662(n1878 ,n1365 ,n1085);
    or g663(n1877 ,n1520 ,n1590);
    or g664(n1876 ,n1519 ,n1459);
    or g665(n1875 ,n1518 ,n1426);
    or g666(n1874 ,n1277 ,n913);
    or g667(n1873 ,n1521 ,n1515);
    or g668(n1872 ,n1356 ,n1102);
    or g669(n1871 ,n1353 ,n1056);
    or g670(n1870 ,n1342 ,n1052);
    or g671(n1869 ,n1352 ,n1053);
    or g672(n1868 ,n1351 ,n1054);
    or g673(n1867 ,n1349 ,n1051);
    or g674(n1866 ,n1348 ,n1048);
    or g675(n1865 ,n1347 ,n1049);
    or g676(n1864 ,n1340 ,n1042);
    or g677(n1863 ,n1345 ,n1046);
    or g678(n1862 ,n1344 ,n1043);
    or g679(n1861 ,n1343 ,n1045);
    or g680(n1860 ,n1341 ,n1044);
    or g681(n1859 ,n1338 ,n1041);
    or g682(n1858 ,n1339 ,n1040);
    or g683(n1857 ,n1337 ,n1037);
    or g684(n1856 ,n1332 ,n1028);
    or g685(n1855 ,n1335 ,n1032);
    or g686(n1854 ,n1336 ,n1034);
    or g687(n1853 ,n1333 ,n1033);
    or g688(n1852 ,n1330 ,n1030);
    or g689(n1851 ,n1331 ,n1031);
    or g690(n1850 ,n1327 ,n1029);
    or g691(n1849 ,n1325 ,n1025);
    or g692(n1848 ,n1326 ,n1026);
    or g693(n1847 ,n1321 ,n1016);
    or g694(n1846 ,n1322 ,n1023);
    or g695(n1845 ,n1318 ,n1021);
    or g696(n1844 ,n1316 ,n1017);
    or g697(n1843 ,n1319 ,n1022);
    or g698(n1842 ,n1480 ,n1481);
    or g699(n1841 ,n1314 ,n1012);
    or g700(n1840 ,n1315 ,n1014);
    or g701(n1839 ,n1312 ,n1011);
    or g702(n1838 ,n1306 ,n1007);
    or g703(n1837 ,n1309 ,n1009);
    or g704(n1836 ,n1308 ,n1008);
    or g705(n1835 ,n1307 ,n1006);
    or g706(n1834 ,n1303 ,n1002);
    or g707(n1833 ,n1304 ,n1003);
    or g708(n1832 ,n1302 ,n1013);
    or g709(n1831 ,n1301 ,n999);
    or g710(n1830 ,n1300 ,n1010);
    or g711(n1829 ,n1299 ,n998);
    or g712(n1828 ,n1305 ,n1000);
    or g713(n1827 ,n1295 ,n1047);
    or g714(n1826 ,n1297 ,n996);
    or g715(n1825 ,n1298 ,n997);
    or g716(n1824 ,n1294 ,n1024);
    or g717(n1823 ,n1293 ,n993);
    or g718(n1822 ,n1292 ,n995);
    or g719(n1821 ,n1287 ,n1060);
    or g720(n1820 ,n1290 ,n994);
    or g721(n1819 ,n1289 ,n991);
    or g722(n1818 ,n1288 ,n992);
    or g723(n1817 ,n1286 ,n989);
    not g724(n1816 ,n1815);
    or g725(n1814 ,n1183 ,n887);
    or g726(n1813 ,n1320 ,n975);
    or g727(n1812 ,n1274 ,n979);
    or g728(n1811 ,n1282 ,n984);
    or g729(n1810 ,n1281 ,n985);
    or g730(n1809 ,n1273 ,n954);
    or g731(n1808 ,n1279 ,n982);
    or g732(n1807 ,n1276 ,n980);
    or g733(n1806 ,n1375 ,n981);
    or g734(n1805 ,n1275 ,n1081);
    or g735(n1804 ,n1272 ,n973);
    or g736(n1803 ,n1271 ,n976);
    or g737(n1802 ,n1268 ,n974);
    or g738(n1801 ,n1269 ,n972);
    or g739(n1800 ,n1267 ,n1091);
    or g740(n1799 ,n1266 ,n969);
    or g741(n1798 ,n1264 ,n970);
    or g742(n1797 ,n1259 ,n964);
    or g743(n1796 ,n1261 ,n857);
    or g744(n1795 ,n1262 ,n968);
    or g745(n1794 ,n1260 ,n966);
    or g746(n1793 ,n1258 ,n965);
    or g747(n1792 ,n1256 ,n963);
    or g748(n1791 ,n1255 ,n962);
    or g749(n1790 ,n1247 ,n934);
    or g750(n1789 ,n1253 ,n955);
    or g751(n1788 ,n1254 ,n858);
    or g752(n1787 ,n1252 ,n960);
    or g753(n1786 ,n1251 ,n961);
    or g754(n1785 ,n1242 ,n950);
    or g755(n1784 ,n1250 ,n958);
    or g756(n1783 ,n1249 ,n957);
    or g757(n1782 ,n1248 ,n956);
    or g758(n1781 ,n1244 ,n951);
    or g759(n1780 ,n1246 ,n953);
    or g760(n1779 ,n1245 ,n952);
    or g761(n1778 ,n1243 ,n867);
    or g762(n1777 ,n1241 ,n949);
    or g763(n1776 ,n1240 ,n871);
    or g764(n1775 ,n1621 ,n945);
    or g765(n1774 ,n1620 ,n948);
    or g766(n1773 ,n1238 ,n946);
    or g767(n1772 ,n1237 ,n878);
    or g768(n1771 ,n1236 ,n943);
    or g769(n1770 ,n1235 ,n944);
    or g770(n1769 ,n1619 ,n942);
    or g771(n1768 ,n1232 ,n940);
    or g772(n1767 ,n1234 ,n880);
    or g773(n1766 ,n1233 ,n941);
    or g774(n1765 ,n1231 ,n939);
    or g775(n1764 ,n1229 ,n938);
    or g776(n1763 ,n1230 ,n936);
    or g777(n1762 ,n1228 ,n935);
    or g778(n1761 ,n1227 ,n925);
    or g779(n1760 ,n1224 ,n931);
    or g780(n1759 ,n1226 ,n933);
    or g781(n1758 ,n1222 ,n932);
    or g782(n1757 ,n1220 ,n930);
    or g783(n1756 ,n1221 ,n928);
    or g784(n1755 ,n1219 ,n929);
    or g785(n1754 ,n1218 ,n924);
    or g786(n1753 ,n1217 ,n926);
    or g787(n1752 ,n1216 ,n923);
    or g788(n1751 ,n1215 ,n922);
    or g789(n1750 ,n1214 ,n921);
    or g790(n1749 ,n1213 ,n920);
    or g791(n1748 ,n1211 ,n918);
    or g792(n1747 ,n1212 ,n919);
    or g793(n1746 ,n1210 ,n917);
    or g794(n1745 ,n1223 ,n910);
    or g795(n1744 ,n1209 ,n914);
    or g796(n1743 ,n1208 ,n916);
    or g797(n1742 ,n1204 ,n899);
    or g798(n1741 ,n1207 ,n915);
    or g799(n1740 ,n1205 ,n911);
    or g800(n1739 ,n1206 ,n912);
    or g801(n1738 ,n1203 ,n909);
    or g802(n1737 ,n1201 ,n907);
    or g803(n1736 ,n1196 ,n888);
    or g804(n1735 ,n1200 ,n906);
    or g805(n1734 ,n1202 ,n908);
    or g806(n1733 ,n1198 ,n903);
    or g807(n1732 ,n1199 ,n904);
    or g808(n1731 ,n1197 ,n902);
    or g809(n1730 ,n1195 ,n901);
    or g810(n1729 ,n1194 ,n900);
    or g811(n1728 ,n1193 ,n898);
    or g812(n1727 ,n1192 ,n897);
    or g813(n1726 ,n1191 ,n896);
    or g814(n1725 ,n1190 ,n894);
    or g815(n1724 ,n1189 ,n893);
    or g816(n1723 ,n1188 ,n892);
    or g817(n1722 ,n1186 ,n889);
    or g818(n1721 ,n1187 ,n891);
    or g819(n1720 ,n1185 ,n890);
    or g820(n1719 ,n1184 ,n879);
    or g821(n1718 ,n1500 ,n1499);
    or g822(n1717 ,n1283 ,n986);
    or g823(n1716 ,n1265 ,n859);
    or g824(n1715 ,n1498 ,n1502);
    or g825(n1714 ,n1182 ,n885);
    or g826(n1713 ,n1291 ,n870);
    or g827(n1712 ,n1179 ,n977);
    or g828(n1711 ,n1497 ,n1496);
    or g829(n1710 ,n1181 ,n884);
    or g830(n1709 ,n1495 ,n1494);
    or g831(n1708 ,n1178 ,n978);
    or g832(n1707 ,n1493 ,n1492);
    or g833(n1706 ,n1491 ,n1490);
    or g834(n1705 ,n1278 ,n882);
    or g835(n1704 ,n1489 ,n1488);
    or g836(n1703 ,n1176 ,n1019);
    or g837(n1702 ,n1177 ,n881);
    or g838(n1701 ,n1487 ,n1486);
    or g839(n1700 ,n1542 ,n1522);
    or g840(n1699 ,n1175 ,n1015);
    or g841(n1698 ,n1484 ,n1483);
    or g842(n1697 ,n1482 ,n1506);
    or g843(n1696 ,n1516 ,n1517);
    or g844(n1695 ,n1311 ,n1050);
    or g845(n1694 ,n1313 ,n1067);
    or g846(n1693 ,n1478 ,n1479);
    or g847(n1692 ,n1172 ,n1055);
    or g848(n1691 ,n1324 ,n1039);
    or g849(n1690 ,n1477 ,n1476);
    or g850(n1689 ,n1474 ,n1475);
    or g851(n1688 ,n1473 ,n1510);
    or g852(n1687 ,n1173 ,n875);
    or g853(n1686 ,n1511 ,n1471);
    or g854(n1685 ,n1363 ,n1108);
    or g855(n1684 ,n1350 ,n873);
    or g856(n1683 ,n1513 ,n1469);
    or g857(n1682 ,n1468 ,n1514);
    or g858(n1681 ,n1359 ,n872);
    or g859(n1680 ,n1467 ,n1466);
    or g860(n1679 ,n1362 ,n1064);
    or g861(n1678 ,n1465 ,n1524);
    or g862(n1677 ,n1464 ,n1463);
    or g863(n1676 ,n1462 ,n1534);
    or g864(n1675 ,n1171 ,n1077);
    or g865(n1674 ,n1366 ,n1066);
    or g866(n1673 ,n1461 ,n1537);
    or g867(n1672 ,n1460 ,n1541);
    or g868(n1671 ,n1170 ,n869);
    or g869(n1670 ,n1364 ,n862);
    or g870(n1669 ,n1457 ,n1458);
    or g871(n1668 ,n1456 ,n1455);
    or g872(n1667 ,n1376 ,n866);
    or g873(n1666 ,n1369 ,n868);
    or g874(n1665 ,n1454 ,n1453);
    or g875(n1664 ,n1452 ,n1451);
    or g876(n1663 ,n1377 ,n1079);
    or g877(n1662 ,n1449 ,n1450);
    or g878(n1661 ,n1550 ,n1448);
    or g879(n1660 ,n1168 ,n1072);
    or g880(n1659 ,n1447 ,n1446);
    or g881(n1658 ,n1385 ,n1082);
    or g882(n1657 ,n1445 ,n1574);
    or g883(n1656 ,n1165 ,n1087);
    or g884(n1655 ,n1166 ,n1099);
    or g885(n1654 ,n1444 ,n1443);
    or g886(n1653 ,n1442 ,n1581);
    or g887(n1652 ,n1384 ,n863);
    or g888(n1651 ,n1441 ,n1586);
    or g889(n1650 ,n1389 ,n1096);
    or g890(n1649 ,n1440 ,n1439);
    or g891(n1648 ,n1392 ,n1093);
    or g892(n1647 ,n1587 ,n1437);
    or g893(n1646 ,n1436 ,n1588);
    or g894(n1645 ,n1434 ,n1589);
    or g895(n1644 ,n1164 ,n861);
    or g896(n1643 ,n1432 ,n1431);
    or g897(n1642 ,n1163 ,n860);
    or g898(n1641 ,n1400 ,n1103);
    or g899(n1640 ,n1428 ,n1429);
    or g900(n1639 ,n1592 ,n1427);
    or g901(n1638 ,n1598 ,n1425);
    or g902(n1637 ,n1407 ,n1106);
    or g903(n1636 ,n1424 ,n1423);
    or g904(n1635 ,n1421 ,n1609);
    or g905(n1634 ,n1405 ,n856);
    or g906(n1633 ,n1161 ,n1107);
    or g907(n1632 ,n1158 ,n883);
    or g908(n1631 ,n1419 ,n1418);
    or g909(n1630 ,n1417 ,n1416);
    or g910(n1629 ,n1354 ,n1057);
    or g911(n1628 ,n1167 ,n855);
    or g912(n1627 ,n1329 ,n1062);
    or g913(n1626 ,n1409 ,n1073);
    or g914(n1625 ,n1415 ,n1472);
    or g915(n1624 ,n1414 ,n1413);
    or g916(n1623 ,n1412 ,n1411);
    or g917(n1622 ,n1410 ,n1532);
    nor g918(n1815 ,n1 ,n1157);
    nor g919(n1621 ,n474 ,n831);
    nor g920(n1620 ,n478 ,n803);
    nor g921(n1619 ,n170 ,n813);
    nor g922(n1618 ,n256 ,n833);
    nor g923(n1617 ,n421 ,n822);
    nor g924(n1616 ,n211 ,n827);
    nor g925(n1615 ,n415 ,n821);
    nor g926(n1614 ,n246 ,n819);
    nor g927(n1613 ,n165 ,n849);
    nor g928(n1612 ,n247 ,n825);
    nor g929(n1611 ,n416 ,n846);
    nor g930(n1610 ,n213 ,n824);
    nor g931(n1609 ,n212 ,n821);
    nor g932(n1608 ,n486 ,n822);
    nor g933(n1607 ,n436 ,n823);
    nor g934(n1606 ,n429 ,n822);
    nor g935(n1605 ,n475 ,n847);
    nor g936(n1604 ,n462 ,n821);
    nor g937(n1603 ,n445 ,n818);
    nor g938(n1602 ,n427 ,n846);
    nor g939(n1601 ,n250 ,n827);
    nor g940(n1600 ,n251 ,n849);
    nor g941(n1599 ,n181 ,n819);
    nor g942(n1598 ,n392 ,n827);
    nor g943(n1597 ,n202 ,n816);
    nor g944(n1596 ,n331 ,n826);
    nor g945(n1595 ,n230 ,n817);
    nor g946(n1594 ,n195 ,n848);
    nor g947(n1593 ,n205 ,n823);
    nor g948(n1592 ,n373 ,n847);
    nor g949(n1591 ,n396 ,n826);
    nor g950(n1590 ,n249 ,n822);
    nor g951(n1589 ,n245 ,n816);
    nor g952(n1588 ,n375 ,n847);
    nor g953(n1587 ,n198 ,n849);
    nor g954(n1586 ,n186 ,n846);
    nor g955(n1585 ,n234 ,n818);
    nor g956(n1584 ,n337 ,n849);
    nor g957(n1583 ,n456 ,n827);
    nor g958(n1582 ,n491 ,n848);
    nor g959(n1581 ,n443 ,n824);
    nor g960(n1580 ,n484 ,n824);
    nor g961(n1579 ,n364 ,n818);
    nor g962(n1578 ,n454 ,n825);
    nor g963(n1577 ,n380 ,n821);
    nor g964(n1576 ,n447 ,n822);
    nor g965(n1575 ,n347 ,n820);
    nor g966(n1574 ,n225 ,n823);
    nor g967(n1573 ,n369 ,n819);
    nor g968(n1572 ,n382 ,n817);
    nor g969(n1571 ,n460 ,n823);
    nor g970(n1570 ,n267 ,n847);
    nor g971(n1569 ,n237 ,n820);
    nor g972(n1568 ,n175 ,n825);
    nor g973(n1567 ,n450 ,n847);
    nor g974(n1566 ,n226 ,n824);
    nor g975(n1565 ,n349 ,n816);
    nor g976(n1564 ,n467 ,n821);
    nor g977(n1563 ,n169 ,n822);
    nor g978(n1562 ,n477 ,n849);
    nor g979(n1561 ,n494 ,n826);
    nor g980(n1560 ,n319 ,n817);
    nor g981(n1559 ,n441 ,n827);
    nor g982(n1558 ,n466 ,n848);
    nor g983(n1557 ,n442 ,n820);
    nor g984(n1556 ,n362 ,n818);
    nor g985(n1555 ,n374 ,n819);
    nor g986(n1554 ,n434 ,n822);
    nor g987(n1553 ,n256 ,n848);
    nor g988(n1552 ,n385 ,n818);
    nor g989(n1551 ,n412 ,n825);
    nor g990(n1550 ,n330 ,n820);
    nor g991(n1549 ,n403 ,n827);
    nor g992(n1548 ,n391 ,n823);
    nor g993(n1547 ,n489 ,n826);
    nor g994(n1546 ,n482 ,n820);
    nor g995(n1545 ,n465 ,n849);
    nor g996(n1544 ,n209 ,n816);
    nor g997(n1543 ,n345 ,n817);
    nor g998(n1542 ,n402 ,n820);
    nor g999(n1541 ,n218 ,n818);
    nor g1000(n1540 ,n401 ,n849);
    nor g1001(n1539 ,n410 ,n848);
    nor g1002(n1538 ,n196 ,n847);
    nor g1003(n1537 ,n274 ,n823);
    nor g1004(n1536 ,n210 ,n816);
    nor g1005(n1535 ,n469 ,n821);
    nor g1006(n1534 ,n471 ,n816);
    nor g1007(n1533 ,n383 ,n821);
    nor g1008(n1532 ,n406 ,n816);
    nor g1009(n1531 ,n389 ,n847);
    nor g1010(n1530 ,n399 ,n825);
    nor g1011(n1529 ,n321 ,n817);
    nor g1012(n1528 ,n338 ,n824);
    nor g1013(n1527 ,n451 ,n846);
    nor g1014(n1526 ,n190 ,n827);
    nor g1015(n1525 ,n189 ,n827);
    nor g1016(n1524 ,n278 ,n826);
    nor g1017(n1523 ,n457 ,n848);
    nor g1018(n1522 ,n352 ,n817);
    nor g1019(n1521 ,n328 ,n846);
    nor g1020(n1520 ,n240 ,n826);
    nor g1021(n1519 ,n359 ,n849);
    nor g1022(n1518 ,n390 ,n825);
    nor g1023(n1517 ,n229 ,n823);
    nor g1024(n1516 ,n253 ,n816);
    nor g1025(n1515 ,n259 ,n818);
    nor g1026(n1514 ,n468 ,n824);
    nor g1027(n1513 ,n159 ,n825);
    nor g1028(n1512 ,n409 ,n824);
    nor g1029(n1511 ,n236 ,n816);
    nor g1030(n1510 ,n407 ,n817);
    nor g1031(n1509 ,n242 ,n823);
    nor g1032(n1508 ,n262 ,n846);
    nor g1033(n1507 ,n370 ,n819);
    nor g1034(n1506 ,n206 ,n823);
    nor g1035(n1505 ,n473 ,n846);
    nor g1036(n1504 ,n325 ,n816);
    nor g1037(n1503 ,n340 ,n826);
    nor g1038(n1502 ,n426 ,n823);
    nor g1039(n1501 ,n487 ,n826);
    nor g1040(n1500 ,n188 ,n819);
    nor g1041(n1499 ,n207 ,n824);
    nor g1042(n1498 ,n255 ,n816);
    nor g1043(n1497 ,n384 ,n822);
    nor g1044(n1496 ,n366 ,n817);
    nor g1045(n1495 ,n176 ,n825);
    nor g1046(n1494 ,n203 ,n820);
    nor g1047(n1493 ,n493 ,n849);
    nor g1048(n1492 ,n243 ,n826);
    nor g1049(n1491 ,n397 ,n827);
    nor g1050(n1490 ,n170 ,n846);
    nor g1051(n1489 ,n219 ,n821);
    nor g1052(n1488 ,n244 ,n848);
    nor g1053(n1487 ,n372 ,n847);
    nor g1054(n1486 ,n419 ,n818);
    nor g1055(n1485 ,n459 ,n847);
    nor g1056(n1484 ,n233 ,n820);
    nor g1057(n1483 ,n368 ,n824);
    nor g1058(n1482 ,n408 ,n848);
    nor g1059(n1481 ,n356 ,n825);
    nor g1060(n1480 ,n266 ,n849);
    nor g1061(n1479 ,n343 ,n827);
    nor g1062(n1478 ,n363 ,n826);
    nor g1063(n1477 ,n200 ,n821);
    nor g1064(n1476 ,n248 ,n819);
    nor g1065(n1475 ,n265 ,n818);
    nor g1066(n1474 ,n453 ,n822);
    nor g1067(n1473 ,n217 ,n847);
    nor g1068(n1472 ,n458 ,n817);
    nor g1069(n1471 ,n238 ,n846);
    nor g1070(n1470 ,n439 ,n824);
    nor g1071(n1469 ,n400 ,n817);
    nor g1072(n1468 ,n271 ,n848);
    nor g1073(n1467 ,n326 ,n822);
    nor g1074(n1466 ,n420 ,n847);
    nor g1075(n1465 ,n276 ,n849);
    nor g1076(n1464 ,n194 ,n821);
    nor g1077(n1463 ,n336 ,n827);
    nor g1078(n1462 ,n197 ,n820);
    nor g1079(n1461 ,n172 ,n819);
    nor g1080(n1460 ,n485 ,n846);
    nor g1081(n1459 ,n158 ,n821);
    nor g1082(n1458 ,n220 ,n824);
    nor g1083(n1457 ,n463 ,n849);
    nor g1084(n1456 ,n241 ,n822);
    nor g1085(n1455 ,n481 ,n818);
    nor g1086(n1454 ,n180 ,n827);
    nor g1087(n1453 ,n269 ,n819);
    nor g1088(n1452 ,n232 ,n821);
    nor g1089(n1451 ,n273 ,n847);
    nor g1090(n1450 ,n472 ,n848);
    nor g1091(n1449 ,n174 ,n825);
    nor g1092(n1448 ,n222 ,n816);
    nor g1093(n1447 ,n449 ,n826);
    nor g1094(n1446 ,n227 ,n817);
    nor g1095(n1445 ,n438 ,n846);
    nor g1096(n1444 ,n452 ,n827);
    nor g1097(n1443 ,n394 ,n848);
    nor g1098(n1442 ,n346 ,n825);
    nor g1099(n1441 ,n387 ,n822);
    nor g1100(n1440 ,n187 ,n817);
    nor g1101(n1439 ,n333 ,n823);
    nor g1102(n1438 ,n272 ,n819);
    nor g1103(n1437 ,n418 ,n821);
    nor g1104(n1436 ,n323 ,n826);
    nor g1105(n1435 ,n177 ,n825);
    nor g1106(n1434 ,n425 ,n819);
    nor g1107(n1433 ,n268 ,n820);
    nor g1108(n1432 ,n182 ,n820);
    nor g1109(n1431 ,n235 ,n818);
    nor g1110(n1430 ,n260 ,n846);
    nor g1111(n1429 ,n398 ,n816);
    nor g1112(n1428 ,n348 ,n820);
    nor g1113(n1427 ,n483 ,n818);
    nor g1114(n1426 ,n492 ,n819);
    nor g1115(n1425 ,n166 ,n817);
    nor g1116(n1424 ,n379 ,n825);
    nor g1117(n1423 ,n320 ,n848);
    nor g1118(n1422 ,n461 ,n824);
    nor g1119(n1421 ,n258 ,n849);
    nor g1120(n1420 ,n191 ,n819);
    nor g1121(n1419 ,n353 ,n822);
    nor g1122(n1418 ,n332 ,n823);
    nor g1123(n1417 ,n490 ,n824);
    nor g1124(n1416 ,n339 ,n846);
    nor g1125(n1415 ,n367 ,n848);
    nor g1126(n1414 ,n479 ,n820);
    nor g1127(n1413 ,n214 ,n823);
    nor g1128(n1412 ,n184 ,n826);
    nor g1129(n1411 ,n480 ,n818);
    nor g1130(n1410 ,n335 ,n847);
    nor g1131(n1409 ,n390 ,n829);
    nor g1132(n1408 ,n389 ,n811);
    nor g1133(n1407 ,n412 ,n829);
    nor g1134(n1406 ,n408 ,n833);
    nor g1135(n1405 ,n267 ,n811);
    nor g1136(n1404 ,n368 ,n845);
    nor g1137(n1403 ,n205 ,n805);
    nor g1138(n1402 ,n271 ,n833);
    nor g1139(n1401 ,n320 ,n833);
    nor g1140(n1400 ,n175 ,n829);
    nor g1141(n1399 ,n367 ,n833);
    nor g1142(n1398 ,n459 ,n811);
    nor g1143(n1397 ,n195 ,n833);
    nor g1144(n1396 ,n228 ,n833);
    nor g1145(n1395 ,n426 ,n805);
    nor g1146(n1394 ,n329 ,n833);
    nor g1147(n1393 ,n491 ,n833);
    nor g1148(n1392 ,n378 ,n829);
    nor g1149(n1391 ,n391 ,n805);
    nor g1150(n1390 ,n380 ,n835);
    nor g1151(n1389 ,n476 ,n811);
    nor g1152(n1388 ,n234 ,n807);
    nor g1153(n1387 ,n324 ,n833);
    nor g1154(n1386 ,n274 ,n805);
    nor g1155(n1385 ,n247 ,n829);
    nor g1156(n1384 ,n261 ,n829);
    nor g1157(n1383 ,n219 ,n835);
    nor g1158(n1382 ,n259 ,n807);
    nor g1159(n1381 ,n200 ,n835);
    nor g1160(n1380 ,n332 ,n805);
    nor g1161(n1379 ,n460 ,n805);
    nor g1162(n1378 ,n214 ,n805);
    nor g1163(n1377 ,n379 ,n829);
    nor g1164(n1376 ,n335 ,n811);
    nor g1165(n1375 ,n250 ,n837);
    nor g1166(n1374 ,n462 ,n835);
    nor g1167(n1373 ,n172 ,n839);
    nor g1168(n1372 ,n192 ,n835);
    nor g1169(n1371 ,n207 ,n845);
    nor g1170(n1370 ,n357 ,n805);
    nor g1171(n1369 ,n346 ,n829);
    nor g1172(n1368 ,n467 ,n835);
    nor g1173(n1367 ,n422 ,n805);
    nor g1174(n1366 ,n159 ,n829);
    nor g1175(n1365 ,n248 ,n839);
    nor g1176(n1364 ,n364 ,n807);
    nor g1177(n1363 ,n244 ,n833);
    nor g1178(n1362 ,n356 ,n829);
    nor g1179(n1361 ,n419 ,n807);
    nor g1180(n1360 ,n188 ,n839);
    nor g1181(n1359 ,n375 ,n811);
    nor g1182(n1358 ,n242 ,n805);
    nor g1183(n1357 ,n196 ,n811);
    nor g1184(n1356 ,n269 ,n839);
    nor g1185(n1355 ,n415 ,n835);
    nor g1186(n1354 ,n254 ,n805);
    nor g1187(n1353 ,n425 ,n839);
    nor g1188(n1352 ,n436 ,n805);
    nor g1189(n1351 ,n191 ,n839);
    nor g1190(n1350 ,n176 ,n829);
    nor g1191(n1349 ,n246 ,n839);
    nor g1192(n1348 ,n229 ,n805);
    nor g1193(n1347 ,n181 ,n839);
    nor g1194(n1346 ,n212 ,n835);
    nor g1195(n1345 ,n430 ,n839);
    nor g1196(n1344 ,n203 ,n843);
    nor g1197(n1343 ,n354 ,n839);
    nor g1198(n1342 ,n220 ,n845);
    nor g1199(n1341 ,n369 ,n839);
    nor g1200(n1340 ,n443 ,n845);
    nor g1201(n1339 ,n233 ,n843);
    nor g1202(n1338 ,n370 ,n839);
    nor g1203(n1337 ,n374 ,n839);
    nor g1204(n1336 ,n361 ,n839);
    nor g1205(n1335 ,n197 ,n843);
    nor g1206(n1334 ,n158 ,n835);
    nor g1207(n1333 ,n272 ,n839);
    nor g1208(n1332 ,n490 ,n845);
    nor g1209(n1331 ,n492 ,n839);
    nor g1210(n1330 ,n330 ,n843);
    nor g1211(n1329 ,n450 ,n811);
    nor g1212(n1328 ,n418 ,n835);
    nor g1213(n1327 ,n243 ,n841);
    nor g1214(n1326 ,n363 ,n841);
    nor g1215(n1325 ,n182 ,n843);
    nor g1216(n1324 ,n210 ,n809);
    nor g1217(n1323 ,n232 ,n835);
    nor g1218(n1322 ,n278 ,n841);
    nor g1219(n1321 ,n213 ,n845);
    nor g1220(n1320 ,n265 ,n807);
    nor g1221(n1319 ,n348 ,n843);
    nor g1222(n1318 ,n449 ,n841);
    nor g1223(n1317 ,n404 ,n835);
    nor g1224(n1316 ,n323 ,n841);
    nor g1225(n1315 ,n487 ,n841);
    nor g1226(n1314 ,n479 ,n843);
    nor g1227(n1313 ,n327 ,n809);
    nor g1228(n1312 ,n184 ,n841);
    nor g1229(n1311 ,n420 ,n811);
    nor g1230(n1310 ,n194 ,n835);
    nor g1231(n1309 ,n268 ,n843);
    nor g1232(n1308 ,n331 ,n841);
    nor g1233(n1307 ,n199 ,n841);
    nor g1234(n1306 ,n439 ,n845);
    nor g1235(n1305 ,n428 ,n845);
    nor g1236(n1304 ,n215 ,n841);
    nor g1237(n1303 ,n216 ,n843);
    nor g1238(n1302 ,n340 ,n841);
    nor g1239(n1301 ,n432 ,n843);
    nor g1240(n1300 ,n494 ,n841);
    nor g1241(n1299 ,n489 ,n841);
    nor g1242(n1298 ,n405 ,n841);
    nor g1243(n1297 ,n347 ,n843);
    nor g1244(n1296 ,n333 ,n805);
    nor g1245(n1295 ,n163 ,n845);
    nor g1246(n1294 ,n396 ,n841);
    nor g1247(n1293 ,n442 ,n843);
    nor g1248(n1292 ,n240 ,n841);
    nor g1249(n1291 ,n488 ,n807);
    nor g1250(n1290 ,n397 ,n837);
    nor g1251(n1289 ,n482 ,n843);
    nor g1252(n1288 ,n343 ,n837);
    nor g1253(n1287 ,n484 ,n845);
    nor g1254(n1286 ,n336 ,n837);
    nor g1255(n1285 ,n185 ,n843);
    nor g1256(n1284 ,n180 ,n837);
    nor g1257(n1283 ,n452 ,n837);
    nor g1258(n1282 ,n237 ,n843);
    nor g1259(n1281 ,n392 ,n837);
    nor g1260(n1280 ,n225 ,n805);
    nor g1261(n1279 ,n211 ,n837);
    nor g1262(n1278 ,n325 ,n809);
    nor g1263(n1277 ,n468 ,n845);
    nor g1264(n1276 ,n402 ,n843);
    nor g1265(n1275 ,n193 ,n837);
    nor g1266(n1274 ,n226 ,n845);
    nor g1267(n1273 ,n218 ,n807);
    nor g1268(n1272 ,n366 ,n831);
    nor g1269(n1271 ,n377 ,n837);
    nor g1270(n1270 ,n457 ,n833);
    nor g1271(n1269 ,n409 ,n845);
    nor g1272(n1268 ,n456 ,n837);
    nor g1273(n1267 ,n441 ,n837);
    nor g1274(n1266 ,n407 ,n831);
    nor g1275(n1265 ,n328 ,n813);
    nor g1276(n1264 ,n403 ,n837);
    nor g1277(n1263 ,n161 ,n835);
    nor g1278(n1262 ,n464 ,n837);
    nor g1279(n1261 ,n400 ,n831);
    nor g1280(n1260 ,n190 ,n837);
    nor g1281(n1259 ,n275 ,n845);
    nor g1282(n1258 ,n189 ,n837);
    nor g1283(n1257 ,n410 ,n833);
    nor g1284(n1256 ,n227 ,n831);
    nor g1285(n1255 ,n493 ,n803);
    nor g1286(n1254 ,n266 ,n803);
    nor g1287(n1253 ,n338 ,n845);
    nor g1288(n1252 ,n187 ,n831);
    nor g1289(n1251 ,n276 ,n803);
    nor g1290(n1250 ,n463 ,n803);
    nor g1291(n1249 ,n166 ,n831);
    nor g1292(n1248 ,n198 ,n803);
    nor g1293(n1247 ,n481 ,n807);
    nor g1294(n1246 ,n258 ,n803);
    nor g1295(n1245 ,n165 ,n803);
    nor g1296(n1244 ,n458 ,n831);
    nor g1297(n1243 ,n251 ,n803);
    nor g1298(n1242 ,n461 ,n845);
    nor g1299(n1241 ,n230 ,n831);
    nor g1300(n1240 ,n411 ,n803);
    nor g1301(n1239 ,n206 ,n805);
    nor g1302(n1238 ,n337 ,n803);
    nor g1303(n1237 ,n477 ,n803);
    nor g1304(n1236 ,n342 ,n831);
    nor g1305(n1235 ,n465 ,n803);
    nor g1306(n1234 ,n381 ,n803);
    nor g1307(n1233 ,n401 ,n803);
    nor g1308(n1232 ,n382 ,n831);
    nor g1309(n1231 ,n359 ,n803);
    nor g1310(n1230 ,n238 ,n813);
    nor g1311(n1229 ,n319 ,n831);
    nor g1312(n1228 ,n345 ,n831);
    nor g1313(n1227 ,n235 ,n807);
    nor g1314(n1226 ,n355 ,n831);
    nor g1315(n1225 ,n466 ,n833);
    nor g1316(n1224 ,n485 ,n813);
    nor g1317(n1223 ,n483 ,n807);
    nor g1318(n1222 ,n321 ,n831);
    nor g1319(n1221 ,n438 ,n813);
    nor g1320(n1220 ,n352 ,n831);
    nor g1321(n1219 ,n384 ,n815);
    nor g1322(n1218 ,n186 ,n813);
    nor g1323(n1217 ,n453 ,n815);
    nor g1324(n1216 ,n326 ,n815);
    nor g1325(n1215 ,n339 ,n813);
    nor g1326(n1214 ,n241 ,n815);
    nor g1327(n1213 ,n387 ,n815);
    nor g1328(n1212 ,n353 ,n815);
    nor g1329(n1211 ,n416 ,n813);
    nor g1330(n1210 ,n421 ,n815);
    nor g1331(n1209 ,n427 ,n813);
    nor g1332(n1208 ,n429 ,n815);
    nor g1333(n1207 ,n178 ,n815);
    nor g1334(n1206 ,n264 ,n815);
    nor g1335(n1205 ,n440 ,n813);
    nor g1336(n1204 ,n480 ,n807);
    nor g1337(n1203 ,n447 ,n815);
    nor g1338(n1202 ,n437 ,n813);
    nor g1339(n1201 ,n169 ,n815);
    nor g1340(n1200 ,n434 ,n815);
    nor g1341(n1199 ,n414 ,n815);
    nor g1342(n1198 ,n473 ,n813);
    nor g1343(n1197 ,n486 ,n815);
    nor g1344(n1196 ,n445 ,n807);
    nor g1345(n1195 ,n262 ,n813);
    nor g1346(n1194 ,n249 ,n815);
    nor g1347(n1193 ,n255 ,n809);
    nor g1348(n1192 ,n451 ,n813);
    nor g1349(n1191 ,n236 ,n809);
    nor g1350(n1190 ,n471 ,n809);
    nor g1351(n1189 ,n239 ,n813);
    nor g1352(n1188 ,n222 ,n809);
    nor g1353(n1187 ,n245 ,n809);
    nor g1354(n1186 ,n260 ,n813);
    nor g1355(n1185 ,n398 ,n809);
    nor g1356(n1184 ,n224 ,n807);
    nor g1357(n1183 ,n406 ,n809);
    nor g1358(n1182 ,n202 ,n809);
    nor g1359(n1181 ,n431 ,n809);
    nor g1360(n1180 ,n469 ,n835);
    nor g1361(n1179 ,n372 ,n811);
    nor g1362(n1178 ,n395 ,n809);
    nor g1363(n1177 ,n349 ,n809);
    nor g1364(n1176 ,n217 ,n811);
    nor g1365(n1175 ,n209 ,n809);
    nor g1366(n1174 ,n433 ,n807);
    nor g1367(n1173 ,n253 ,n809);
    nor g1368(n1172 ,n273 ,n811);
    nor g1369(n1171 ,n373 ,n811);
    nor g1370(n1170 ,n174 ,n829);
    nor g1371(n1169 ,n394 ,n833);
    nor g1372(n1168 ,n362 ,n807);
    nor g1373(n1167 ,n399 ,n829);
    nor g1374(n1166 ,n177 ,n829);
    nor g1375(n1165 ,n475 ,n811);
    nor g1376(n1164 ,n454 ,n829);
    nor g1377(n1163 ,n413 ,n811);
    nor g1378(n1162 ,n472 ,n833);
    nor g1379(n1161 ,n417 ,n829);
    nor g1380(n1160 ,n383 ,n835);
    nor g1381(n1159 ,n322 ,n811);
    nor g1382(n1158 ,n385 ,n807);
    nor g1383(n1157 ,n26[4] ,n850);
    nor g1384(n1156 ,n18[13] ,n848);
    nor g1385(n1155 ,n23[8] ,n849);
    nor g1386(n1154 ,n13[8] ,n820);
    nor g1387(n1153 ,n21[8] ,n826);
    nor g1388(n1152 ,n22[8] ,n827);
    nor g1389(n1151 ,n14[8] ,n817);
    nor g1390(n1150 ,n18[8] ,n848);
    nor g1391(n1149 ,n10[8] ,n846);
    nor g1392(n1148 ,n8[8] ,n818);
    nor g1393(n1147 ,n15[9] ,n822);
    nor g1394(n1146 ,n23[9] ,n849);
    nor g1395(n1145 ,n18[9] ,n848);
    nor g1396(n1144 ,n21[9] ,n826);
    nor g1397(n1143 ,n10[13] ,n846);
    nor g1398(n1142 ,n17[9] ,n825);
    nor g1399(n1141 ,n11[9] ,n847);
    nor g1400(n1140 ,n8[9] ,n818);
    nor g1401(n1139 ,n14[13] ,n817);
    nor g1402(n1138 ,n9[13] ,n824);
    nor g1403(n1137 ,n12[13] ,n823);
    nor g1404(n1136 ,n11[13] ,n847);
    nor g1405(n1135 ,n17[13] ,n825);
    nor g1406(n1134 ,n8[13] ,n818);
    nor g1407(n1133 ,n13[13] ,n820);
    nor g1408(n1132 ,n21[13] ,n826);
    nor g1409(n1131 ,n16[13] ,n816);
    nor g1410(n1130 ,n23[13] ,n849);
    nor g1411(n1129 ,n22[13] ,n827);
    nor g1412(n1128 ,n20[13] ,n819);
    nor g1413(n1127 ,n12[9] ,n823);
    nor g1414(n1126 ,n15[13] ,n822);
    nor g1415(n1125 ,n16[9] ,n816);
    nor g1416(n1124 ,n10[9] ,n846);
    nor g1417(n1123 ,n19[8] ,n821);
    nor g1418(n1122 ,n14[9] ,n817);
    nor g1419(n1121 ,n20[9] ,n819);
    nor g1420(n1120 ,n19[9] ,n821);
    nor g1421(n1119 ,n13[9] ,n820);
    nor g1422(n1118 ,n9[8] ,n824);
    nor g1423(n1117 ,n9[9] ,n824);
    nor g1424(n1116 ,n19[13] ,n821);
    nor g1425(n1115 ,n12[8] ,n823);
    nor g1426(n1114 ,n22[9] ,n827);
    nor g1427(n1113 ,n11[8] ,n847);
    nor g1428(n1112 ,n15[8] ,n822);
    nor g1429(n1111 ,n20[8] ,n819);
    nor g1430(n1110 ,n16[8] ,n816);
    nor g1431(n1109 ,n17[8] ,n825);
    nor g1432(n1108 ,n571 ,n832);
    nor g1433(n1107 ,n562 ,n828);
    nor g1434(n1106 ,n560 ,n828);
    nor g1435(n1105 ,n567 ,n832);
    nor g1436(n1104 ,n562 ,n810);
    nor g1437(n1103 ,n566 ,n828);
    nor g1438(n1102 ,n567 ,n838);
    nor g1439(n1101 ,n570 ,n832);
    nor g1440(n1100 ,n569 ,n832);
    nor g1441(n1099 ,n569 ,n828);
    nor g1442(n1098 ,n564 ,n804);
    nor g1443(n1097 ,n563 ,n832);
    nor g1444(n1096 ,n564 ,n810);
    nor g1445(n1095 ,n559 ,n832);
    nor g1446(n1094 ,n565 ,n832);
    nor g1447(n1093 ,n563 ,n828);
    nor g1448(n1092 ,n566 ,n832);
    nor g1449(n1091 ,n566 ,n836);
    nor g1450(n1090 ,n561 ,n832);
    nor g1451(n1089 ,n562 ,n832);
    nor g1452(n1088 ,n560 ,n810);
    nor g1453(n1087 ,n569 ,n810);
    nor g1454(n1086 ,n563 ,n834);
    nor g1455(n1085 ,n559 ,n838);
    nor g1456(n1084 ,n571 ,n834);
    nor g1457(n1083 ,n568 ,n834);
    nor g1458(n1082 ,n570 ,n828);
    nor g1459(n1081 ,n564 ,n836);
    nor g1460(n1080 ,n561 ,n834);
    nor g1461(n1079 ,n573 ,n828);
    nor g1462(n1078 ,n570 ,n804);
    nor g1463(n1077 ,n573 ,n810);
    nor g1464(n1076 ,n571 ,n844);
    nor g1465(n1075 ,n569 ,n804);
    nor g1466(n1074 ,n564 ,n834);
    nor g1467(n1073 ,n561 ,n828);
    nor g1468(n1072 ,n566 ,n806);
    nor g1469(n1071 ,n565 ,n834);
    nor g1470(n1070 ,n565 ,n804);
    nor g1471(n1069 ,n566 ,n834);
    nor g1472(n1068 ,n563 ,n804);
    nor g1473(n1067 ,n562 ,n808);
    nor g1474(n1066 ,n568 ,n828);
    nor g1475(n1065 ,n574 ,n834);
    nor g1476(n1064 ,n559 ,n828);
    nor g1477(n1063 ,n566 ,n804);
    nor g1478(n1062 ,n566 ,n810);
    nor g1479(n1061 ,n568 ,n832);
    nor g1480(n1060 ,n565 ,n844);
    nor g1481(n1059 ,n570 ,n834);
    nor g1482(n1058 ,n573 ,n834);
    nor g1483(n1057 ,n562 ,n804);
    nor g1484(n1056 ,n572 ,n838);
    nor g1485(n1055 ,n567 ,n810);
    nor g1486(n1054 ,n573 ,n838);
    nor g1487(n1053 ,n574 ,n804);
    nor g1488(n1052 ,n567 ,n844);
    nor g1489(n1051 ,n570 ,n838);
    nor g1490(n1050 ,n568 ,n810);
    nor g1491(n1049 ,n569 ,n838);
    nor g1492(n1048 ,n561 ,n804);
    nor g1493(n1047 ,n563 ,n844);
    nor g1494(n1046 ,n564 ,n838);
    nor g1495(n1045 ,n563 ,n838);
    nor g1496(n1044 ,n565 ,n838);
    nor g1497(n1043 ,n571 ,n842);
    nor g1498(n1042 ,n572 ,n844);
    nor g1499(n1041 ,n566 ,n838);
    nor g1500(n1040 ,n559 ,n842);
    nor g1501(n1039 ,n574 ,n808);
    nor g1502(n1038 ,n572 ,n834);
    nor g1503(n1037 ,n560 ,n838);
    nor g1504(n1036 ,n561 ,n806);
    nor g1505(n1035 ,n573 ,n804);
    nor g1506(n1034 ,n562 ,n838);
    nor g1507(n1033 ,n574 ,n838);
    nor g1508(n1032 ,n568 ,n842);
    nor g1509(n1031 ,n561 ,n838);
    nor g1510(n1030 ,n567 ,n842);
    nor g1511(n1029 ,n571 ,n840);
    nor g1512(n1028 ,n573 ,n844);
    nor g1513(n1027 ,n567 ,n834);
    nor g1514(n1026 ,n559 ,n840);
    nor g1515(n1025 ,n572 ,n842);
    nor g1516(n1024 ,n574 ,n840);
    nor g1517(n1023 ,n568 ,n840);
    nor g1518(n1022 ,n573 ,n842);
    nor g1519(n1021 ,n567 ,n840);
    nor g1520(n1020 ,n560 ,n804);
    nor g1521(n1019 ,n559 ,n810);
    nor g1522(n1018 ,n569 ,n834);
    nor g1523(n1017 ,n572 ,n840);
    nor g1524(n1016 ,n570 ,n844);
    nor g1525(n1015 ,n560 ,n808);
    nor g1526(n1014 ,n573 ,n840);
    nor g1527(n1013 ,n565 ,n840);
    nor g1528(n1012 ,n570 ,n842);
    nor g1529(n1011 ,n570 ,n840);
    nor g1530(n1010 ,n566 ,n840);
    nor g1531(n1009 ,n569 ,n842);
    nor g1532(n1008 ,n569 ,n840);
    nor g1533(n1007 ,n569 ,n844);
    nor g1534(n1006 ,n564 ,n840);
    nor g1535(n1005 ,n571 ,n806);
    nor g1536(n1004 ,n572 ,n804);
    nor g1537(n1003 ,n563 ,n840);
    nor g1538(n1002 ,n564 ,n842);
    nor g1539(n1001 ,n559 ,n834);
    nor g1540(n1000 ,n564 ,n844);
    nor g1541(n999 ,n563 ,n842);
    nor g1542(n998 ,n560 ,n840);
    nor g1543(n997 ,n562 ,n840);
    nor g1544(n996 ,n565 ,n842);
    nor g1545(n995 ,n561 ,n840);
    nor g1546(n994 ,n571 ,n836);
    nor g1547(n993 ,n566 ,n842);
    nor g1548(n992 ,n559 ,n836);
    nor g1549(n991 ,n560 ,n842);
    nor g1550(n990 ,n567 ,n804);
    nor g1551(n989 ,n568 ,n836);
    nor g1552(n988 ,n567 ,n836);
    nor g1553(n987 ,n562 ,n842);
    nor g1554(n986 ,n572 ,n836);
    nor g1555(n985 ,n573 ,n836);
    nor g1556(n984 ,n574 ,n842);
    nor g1557(n983 ,n574 ,n806);
    nor g1558(n982 ,n570 ,n836);
    nor g1559(n981 ,n569 ,n836);
    nor g1560(n980 ,n561 ,n842);
    nor g1561(n979 ,n566 ,n844);
    nor g1562(n978 ,n563 ,n808);
    nor g1563(n977 ,n571 ,n810);
    nor g1564(n976 ,n563 ,n836);
    nor g1565(n975 ,n559 ,n806);
    nor g1566(n974 ,n565 ,n836);
    nor g1567(n973 ,n571 ,n830);
    nor g1568(n972 ,n560 ,n844);
    nor g1569(n971 ,n574 ,n832);
    nor g1570(n970 ,n560 ,n836);
    nor g1571(n969 ,n559 ,n830);
    nor g1572(n968 ,n562 ,n836);
    nor g1573(n967 ,n571 ,n838);
    nor g1574(n966 ,n574 ,n836);
    nor g1575(n965 ,n561 ,n836);
    nor g1576(n964 ,n562 ,n844);
    nor g1577(n963 ,n567 ,n830);
    nor g1578(n962 ,n571 ,n802);
    nor g1579(n961 ,n568 ,n802);
    nor g1580(n960 ,n572 ,n830);
    nor g1581(n959 ,n562 ,n806);
    nor g1582(n958 ,n567 ,n802);
    nor g1583(n957 ,n573 ,n830);
    nor g1584(n956 ,n572 ,n802);
    nor g1585(n955 ,n574 ,n844);
    nor g1586(n954 ,n568 ,n806);
    nor g1587(n953 ,n573 ,n802);
    nor g1588(n952 ,n570 ,n802);
    nor g1589(n951 ,n570 ,n830);
    nor g1590(n950 ,n561 ,n844);
    nor g1591(n949 ,n569 ,n830);
    nor g1592(n948 ,n563 ,n802);
    nor g1593(n947 ,n559 ,n804);
    nor g1594(n946 ,n565 ,n802);
    nor g1595(n945 ,n564 ,n830);
    nor g1596(n944 ,n560 ,n802);
    nor g1597(n943 ,n563 ,n830);
    nor g1598(n942 ,n571 ,n812);
    nor g1599(n941 ,n574 ,n802);
    nor g1600(n940 ,n565 ,n830);
    nor g1601(n939 ,n561 ,n802);
    nor g1602(n938 ,n566 ,n830);
    nor g1603(n937 ,n571 ,n804);
    nor g1604(n936 ,n559 ,n812);
    nor g1605(n935 ,n560 ,n830);
    nor g1606(n934 ,n567 ,n806);
    nor g1607(n933 ,n562 ,n830);
    nor g1608(n932 ,n574 ,n830);
    nor g1609(n931 ,n568 ,n812);
    nor g1610(n930 ,n561 ,n830);
    nor g1611(n929 ,n571 ,n814);
    nor g1612(n928 ,n567 ,n812);
    nor g1613(n927 ,n559 ,n844);
    nor g1614(n926 ,n559 ,n814);
    nor g1615(n925 ,n572 ,n806);
    nor g1616(n924 ,n572 ,n812);
    nor g1617(n923 ,n568 ,n814);
    nor g1618(n922 ,n573 ,n812);
    nor g1619(n921 ,n567 ,n814);
    nor g1620(n920 ,n572 ,n814);
    nor g1621(n919 ,n573 ,n814);
    nor g1622(n918 ,n570 ,n812);
    nor g1623(n917 ,n570 ,n814);
    nor g1624(n916 ,n569 ,n814);
    nor g1625(n915 ,n564 ,n814);
    nor g1626(n914 ,n569 ,n812);
    nor g1627(n913 ,n568 ,n844);
    nor g1628(n912 ,n563 ,n814);
    nor g1629(n911 ,n564 ,n812);
    nor g1630(n910 ,n573 ,n806);
    nor g1631(n909 ,n565 ,n814);
    nor g1632(n908 ,n563 ,n812);
    nor g1633(n907 ,n566 ,n814);
    nor g1634(n906 ,n560 ,n814);
    nor g1635(n905 ,n564 ,n832);
    nor g1636(n904 ,n562 ,n814);
    nor g1637(n903 ,n565 ,n812);
    nor g1638(n902 ,n574 ,n814);
    nor g1639(n901 ,n566 ,n812);
    nor g1640(n900 ,n561 ,n814);
    nor g1641(n899 ,n570 ,n806);
    nor g1642(n898 ,n571 ,n808);
    nor g1643(n897 ,n560 ,n812);
    nor g1644(n896 ,n559 ,n808);
    nor g1645(n895 ,n561 ,n810);
    nor g1646(n894 ,n568 ,n808);
    nor g1647(n893 ,n562 ,n812);
    nor g1648(n892 ,n567 ,n808);
    nor g1649(n891 ,n572 ,n808);
    nor g1650(n890 ,n573 ,n808);
    nor g1651(n889 ,n574 ,n812);
    nor g1652(n888 ,n569 ,n806);
    nor g1653(n887 ,n570 ,n808);
    nor g1654(n886 ,n572 ,n832);
    nor g1655(n885 ,n569 ,n808);
    nor g1656(n884 ,n564 ,n808);
    nor g1657(n883 ,n560 ,n806);
    nor g1658(n882 ,n565 ,n808);
    nor g1659(n881 ,n566 ,n808);
    nor g1660(n880 ,n562 ,n802);
    nor g1661(n879 ,n564 ,n806);
    nor g1662(n878 ,n566 ,n802);
    nor g1663(n877 ,n573 ,n832);
    nor g1664(n876 ,n574 ,n810);
    nor g1665(n875 ,n561 ,n808);
    nor g1666(n874 ,n560 ,n832);
    nor g1667(n873 ,n571 ,n828);
    nor g1668(n872 ,n572 ,n810);
    nor g1669(n871 ,n564 ,n802);
    nor g1670(n870 ,n563 ,n806);
    nor g1671(n869 ,n567 ,n828);
    nor g1672(n868 ,n572 ,n828);
    nor g1673(n867 ,n569 ,n802);
    nor g1674(n866 ,n570 ,n810);
    nor g1675(n865 ,n568 ,n838);
    nor g1676(n864 ,n562 ,n834);
    nor g1677(n863 ,n564 ,n828);
    nor g1678(n862 ,n565 ,n806);
    nor g1679(n861 ,n565 ,n828);
    nor g1680(n860 ,n563 ,n810);
    nor g1681(n859 ,n561 ,n812);
    nor g1682(n858 ,n559 ,n802);
    nor g1683(n857 ,n568 ,n830);
    nor g1684(n856 ,n565 ,n810);
    nor g1685(n855 ,n574 ,n828);
    nor g1686(n854 ,n560 ,n834);
    nor g1687(n853 ,n568 ,n804);
    or g1688(n852 ,n702 ,n800);
    or g1689(n851 ,n712 ,n801);
    not g1690(n844 ,n845);
    not g1691(n842 ,n843);
    not g1692(n840 ,n841);
    not g1693(n838 ,n839);
    not g1694(n836 ,n837);
    not g1695(n834 ,n835);
    not g1696(n832 ,n833);
    not g1697(n830 ,n831);
    not g1698(n828 ,n829);
    or g1699(n850 ,n506 ,n769);
    or g1700(n849 ,n590 ,n774);
    or g1701(n848 ,n591 ,n772);
    or g1702(n847 ,n591 ,n777);
    or g1703(n846 ,n591 ,n775);
    nor g1704(n845 ,n520 ,n773);
    nor g1705(n843 ,n520 ,n794);
    nor g1706(n841 ,n522 ,n794);
    nor g1707(n839 ,n519 ,n794);
    nor g1708(n837 ,n519 ,n795);
    nor g1709(n835 ,n522 ,n776);
    nor g1710(n833 ,n519 ,n776);
    nor g1711(n831 ,n521 ,n795);
    nor g1712(n829 ,n522 ,n773);
    not g1713(n814 ,n815);
    not g1714(n812 ,n813);
    not g1715(n810 ,n811);
    not g1716(n808 ,n809);
    not g1717(n806 ,n807);
    not g1718(n804 ,n805);
    not g1719(n802 ,n803);
    nor g1720(n801 ,n753 ,n767);
    nor g1721(n800 ,n752 ,n768);
    or g1722(n799 ,n690 ,n757);
    or g1723(n798 ,n697 ,n758);
    or g1724(n797 ,n664 ,n756);
    or g1725(n796 ,n665 ,n766);
    or g1726(n827 ,n590 ,n772);
    or g1727(n826 ,n592 ,n774);
    or g1728(n825 ,n589 ,n774);
    or g1729(n824 ,n589 ,n777);
    or g1730(n823 ,n592 ,n775);
    or g1731(n822 ,n590 ,n777);
    or g1732(n821 ,n591 ,n774);
    or g1733(n820 ,n592 ,n777);
    or g1734(n819 ,n592 ,n772);
    or g1735(n818 ,n589 ,n775);
    or g1736(n817 ,n590 ,n775);
    or g1737(n816 ,n589 ,n772);
    nor g1738(n815 ,n520 ,n795);
    nor g1739(n813 ,n521 ,n776);
    nor g1740(n811 ,n520 ,n776);
    nor g1741(n809 ,n519 ,n773);
    nor g1742(n807 ,n521 ,n773);
    nor g1743(n805 ,n521 ,n794);
    nor g1744(n803 ,n522 ,n795);
    nor g1745(n793 ,n455 ,n747);
    nor g1746(n792 ,n334 ,n747);
    nor g1747(n791 ,n446 ,n747);
    nor g1748(n790 ,n423 ,n747);
    nor g1749(n789 ,n277 ,n747);
    nor g1750(n788 ,n376 ,n747);
    nor g1751(n787 ,n157 ,n747);
    nor g1752(n786 ,n371 ,n747);
    nor g1753(n785 ,n424 ,n747);
    nor g1754(n784 ,n470 ,n747);
    nor g1755(n783 ,n444 ,n747);
    nor g1756(n782 ,n435 ,n747);
    nor g1757(n781 ,n263 ,n747);
    nor g1758(n780 ,n257 ,n747);
    nor g1759(n779 ,n388 ,n747);
    nor g1760(n778 ,n448 ,n747);
    or g1761(n795 ,n307 ,n750);
    or g1762(n794 ,n307 ,n749);
    or g1763(n771 ,n700 ,n726);
    xnor g1764(n770 ,n498 ,n663);
    or g1765(n769 ,n508 ,n745);
    nor g1766(n768 ,n511 ,n730);
    nor g1767(n767 ,n512 ,n728);
    or g1768(n766 ,n713 ,n742);
    or g1769(n765 ,n703 ,n721);
    or g1770(n764 ,n716 ,n722);
    or g1771(n763 ,n686 ,n732);
    or g1772(n762 ,n718 ,n723);
    or g1773(n761 ,n707 ,n727);
    or g1774(n760 ,n705 ,n725);
    or g1775(n759 ,n714 ,n720);
    or g1776(n758 ,n719 ,n743);
    or g1777(n757 ,n709 ,n740);
    or g1778(n756 ,n711 ,n741);
    or g1779(n755 ,n642 ,n744);
    or g1780(n754 ,n694 ,n724);
    nor g1781(n753 ,n29[3] ,n729);
    nor g1782(n752 ,n29[2] ,n731);
    or g1783(n777 ,n27[3] ,n751);
    or g1784(n776 ,n28[2] ,n750);
    or g1785(n775 ,n27[3] ,n748);
    or g1786(n774 ,n306 ,n751);
    or g1787(n773 ,n28[2] ,n749);
    or g1788(n772 ,n306 ,n748);
    not g1789(n746 ,n747);
    or g1790(n745 ,n579 ,n691);
    nor g1791(n744 ,n582 ,n688);
    nor g1792(n743 ,n549 ,n681);
    nor g1793(n742 ,n551 ,n684);
    nor g1794(n741 ,n550 ,n683);
    nor g1795(n740 ,n547 ,n682);
    or g1796(n751 ,n309 ,n698);
    or g1797(n750 ,n310 ,n699);
    or g1798(n749 ,n28[1] ,n699);
    or g1799(n748 ,n27[0] ,n698);
    nor g1800(n747 ,n27[6] ,n698);
    or g1801(n739 ,n643 ,n677);
    or g1802(n738 ,n637 ,n678);
    or g1803(n737 ,n638 ,n687);
    or g1804(n736 ,n650 ,n673);
    or g1805(n735 ,n651 ,n672);
    or g1806(n734 ,n649 ,n671);
    or g1807(n733 ,n652 ,n670);
    or g1808(n732 ,n706 ,n689);
    or g1809(n731 ,n654 ,n717);
    or g1810(n730 ,n576 ,n680);
    or g1811(n729 ,n655 ,n715);
    or g1812(n728 ,n575 ,n685);
    or g1813(n727 ,n661 ,n692);
    or g1814(n726 ,n658 ,n693);
    or g1815(n725 ,n656 ,n696);
    or g1816(n724 ,n657 ,n701);
    or g1817(n723 ,n659 ,n704);
    or g1818(n722 ,n653 ,n708);
    or g1819(n721 ,n660 ,n695);
    or g1820(n720 ,n662 ,n710);
    nor g1821(n719 ,n150 ,n625);
    nor g1822(n718 ,n285 ,n623);
    nor g1823(n717 ,n173 ,n623);
    nor g1824(n716 ,n288 ,n623);
    nor g1825(n715 ,n231 ,n623);
    nor g1826(n714 ,n287 ,n623);
    nor g1827(n713 ,n315 ,n625);
    nor g1828(n712 ,n314 ,n625);
    nor g1829(n711 ,n153 ,n625);
    nor g1830(n710 ,n151 ,n625);
    nor g1831(n709 ,n155 ,n625);
    nor g1832(n708 ,n311 ,n625);
    nor g1833(n707 ,n156 ,n625);
    nor g1834(n706 ,n154 ,n625);
    nor g1835(n705 ,n152 ,n625);
    nor g1836(n704 ,n313 ,n625);
    nor g1837(n703 ,n312 ,n625);
    nor g1838(n702 ,n317 ,n625);
    nor g1839(n701 ,n149 ,n625);
    nor g1840(n700 ,n318 ,n625);
    nor g1841(n697 ,n585 ,n606);
    nor g1842(n696 ,n293 ,n623);
    nor g1843(n695 ,n297 ,n623);
    nor g1844(n694 ,n295 ,n623);
    nor g1845(n693 ,n301 ,n623);
    nor g1846(n692 ,n280 ,n623);
    or g1847(n691 ,n517 ,n620);
    nor g1848(n690 ,n585 ,n605);
    nor g1849(n689 ,n627 ,n623);
    or g1850(n688 ,n513 ,n628);
    nor g1851(n687 ,n580 ,n616);
    nor g1852(n686 ,n626 ,n628);
    nor g1853(n685 ,n2248 ,n623);
    or g1854(n684 ,n502 ,n623);
    or g1855(n683 ,n518 ,n623);
    or g1856(n682 ,n514 ,n623);
    or g1857(n681 ,n516 ,n623);
    nor g1858(n680 ,n2249 ,n623);
    or g1859(n679 ,n630 ,n639);
    nor g1860(n678 ,n585 ,n610);
    nor g1861(n677 ,n585 ,n602);
    or g1862(n676 ,n622 ,n644);
    or g1863(n675 ,n631 ,n641);
    or g1864(n674 ,n629 ,n640);
    nor g1865(n673 ,n587 ,n597);
    nor g1866(n672 ,n587 ,n599);
    nor g1867(n671 ,n587 ,n598);
    nor g1868(n670 ,n587 ,n594);
    or g1869(n669 ,n633 ,n648);
    or g1870(n668 ,n634 ,n645);
    or g1871(n667 ,n636 ,n647);
    or g1872(n666 ,n635 ,n646);
    nor g1873(n665 ,n585 ,n604);
    nor g1874(n664 ,n585 ,n607);
    nor g1875(n663 ,n29[0] ,n624);
    or g1876(n699 ,n510 ,n632);
    or g1877(n698 ,n515 ,n619);
    nor g1878(n662 ,n286 ,n588);
    nor g1879(n661 ,n291 ,n588);
    nor g1880(n660 ,n290 ,n588);
    nor g1881(n659 ,n279 ,n588);
    nor g1882(n658 ,n282 ,n588);
    nor g1883(n657 ,n299 ,n588);
    nor g1884(n656 ,n296 ,n588);
    nor g1885(n655 ,n164 ,n588);
    nor g1886(n654 ,n167 ,n588);
    nor g1887(n653 ,n284 ,n588);
    nor g1888(n652 ,n350 ,n586);
    nor g1889(n651 ,n351 ,n586);
    nor g1890(n650 ,n208 ,n586);
    nor g1891(n649 ,n270 ,n586);
    nor g1892(n648 ,n252 ,n586);
    nor g1893(n647 ,n201 ,n586);
    nor g1894(n646 ,n341 ,n586);
    nor g1895(n645 ,n221 ,n586);
    nor g1896(n644 ,n223 ,n584);
    nor g1897(n643 ,n358 ,n584);
    nor g1898(n642 ,n344 ,n584);
    nor g1899(n641 ,n386 ,n584);
    nor g1900(n640 ,n365 ,n584);
    nor g1901(n639 ,n393 ,n584);
    nor g1902(n638 ,n360 ,n584);
    nor g1903(n637 ,n204 ,n584);
    nor g1904(n636 ,n146 ,n587);
    nor g1905(n635 ,n143 ,n587);
    nor g1906(n634 ,n145 ,n587);
    nor g1907(n633 ,n144 ,n587);
    or g1908(n632 ,n501 ,n577);
    nor g1909(n631 ,n133 ,n585);
    nor g1910(n630 ,n136 ,n585);
    nor g1911(n629 ,n134 ,n585);
    not g1912(n627 ,n626);
    not g1913(n625 ,n624);
    nor g1914(n622 ,n135 ,n585);
    xnor g1915(n621 ,n145 ,n497);
    or g1916(n620 ,n26[15] ,n578);
    or g1917(n619 ,n27[7] ,n588);
    xnor g1918(n618 ,n143 ,n495);
    xnor g1919(n617 ,n144 ,n537);
    or g1920(n616 ,n585 ,n583);
    xnor g1921(n615 ,n146 ,n526);
    xnor g1922(n614 ,n131 ,n529);
    xnor g1923(n613 ,n132 ,n532);
    xnor g1924(n612 ,n133 ,n528);
    xnor g1925(n611 ,n136 ,n543);
    xnor g1926(n610 ,n29[0] ,n500);
    xnor g1927(n609 ,n134 ,n545);
    xnor g1928(n608 ,n135 ,n538);
    xnor g1929(n607 ,n29[5] ,n546);
    xnor g1930(n606 ,n29[7] ,n534);
    xnor g1931(n605 ,n29[6] ,n496);
    xnor g1932(n604 ,n29[4] ,n531);
    xnor g1933(n603 ,n137 ,n544);
    xnor g1934(n602 ,n29[2] ,n527);
    xnor g1935(n601 ,n138 ,n536);
    xnor g1936(n600 ,n141 ,n541);
    xnor g1937(n599 ,n29[9] ,n539);
    xnor g1938(n598 ,n29[10] ,n540);
    xnor g1939(n597 ,n29[8] ,n499);
    xnor g1940(n596 ,n139 ,n535);
    xnor g1941(n595 ,n140 ,n530);
    xnor g1942(n594 ,n29[11] ,n542);
    xnor g1943(n593 ,n142 ,n533);
    or g1944(n628 ,n509 ,n585);
    nor g1945(n626 ,n548 ,n581);
    nor g1946(n624 ,n552 ,n586);
    or g1947(n623 ,n555 ,n584);
    not g1948(n586 ,n587);
    not g1949(n584 ,n585);
    nor g1950(n583 ,n29[3] ,n557);
    nor g1951(n582 ,n168 ,n525);
    nor g1952(n581 ,n2250 ,n524);
    nor g1953(n580 ,n138 ,n558);
    or g1954(n579 ,n507 ,n504);
    or g1955(n578 ,n505 ,n503);
    or g1956(n577 ,n28[6] ,n555);
    nor g1957(n576 ,n2240 ,n553);
    nor g1958(n575 ,n2239 ,n553);
    or g1959(n592 ,n148 ,n523);
    or g1960(n591 ,n27[2] ,n556);
    or g1961(n590 ,n148 ,n556);
    or g1962(n589 ,n27[2] ,n523);
    or g1963(n588 ,n1 ,n553);
    nor g1964(n587 ,n1 ,n554);
    nor g1965(n585 ,n1 ,n552);
    xnor g1966(n574 ,n4[14] ,n29[14]);
    xnor g1967(n573 ,n4[5] ,n29[5]);
    xnor g1968(n572 ,n4[4] ,n29[4]);
    xnor g1969(n571 ,n4[0] ,n29[0]);
    xnor g1970(n570 ,n4[6] ,n29[6]);
    xnor g1971(n569 ,n4[7] ,n29[7]);
    xnor g1972(n568 ,n4[2] ,n29[2]);
    xnor g1973(n567 ,n4[3] ,n29[3]);
    xnor g1974(n566 ,n4[11] ,n29[11]);
    xnor g1975(n565 ,n4[10] ,n29[10]);
    xnor g1976(n564 ,n4[8] ,n29[8]);
    xnor g1977(n563 ,n4[9] ,n29[9]);
    xnor g1978(n562 ,n4[13] ,n29[13]);
    xnor g1979(n561 ,n4[15] ,n29[15]);
    xnor g1980(n560 ,n4[12] ,n29[12]);
    xnor g1981(n559 ,n4[1] ,n29[1]);
    not g1982(n558 ,n557);
    not g1983(n555 ,n554);
    not g1984(n553 ,n552);
    nor g1985(n551 ,n135 ,n179);
    nor g1986(n550 ,n133 ,n183);
    nor g1987(n549 ,n136 ,n160);
    nor g1988(n548 ,n131 ,n171);
    nor g1989(n547 ,n134 ,n162);
    nor g1990(n546 ,n283 ,n1);
    nor g1991(n545 ,n365 ,n1);
    nor g1992(n544 ,n358 ,n1);
    nor g1993(n543 ,n393 ,n1);
    nor g1994(n542 ,n300 ,n1);
    nor g1995(n541 ,n208 ,n1);
    nor g1996(n540 ,n304 ,n1);
    nor g1997(n539 ,n303 ,n1);
    nor g1998(n557 ,n294 ,n1);
    nor g1999(n538 ,n223 ,n1);
    nor g2000(n537 ,n252 ,n1);
    nor g2001(n536 ,n360 ,n1);
    nor g2002(n535 ,n350 ,n1);
    nor g2003(n534 ,n281 ,n1);
    nor g2004(n533 ,n270 ,n1);
    nor g2005(n532 ,n204 ,n1);
    nor g2006(n531 ,n289 ,n1);
    or g2007(n556 ,n316 ,n27[6]);
    nor g2008(n530 ,n351 ,n1);
    nor g2009(n529 ,n344 ,n1);
    nor g2010(n528 ,n386 ,n1);
    nor g2011(n527 ,n302 ,n1);
    nor g2012(n526 ,n201 ,n1);
    nor g2013(n554 ,n292 ,n7);
    nor g2014(n552 ,n298 ,n6);
    not g2015(n525 ,n524);
    nor g2016(n518 ,n29[5] ,n2246);
    or g2017(n517 ,n26[13] ,n26[14]);
    nor g2018(n516 ,n29[7] ,n2244);
    or g2019(n515 ,n27[4] ,n27[5]);
    nor g2020(n514 ,n29[6] ,n2245);
    nor g2021(n513 ,n29[1] ,n2243);
    or g2022(n512 ,n138 ,n1);
    or g2023(n511 ,n137 ,n1);
    or g2024(n510 ,n28[4] ,n1);
    nor g2025(n509 ,n130 ,n29[1]);
    or g2026(n508 ,n26[5] ,n26[6]);
    or g2027(n507 ,n26[0] ,n26[1]);
    or g2028(n506 ,n26[7] ,n26[8]);
    or g2029(n505 ,n26[9] ,n26[10]);
    or g2030(n504 ,n26[2] ,n26[3]);
    or g2031(n503 ,n26[11] ,n26[12]);
    nor g2032(n502 ,n29[4] ,n2247);
    or g2033(n501 ,n28[5] ,n28[7]);
    nor g2034(n500 ,n27[0] ,n1);
    nor g2035(n499 ,n28[0] ,n1);
    nor g2036(n498 ,n26[0] ,n1);
    nor g2037(n524 ,n131 ,n1);
    or g2038(n523 ,n27[1] ,n27[6]);
    nor g2039(n497 ,n221 ,n1);
    nor g2040(n496 ,n305 ,n1);
    nor g2041(n495 ,n341 ,n1);
    or g2042(n522 ,n147 ,n308);
    or g2043(n521 ,n28[0] ,n28[3]);
    or g2044(n520 ,n147 ,n28[3]);
    or g2045(n519 ,n308 ,n28[0]);
    not g2046(n494 ,n21[11]);
    not g2047(n493 ,n23[0]);
    not g2048(n492 ,n20[15]);
    not g2049(n491 ,n18[10]);
    not g2050(n490 ,n9[5]);
    not g2051(n489 ,n21[12]);
    not g2052(n488 ,n8[9]);
    not g2053(n487 ,n21[5]);
    not g2054(n486 ,n15[14]);
    not g2055(n485 ,n10[2]);
    not g2056(n484 ,n9[10]);
    not g2057(n483 ,n8[5]);
    not g2058(n482 ,n13[12]);
    not g2059(n481 ,n8[3]);
    not g2060(n480 ,n8[6]);
    not g2061(n479 ,n13[6]);
    not g2062(n478 ,n23[9]);
    not g2063(n477 ,n23[11]);
    not g2064(n476 ,n11[8]);
    not g2065(n475 ,n11[7]);
    not g2066(n474 ,n14[8]);
    not g2067(n473 ,n10[10]);
    not g2068(n472 ,n18[3]);
    not g2069(n471 ,n16[2]);
    not g2070(n470 ,n5[13]);
    not g2071(n469 ,n19[14]);
    not g2072(n468 ,n9[2]);
    not g2073(n467 ,n19[11]);
    not g2074(n466 ,n18[11]);
    not g2075(n465 ,n23[12]);
    not g2076(n464 ,n22[13]);
    not g2077(n463 ,n23[3]);
    not g2078(n462 ,n19[7]);
    not g2079(n461 ,n9[15]);
    not g2080(n460 ,n12[10]);
    not g2081(n459 ,n11[15]);
    not g2082(n458 ,n14[6]);
    not g2083(n457 ,n18[15]);
    not g2084(n456 ,n22[10]);
    not g2085(n455 ,n5[3]);
    not g2086(n454 ,n17[10]);
    not g2087(n453 ,n15[1]);
    not g2088(n452 ,n22[4]);
    not g2089(n451 ,n10[12]);
    not g2090(n450 ,n11[11]);
    not g2091(n449 ,n21[3]);
    not g2092(n448 ,n5[12]);
    not g2093(n447 ,n15[10]);
    not g2094(n446 ,n5[1]);
    not g2095(n445 ,n8[7]);
    not g2096(n444 ,n5[8]);
    not g2097(n443 ,n9[4]);
    not g2098(n442 ,n13[11]);
    not g2099(n441 ,n22[11]);
    not g2100(n440 ,n10[8]);
    not g2101(n439 ,n9[7]);
    not g2102(n438 ,n10[3]);
    not g2103(n437 ,n10[9]);
    not g2104(n436 ,n12[14]);
    not g2105(n435 ,n5[6]);
    not g2106(n434 ,n15[12]);
    not g2107(n433 ,n8[13]);
    not g2108(n432 ,n13[9]);
    not g2109(n431 ,n16[8]);
    not g2110(n430 ,n20[8]);
    not g2111(n429 ,n15[7]);
    not g2112(n428 ,n9[8]);
    not g2113(n427 ,n10[7]);
    not g2114(n426 ,n12[0]);
    not g2115(n425 ,n20[4]);
    not g2116(n424 ,n5[4]);
    not g2117(n423 ,n5[0]);
    not g2118(n422 ,n12[9]);
    not g2119(n421 ,n15[6]);
    not g2120(n420 ,n11[2]);
    not g2121(n419 ,n8[0]);
    not g2122(n418 ,n19[4]);
    not g2123(n417 ,n17[13]);
    not g2124(n416 ,n10[6]);
    not g2125(n415 ,n19[6]);
    not g2126(n414 ,n15[13]);
    not g2127(n413 ,n11[9]);
    not g2128(n412 ,n17[12]);
    not g2129(n411 ,n23[8]);
    not g2130(n410 ,n18[14]);
    not g2131(n409 ,n9[12]);
    not g2132(n408 ,n18[1]);
    not g2133(n407 ,n14[1]);
    not g2134(n406 ,n16[6]);
    not g2135(n405 ,n21[13]);
    not g2136(n404 ,n19[9]);
    not g2137(n403 ,n22[12]);
    not g2138(n402 ,n13[15]);
    not g2139(n401 ,n23[14]);
    not g2140(n400 ,n14[2]);
    not g2141(n399 ,n17[14]);
    not g2142(n398 ,n16[5]);
    not g2143(n397 ,n22[0]);
    not g2144(n396 ,n21[14]);
    not g2145(n395 ,n16[9]);
    not g2146(n394 ,n18[4]);
    not g2147(n393 ,n24[7]);
    not g2148(n392 ,n22[5]);
    not g2149(n391 ,n12[12]);
    not g2150(n390 ,n17[15]);
    not g2151(n389 ,n11[12]);
    not g2152(n388 ,n5[2]);
    not g2153(n387 ,n15[4]);
    not g2154(n386 ,n24[5]);
    not g2155(n385 ,n8[12]);
    not g2156(n384 ,n15[0]);
    not g2157(n383 ,n19[12]);
    not g2158(n382 ,n14[10]);
    not g2159(n381 ,n23[13]);
    not g2160(n380 ,n19[10]);
    not g2161(n379 ,n17[5]);
    not g2162(n378 ,n17[9]);
    not g2163(n377 ,n22[9]);
    not g2164(n376 ,n5[9]);
    not g2165(n375 ,n11[4]);
    not g2166(n374 ,n20[12]);
    not g2167(n373 ,n11[5]);
    not g2168(n372 ,n11[0]);
    not g2169(n371 ,n5[7]);
    not g2170(n370 ,n20[11]);
    not g2171(n369 ,n20[10]);
    not g2172(n368 ,n9[1]);
    not g2173(n367 ,n18[6]);
    not g2174(n366 ,n14[0]);
    not g2175(n365 ,n24[6]);
    not g2176(n364 ,n8[10]);
    not g2177(n363 ,n21[1]);
    not g2178(n362 ,n8[11]);
    not g2179(n361 ,n20[13]);
    not g2180(n360 ,n24[3]);
    not g2181(n359 ,n23[15]);
    not g2182(n358 ,n24[2]);
    not g2183(n357 ,n12[8]);
    not g2184(n356 ,n17[1]);
    not g2185(n355 ,n14[13]);
    not g2186(n354 ,n20[9]);
    not g2187(n353 ,n15[5]);
    not g2188(n352 ,n14[15]);
    not g2189(n351 ,n25[1]);
    not g2190(n350 ,n25[3]);
    not g2191(n349 ,n16[11]);
    not g2192(n348 ,n13[5]);
    not g2193(n347 ,n13[10]);
    not g2194(n346 ,n17[4]);
    not g2195(n345 ,n14[12]);
    not g2196(n344 ,n24[1]);
    not g2197(n343 ,n22[1]);
    not g2198(n342 ,n14[9]);
    not g2199(n341 ,n25[7]);
    not g2200(n340 ,n21[10]);
    not g2201(n339 ,n10[5]);
    not g2202(n338 ,n9[14]);
    not g2203(n337 ,n23[10]);
    not g2204(n336 ,n22[2]);
    not g2205(n335 ,n11[6]);
    not g2206(n334 ,n5[5]);
    not g2207(n333 ,n12[4]);
    not g2208(n332 ,n12[5]);
    not g2209(n331 ,n21[7]);
    not g2210(n330 ,n13[3]);
    not g2211(n329 ,n18[9]);
    not g2212(n328 ,n10[15]);
    not g2213(n327 ,n16[13]);
    not g2214(n326 ,n15[2]);
    not g2215(n325 ,n16[10]);
    not g2216(n324 ,n18[13]);
    not g2217(n323 ,n21[4]);
    not g2218(n322 ,n11[13]);
    not g2219(n321 ,n14[14]);
    not g2220(n320 ,n18[5]);
    not g2221(n319 ,n14[11]);
    not g2222(n318 ,n26[9]);
    not g2223(n317 ,n26[2]);
    not g2224(n316 ,n27[1]);
    not g2225(n315 ,n26[4]);
    not g2226(n314 ,n26[3]);
    not g2227(n313 ,n26[12]);
    not g2228(n312 ,n26[14]);
    not g2229(n311 ,n26[13]);
    not g2230(n310 ,n28[1]);
    not g2231(n309 ,n27[0]);
    not g2232(n308 ,n28[3]);
    not g2233(n307 ,n28[2]);
    not g2234(n306 ,n27[3]);
    not g2235(n305 ,n2236);
    not g2236(n304 ,n2252);
    not g2237(n303 ,n2253);
    not g2238(n302 ,n2242);
    not g2239(n301 ,n2228);
    not g2240(n300 ,n2251);
    not g2241(n299 ,n2222);
    not g2242(n298 ,n3);
    not g2243(n297 ,n2233);
    not g2244(n296 ,n2221);
    not g2245(n295 ,n2230);
    not g2246(n294 ,n2241);
    not g2247(n293 ,n2229);
    not g2248(n292 ,n2);
    not g2249(n291 ,n2219);
    not g2250(n290 ,n2225);
    not g2251(n289 ,n2238);
    not g2252(n288 ,n2232);
    not g2253(n287 ,n2234);
    not g2254(n286 ,n2226);
    not g2255(n285 ,n2231);
    not g2256(n284 ,n2224);
    not g2257(n283 ,n2237);
    not g2258(n282 ,n2220);
    not g2259(n281 ,n2235);
    not g2260(n280 ,n2227);
    not g2261(n279 ,n2223);
    not g2262(n278 ,n21[2]);
    not g2263(n277 ,n5[14]);
    not g2264(n276 ,n23[2]);
    not g2265(n275 ,n9[13]);
    not g2266(n274 ,n12[2]);
    not g2267(n273 ,n11[3]);
    not g2268(n272 ,n20[14]);
    not g2269(n271 ,n18[2]);
    not g2270(n270 ,n25[2]);
    not g2271(n269 ,n20[3]);
    not g2272(n268 ,n13[7]);
    not g2273(n267 ,n11[10]);
    not g2274(n266 ,n23[1]);
    not g2275(n265 ,n8[1]);
    not g2276(n264 ,n15[9]);
    not g2277(n263 ,n5[15]);
    not g2278(n262 ,n10[11]);
    not g2279(n261 ,n17[8]);
    not g2280(n260 ,n10[14]);
    not g2281(n259 ,n8[15]);
    not g2282(n258 ,n23[5]);
    not g2283(n257 ,n5[11]);
    not g2284(n256 ,n18[12]);
    not g2285(n255 ,n16[0]);
    not g2286(n254 ,n12[13]);
    not g2287(n253 ,n16[15]);
    not g2288(n252 ,n25[4]);
    not g2289(n251 ,n23[7]);
    not g2290(n250 ,n22[7]);
    not g2291(n249 ,n15[15]);
    not g2292(n248 ,n20[1]);
    not g2293(n247 ,n17[6]);
    not g2294(n246 ,n20[6]);
    not g2295(n245 ,n16[4]);
    not g2296(n244 ,n18[0]);
    not g2297(n243 ,n21[0]);
    not g2298(n242 ,n12[11]);
    not g2299(n241 ,n15[3]);
    not g2300(n240 ,n21[15]);
    not g2301(n239 ,n10[13]);
    not g2302(n238 ,n10[1]);
    not g2303(n237 ,n13[14]);
    not g2304(n236 ,n16[1]);
    not g2305(n235 ,n8[4]);
    not g2306(n234 ,n8[14]);
    not g2307(n233 ,n13[1]);
    not g2308(n232 ,n19[3]);
    not g2309(n231 ,n2248);
    not g2310(n230 ,n14[7]);
    not g2311(n229 ,n12[15]);
    not g2312(n228 ,n18[8]);
    not g2313(n227 ,n14[3]);
    not g2314(n226 ,n9[11]);
    not g2315(n225 ,n12[3]);
    not g2316(n224 ,n8[8]);
    not g2317(n223 ,n24[4]);
    not g2318(n222 ,n16[3]);
    not g2319(n221 ,n25[5]);
    not g2320(n220 ,n9[3]);
    not g2321(n219 ,n19[0]);
    not g2322(n218 ,n8[2]);
    not g2323(n217 ,n11[1]);
    not g2324(n216 ,n13[8]);
    not g2325(n215 ,n21[9]);
    not g2326(n214 ,n12[6]);
    not g2327(n213 ,n9[6]);
    not g2328(n212 ,n19[5]);
    not g2329(n211 ,n22[6]);
    not g2330(n210 ,n16[14]);
    not g2331(n209 ,n16[12]);
    not g2332(n208 ,n25[0]);
    not g2333(n207 ,n9[0]);
    not g2334(n206 ,n12[1]);
    not g2335(n205 ,n12[7]);
    not g2336(n204 ,n24[0]);
    not g2337(n203 ,n13[0]);
    not g2338(n202 ,n16[7]);
    not g2339(n201 ,n25[6]);
    not g2340(n200 ,n19[1]);
    not g2341(n199 ,n21[8]);
    not g2342(n198 ,n23[4]);
    not g2343(n197 ,n13[2]);
    not g2344(n196 ,n11[14]);
    not g2345(n195 ,n18[7]);
    not g2346(n194 ,n19[2]);
    not g2347(n193 ,n22[8]);
    not g2348(n192 ,n19[8]);
    not g2349(n191 ,n20[5]);
    not g2350(n190 ,n22[14]);
    not g2351(n189 ,n22[15]);
    not g2352(n188 ,n20[0]);
    not g2353(n187 ,n14[4]);
    not g2354(n186 ,n10[4]);
    not g2355(n185 ,n13[13]);
    not g2356(n184 ,n21[6]);
    not g2357(n183 ,n2246);
    not g2358(n182 ,n13[4]);
    not g2359(n181 ,n20[7]);
    not g2360(n180 ,n22[3]);
    not g2361(n179 ,n2247);
    not g2362(n178 ,n15[8]);
    not g2363(n177 ,n17[7]);
    not g2364(n176 ,n17[0]);
    not g2365(n175 ,n17[11]);
    not g2366(n174 ,n17[3]);
    not g2367(n173 ,n2249);
    not g2368(n172 ,n20[2]);
    not g2369(n171 ,n2250);
    not g2370(n170 ,n10[0]);
    not g2371(n169 ,n15[11]);
    not g2372(n168 ,n2243);
    not g2373(n167 ,n2240);
    not g2374(n166 ,n14[5]);
    not g2375(n165 ,n23[6]);
    not g2376(n164 ,n2239);
    not g2377(n163 ,n9[9]);
    not g2378(n162 ,n2245);
    not g2379(n161 ,n19[13]);
    not g2380(n160 ,n2244);
    not g2381(n159 ,n17[2]);
    not g2382(n158 ,n19[15]);
    not g2383(n157 ,n5[10]);
    not g2384(n156 ,n26[8]);
    not g2385(n155 ,n26[6]);
    not g2386(n154 ,n26[1]);
    not g2387(n153 ,n26[5]);
    not g2388(n152 ,n26[10]);
    not g2389(n151 ,n26[15]);
    not g2390(n150 ,n26[7]);
    not g2391(n149 ,n26[11]);
    not g2392(n148 ,n27[2]);
    not g2393(n147 ,n28[0]);
    not g2394(n146 ,n29[14]);
    not g2395(n145 ,n29[13]);
    not g2396(n144 ,n29[12]);
    not g2397(n143 ,n29[15]);
    not g2398(n142 ,n29[10]);
    not g2399(n141 ,n29[8]);
    not g2400(n140 ,n29[9]);
    not g2401(n139 ,n29[11]);
    not g2402(n138 ,n29[3]);
    not g2403(n137 ,n29[2]);
    not g2404(n136 ,n29[7]);
    not g2405(n135 ,n29[4]);
    not g2406(n134 ,n29[6]);
    not g2407(n133 ,n29[5]);
    not g2408(n132 ,n29[0]);
    not g2409(n131 ,n29[1]);
    not g2410(n130 ,n1);
    xor g2411(n2226 ,n26[15] ,n57);
    xor g2412(n2225 ,n26[14] ,n55);
    nor g2413(n57 ,n26[14] ,n56);
    xor g2414(n2224 ,n26[13] ,n53);
    not g2415(n56 ,n55);
    nor g2416(n55 ,n26[13] ,n54);
    xor g2417(n2223 ,n26[12] ,n51);
    not g2418(n54 ,n53);
    nor g2419(n53 ,n26[12] ,n52);
    xor g2420(n2222 ,n26[11] ,n49);
    not g2421(n52 ,n51);
    nor g2422(n51 ,n26[11] ,n50);
    xor g2423(n2221 ,n26[10] ,n47);
    not g2424(n50 ,n49);
    nor g2425(n49 ,n26[10] ,n48);
    xor g2426(n2220 ,n26[9] ,n45);
    not g2427(n48 ,n47);
    nor g2428(n47 ,n26[9] ,n46);
    xor g2429(n2219 ,n26[8] ,n43);
    not g2430(n46 ,n45);
    nor g2431(n45 ,n26[8] ,n44);
    xor g2432(n2235 ,n26[7] ,n41);
    not g2433(n44 ,n43);
    nor g2434(n43 ,n26[7] ,n42);
    xor g2435(n2236 ,n26[6] ,n39);
    not g2436(n42 ,n41);
    nor g2437(n41 ,n26[6] ,n40);
    xor g2438(n2237 ,n26[5] ,n37);
    not g2439(n40 ,n39);
    nor g2440(n39 ,n26[5] ,n38);
    xor g2441(n2238 ,n26[4] ,n35);
    not g2442(n38 ,n37);
    nor g2443(n37 ,n26[4] ,n36);
    xor g2444(n2239 ,n26[3] ,n33);
    not g2445(n36 ,n35);
    nor g2446(n35 ,n26[3] ,n34);
    xor g2447(n2240 ,n26[2] ,n31);
    not g2448(n34 ,n33);
    nor g2449(n33 ,n26[2] ,n32);
    not g2450(n32 ,n31);
    nor g2451(n31 ,n26[1] ,n26[0]);
    xor g2452(n2234 ,n26[15] ,n113);
    nor g2453(n2233 ,n112 ,n113);
    nor g2454(n113 ,n69 ,n111);
    nor g2455(n112 ,n26[14] ,n110);
    nor g2456(n2232 ,n109 ,n110);
    not g2457(n111 ,n110);
    nor g2458(n110 ,n59 ,n108);
    nor g2459(n109 ,n26[13] ,n107);
    nor g2460(n2231 ,n106 ,n107);
    not g2461(n108 ,n107);
    nor g2462(n107 ,n72 ,n105);
    nor g2463(n106 ,n26[12] ,n104);
    nor g2464(n2230 ,n103 ,n104);
    not g2465(n105 ,n104);
    nor g2466(n104 ,n68 ,n102);
    nor g2467(n103 ,n26[11] ,n101);
    nor g2468(n2229 ,n100 ,n101);
    not g2469(n102 ,n101);
    nor g2470(n101 ,n70 ,n99);
    nor g2471(n100 ,n26[10] ,n98);
    nor g2472(n2228 ,n97 ,n98);
    not g2473(n99 ,n98);
    nor g2474(n98 ,n67 ,n96);
    nor g2475(n97 ,n26[9] ,n95);
    nor g2476(n2227 ,n94 ,n95);
    not g2477(n96 ,n95);
    nor g2478(n95 ,n64 ,n93);
    nor g2479(n94 ,n26[8] ,n92);
    nor g2480(n2244 ,n91 ,n92);
    not g2481(n93 ,n92);
    nor g2482(n92 ,n65 ,n90);
    nor g2483(n91 ,n26[7] ,n89);
    nor g2484(n2245 ,n88 ,n89);
    not g2485(n90 ,n89);
    nor g2486(n89 ,n58 ,n87);
    nor g2487(n88 ,n26[6] ,n86);
    nor g2488(n2246 ,n85 ,n86);
    not g2489(n87 ,n86);
    nor g2490(n86 ,n63 ,n84);
    nor g2491(n85 ,n26[5] ,n83);
    nor g2492(n2247 ,n82 ,n83);
    not g2493(n84 ,n83);
    nor g2494(n83 ,n61 ,n81);
    nor g2495(n82 ,n26[4] ,n80);
    nor g2496(n2248 ,n79 ,n80);
    not g2497(n81 ,n80);
    nor g2498(n80 ,n60 ,n78);
    nor g2499(n79 ,n26[3] ,n77);
    nor g2500(n2249 ,n76 ,n77);
    not g2501(n78 ,n77);
    nor g2502(n77 ,n62 ,n75);
    nor g2503(n76 ,n26[2] ,n74);
    nor g2504(n2250 ,n74 ,n73);
    not g2505(n75 ,n74);
    nor g2506(n74 ,n66 ,n71);
    nor g2507(n73 ,n26[1] ,n26[0]);
    not g2508(n72 ,n26[12]);
    not g2509(n71 ,n26[0]);
    not g2510(n70 ,n26[10]);
    not g2511(n69 ,n26[14]);
    not g2512(n68 ,n26[11]);
    not g2513(n67 ,n26[9]);
    not g2514(n66 ,n26[1]);
    not g2515(n65 ,n26[7]);
    not g2516(n64 ,n26[8]);
    not g2517(n63 ,n26[5]);
    not g2518(n62 ,n26[2]);
    not g2519(n61 ,n26[4]);
    not g2520(n60 ,n26[3]);
    not g2521(n59 ,n26[13]);
    not g2522(n58 ,n26[6]);
    xor g2523(n2251 ,n28[3] ,n121);
    nor g2524(n2252 ,n120 ,n121);
    nor g2525(n121 ,n116 ,n119);
    nor g2526(n120 ,n28[2] ,n118);
    nor g2527(n2253 ,n118 ,n117);
    not g2528(n119 ,n118);
    nor g2529(n118 ,n114 ,n115);
    nor g2530(n117 ,n28[1] ,n28[0]);
    not g2531(n116 ,n28[2]);
    not g2532(n115 ,n28[0]);
    not g2533(n114 ,n28[1]);
    xor g2534(n2241 ,n27[3] ,n129);
    nor g2535(n2242 ,n128 ,n129);
    nor g2536(n129 ,n124 ,n127);
    nor g2537(n128 ,n27[2] ,n126);
    nor g2538(n2243 ,n126 ,n125);
    not g2539(n127 ,n126);
    nor g2540(n126 ,n122 ,n123);
    nor g2541(n125 ,n27[1] ,n27[0]);
    not g2542(n124 ,n27[2]);
    not g2543(n123 ,n27[0]);
    not g2544(n122 ,n27[1]);
    xor g2545(n4580 ,n28[0] ,n27[0]);
    xor g2546(n4581 ,n28[1] ,n27[1]);
    or g2547(n29[4] ,n4561 ,n4571);
    or g2548(n29[9] ,n4549 ,n4570);
    or g2549(n29[10] ,n4537 ,n4563);
    or g2550(n29[3] ,n4540 ,n4565);
    or g2551(n29[8] ,n4545 ,n4568);
    or g2552(n29[2] ,n4544 ,n4567);
    or g2553(n29[7] ,n4541 ,n4569);
    or g2554(n29[1] ,n4542 ,n4566);
    or g2555(n29[6] ,n4536 ,n4562);
    or g2556(n29[0] ,n4547 ,n4564);
    or g2557(n29[5] ,n4533 ,n4572);
    or g2558(n29[14] ,n4484 ,n4546);
    or g2559(n29[12] ,n4534 ,n4550);
    or g2560(n29[13] ,n4500 ,n4538);
    or g2561(n29[15] ,n4519 ,n4535);
    or g2562(n29[11] ,n4543 ,n4539);
    or g2563(n4572 ,n4518 ,n4548);
    or g2564(n4571 ,n4513 ,n4560);
    or g2565(n4570 ,n4511 ,n4559);
    or g2566(n4569 ,n4492 ,n4553);
    or g2567(n4568 ,n4502 ,n4556);
    or g2568(n4567 ,n4504 ,n4557);
    or g2569(n4566 ,n4499 ,n4555);
    or g2570(n4565 ,n4508 ,n4558);
    or g2571(n4564 ,n4494 ,n4554);
    or g2572(n4563 ,n4521 ,n4551);
    or g2573(n4562 ,n4522 ,n4552);
    or g2574(n4561 ,n4503 ,n4514);
    nor g2575(n4560 ,n4467 ,n4480);
    nor g2576(n4559 ,n4459 ,n4478);
    nor g2577(n4558 ,n4462 ,n4477);
    nor g2578(n4557 ,n4468 ,n4476);
    nor g2579(n4556 ,n4464 ,n4479);
    nor g2580(n4555 ,n4466 ,n4475);
    nor g2581(n4554 ,n4463 ,n4474);
    nor g2582(n4553 ,n4461 ,n4473);
    nor g2583(n4552 ,n4460 ,n4472);
    nor g2584(n4551 ,n4465 ,n4482);
    or g2585(n4550 ,n4509 ,n4507);
    or g2586(n4549 ,n4515 ,n4531);
    nor g2587(n4548 ,n4469 ,n4481);
    or g2588(n4547 ,n4524 ,n4495);
    or g2589(n4546 ,n4512 ,n4532);
    or g2590(n4545 ,n4506 ,n4527);
    or g2591(n4544 ,n4528 ,n4505);
    or g2592(n4543 ,n4501 ,n4526);
    or g2593(n4542 ,n4510 ,n4525);
    or g2594(n4541 ,n4488 ,n4523);
    or g2595(n4540 ,n4497 ,n4529);
    or g2596(n4539 ,n4496 ,n4493);
    or g2597(n4538 ,n4491 ,n4485);
    or g2598(n4537 ,n4490 ,n4486);
    or g2599(n4536 ,n4489 ,n4487);
    or g2600(n4535 ,n4516 ,n4498);
    or g2601(n4534 ,n4517 ,n4530);
    or g2602(n4533 ,n4483 ,n4520);
    nor g2603(n4532 ,n4400 ,n4458);
    nor g2604(n4531 ,n4418 ,n4471);
    nor g2605(n4530 ,n4416 ,n4471);
    nor g2606(n4529 ,n4417 ,n4471);
    nor g2607(n4528 ,n4389 ,n4471);
    nor g2608(n4527 ,n4390 ,n4471);
    nor g2609(n4526 ,n4385 ,n4471);
    nor g2610(n4525 ,n4410 ,n4471);
    nor g2611(n4524 ,n4397 ,n4471);
    nor g2612(n4523 ,n4384 ,n4471);
    nor g2613(n4522 ,n4419 ,n4471);
    nor g2614(n4521 ,n4387 ,n4471);
    nor g2615(n4520 ,n4388 ,n4471);
    nor g2616(n4519 ,n4406 ,n4457);
    nor g2617(n4518 ,n4432 ,n4457);
    nor g2618(n4517 ,n4394 ,n4458);
    nor g2619(n4516 ,n4405 ,n4470);
    nor g2620(n4515 ,n4441 ,n4458);
    nor g2621(n4514 ,n4433 ,n4457);
    nor g2622(n4513 ,n4412 ,n4458);
    nor g2623(n4512 ,n4399 ,n4470);
    nor g2624(n4511 ,n4404 ,n4457);
    nor g2625(n4510 ,n4443 ,n4458);
    nor g2626(n4509 ,n4437 ,n4470);
    nor g2627(n4508 ,n4445 ,n4457);
    nor g2628(n4507 ,n4398 ,n4457);
    nor g2629(n4506 ,n4434 ,n4458);
    nor g2630(n4505 ,n4409 ,n4457);
    nor g2631(n4504 ,n4402 ,n4458);
    nor g2632(n4503 ,n4386 ,n4471);
    nor g2633(n4502 ,n4395 ,n4457);
    nor g2634(n4501 ,n4436 ,n4470);
    nor g2635(n4500 ,n4414 ,n4470);
    nor g2636(n4499 ,n4411 ,n4457);
    nor g2637(n4498 ,n4430 ,n4458);
    nor g2638(n4497 ,n4440 ,n4458);
    nor g2639(n4496 ,n4429 ,n4458);
    nor g2640(n4495 ,n4408 ,n4457);
    nor g2641(n4494 ,n4407 ,n4458);
    nor g2642(n4493 ,n4444 ,n4457);
    nor g2643(n4492 ,n4403 ,n4457);
    nor g2644(n4491 ,n4442 ,n4458);
    nor g2645(n4490 ,n4439 ,n4458);
    nor g2646(n4489 ,n4438 ,n4458);
    nor g2647(n4488 ,n4428 ,n4458);
    nor g2648(n4487 ,n4435 ,n4457);
    nor g2649(n4486 ,n4431 ,n4457);
    nor g2650(n4485 ,n4413 ,n4457);
    nor g2651(n4484 ,n4396 ,n4457);
    nor g2652(n4483 ,n4401 ,n4458);
    or g2653(n4482 ,n4470 ,n4451);
    or g2654(n4481 ,n4470 ,n4455);
    or g2655(n4480 ,n4470 ,n4453);
    or g2656(n4479 ,n4470 ,n4454);
    or g2657(n4478 ,n4470 ,n4452);
    or g2658(n4477 ,n4470 ,n4456);
    or g2659(n4476 ,n4470 ,n4450);
    or g2660(n4475 ,n4470 ,n4449);
    or g2661(n4474 ,n4470 ,n4448);
    or g2662(n4473 ,n4470 ,n4447);
    or g2663(n4472 ,n4470 ,n4446);
    nor g2664(n4469 ,n4393 ,n4384);
    nor g2665(n4468 ,n4423 ,n4386);
    nor g2666(n4467 ,n4391 ,n4419);
    nor g2667(n4466 ,n4422 ,n4417);
    nor g2668(n4465 ,n4392 ,n4416);
    nor g2669(n4464 ,n4425 ,n4387);
    nor g2670(n4463 ,n4421 ,n4389);
    nor g2671(n4462 ,n4427 ,n4388);
    nor g2672(n4461 ,n4426 ,n4418);
    nor g2673(n4460 ,n4424 ,n4390);
    nor g2674(n4459 ,n4420 ,n4385);
    or g2675(n4471 ,n4415 ,n3);
    or g2676(n4470 ,n4415 ,n4383);
    nor g2677(n4456 ,n4636 ,n30[5]);
    nor g2678(n4455 ,n4634 ,n30[7]);
    nor g2679(n4454 ,n4631 ,n30[10]);
    nor g2680(n4453 ,n4635 ,n30[6]);
    nor g2681(n4452 ,n4630 ,n30[11]);
    nor g2682(n4451 ,n4629 ,n30[12]);
    nor g2683(n4450 ,n4637 ,n30[4]);
    nor g2684(n4449 ,n4638 ,n30[3]);
    nor g2685(n4448 ,n4639 ,n30[2]);
    nor g2686(n4447 ,n4632 ,n30[9]);
    nor g2687(n4446 ,n4633 ,n30[8]);
    or g2688(n4458 ,n4383 ,n2);
    or g2689(n4457 ,n2 ,n3);
    not g2690(n4445 ,n4607);
    not g2691(n4444 ,n4615);
    not g2692(n4443 ,n4589);
    not g2693(n4442 ,n4601);
    not g2694(n4441 ,n4597);
    not g2695(n4440 ,n4591);
    not g2696(n4439 ,n4598);
    not g2697(n4438 ,n4594);
    not g2698(n4437 ,n4576);
    not g2699(n4436 ,n4575);
    not g2700(n4435 ,n4610);
    not g2701(n4434 ,n4596);
    not g2702(n4433 ,n4608);
    not g2703(n4432 ,n4609);
    not g2704(n4431 ,n4614);
    not g2705(n4430 ,n4603);
    not g2706(n4429 ,n4599);
    not g2707(n4428 ,n4595);
    not g2708(n4427 ,n4636);
    not g2709(n4426 ,n4632);
    not g2710(n4425 ,n4631);
    not g2711(n4424 ,n4633);
    not g2712(n4423 ,n4637);
    not g2713(n4422 ,n4638);
    not g2714(n4421 ,n4639);
    not g2715(n4420 ,n4630);
    not g2716(n4419 ,n30[6]);
    not g2717(n4418 ,n30[9]);
    not g2718(n4417 ,n30[3]);
    not g2719(n4416 ,n30[12]);
    not g2720(n4415 ,n2);
    not g2721(n4414 ,n4577);
    not g2722(n4413 ,n4617);
    not g2723(n4412 ,n4592);
    not g2724(n4411 ,n4605);
    not g2725(n4410 ,n4574);
    not g2726(n4409 ,n4606);
    not g2727(n4408 ,n4604);
    not g2728(n4407 ,n4588);
    not g2729(n4406 ,n4619);
    not g2730(n4405 ,n4579);
    not g2731(n4404 ,n4613);
    not g2732(n4403 ,n4611);
    not g2733(n4402 ,n4590);
    not g2734(n4401 ,n4593);
    not g2735(n4400 ,n4602);
    not g2736(n4399 ,n4578);
    not g2737(n4398 ,n4616);
    not g2738(n4397 ,n4573);
    not g2739(n4396 ,n4618);
    not g2740(n4395 ,n4612);
    not g2741(n4394 ,n4600);
    not g2742(n4393 ,n4634);
    not g2743(n4392 ,n4629);
    not g2744(n4391 ,n4635);
    not g2745(n4390 ,n30[8]);
    not g2746(n4389 ,n30[2]);
    not g2747(n4388 ,n30[5]);
    not g2748(n4387 ,n30[10]);
    not g2749(n4386 ,n30[4]);
    not g2750(n4385 ,n30[11]);
    not g2751(n4384 ,n30[7]);
    not g2752(n4383 ,n3);
    xor g2753(n4583 ,n28[3] ,n27[3]);
    xor g2754(n4584 ,n28[4] ,n27[4]);
    xor g2755(n4585 ,n28[5] ,n27[5]);
    xor g2756(n4586 ,n28[6] ,n27[6]);
    xor g2757(n4587 ,n28[7] ,n27[7]);
    xor g2758(n4582 ,n28[2] ,n27[2]);
    xnor g2759(n4619 ,n2774 ,n2824);
    nor g2760(n2824 ,n2782 ,n2823);
    xnor g2761(n4618 ,n2790 ,n2822);
    nor g2762(n2823 ,n2822 ,n2783);
    nor g2763(n2822 ,n2791 ,n2821);
    xnor g2764(n4617 ,n2804 ,n2820);
    nor g2765(n2821 ,n2820 ,n2797);
    nor g2766(n2820 ,n2819 ,n2805);
    xnor g2767(n4616 ,n2808 ,n2818);
    nor g2768(n2819 ,n2807 ,n2818);
    nor g2769(n2818 ,n2792 ,n2817);
    xnor g2770(n4615 ,n2803 ,n2816);
    nor g2771(n2817 ,n2816 ,n2798);
    nor g2772(n2816 ,n2796 ,n2815);
    xnor g2773(n4614 ,n2802 ,n2814);
    nor g2774(n2815 ,n2814 ,n2799);
    nor g2775(n2814 ,n2781 ,n2813);
    xnor g2776(n4613 ,n2789 ,n2812);
    nor g2777(n2813 ,n2785 ,n2812);
    nor g2778(n2812 ,n2811 ,n2768);
    xnor g2779(n4612 ,n2773 ,n2810);
    nor g2780(n2811 ,n2770 ,n2810);
    nor g2781(n2810 ,n2766 ,n2809);
    xnor g2782(n4611 ,n2772 ,n2806);
    nor g2783(n2809 ,n2765 ,n2806);
    xnor g2784(n2808 ,n2795 ,n2800);
    nor g2785(n2807 ,n2801 ,n2795);
    nor g2786(n2806 ,n2750 ,n2793);
    nor g2787(n2805 ,n2800 ,n2794);
    xnor g2788(n2804 ,n2776 ,n2786);
    xnor g2789(n2803 ,n2778 ,n2761);
    xnor g2790(n2802 ,n2779 ,n2751);
    xnor g2791(n4610 ,n2755 ,n2788);
    not g2792(n2801 ,n2800);
    nor g2793(n2799 ,n2752 ,n2779);
    nor g2794(n2798 ,n2762 ,n2778);
    nor g2795(n2797 ,n2787 ,n2776);
    nor g2796(n2796 ,n2751 ,n2780);
    nor g2797(n2800 ,n2771 ,n2784);
    not g2798(n2795 ,n2794);
    nor g2799(n2793 ,n2747 ,n2788);
    nor g2800(n2792 ,n2761 ,n2777);
    nor g2801(n2791 ,n2786 ,n2775);
    xnor g2802(n2790 ,n2764 ,n2757);
    xnor g2803(n2789 ,n2760 ,n2743);
    xnor g2804(n2794 ,n2754 ,n2711);
    not g2805(n2787 ,n2786);
    nor g2806(n2785 ,n2744 ,n2760);
    nor g2807(n2784 ,n2699 ,n2769);
    nor g2808(n2783 ,n2758 ,n2764);
    nor g2809(n2782 ,n2757 ,n2763);
    nor g2810(n2781 ,n2743 ,n2759);
    nor g2811(n2788 ,n2693 ,n2756);
    nor g2812(n2786 ,n2736 ,n2767);
    not g2813(n2780 ,n2779);
    not g2814(n2778 ,n2777);
    not g2815(n2776 ,n2775);
    xnor g2816(n4609 ,n2713 ,n2753);
    xnor g2817(n2774 ,n2714 ,n2745);
    xnor g2818(n2773 ,n2739 ,n2729);
    xnor g2819(n2772 ,n2738 ,n2731);
    xnor g2820(n2779 ,n2735 ,n2685);
    xnor g2821(n2777 ,n2733 ,n2741);
    xnor g2822(n2775 ,n2734 ,n2697);
    nor g2823(n2771 ,n2617 ,n2741);
    nor g2824(n2770 ,n2730 ,n2739);
    nor g2825(n2769 ,n2618 ,n2742);
    nor g2826(n2768 ,n2729 ,n2740);
    nor g2827(n2767 ,n2711 ,n2749);
    nor g2828(n2766 ,n2731 ,n2737);
    nor g2829(n2765 ,n2732 ,n2738);
    not g2830(n2764 ,n2763);
    not g2831(n2762 ,n2761);
    not g2832(n2760 ,n2759);
    not g2833(n2758 ,n2757);
    xnor g2834(n4608 ,n2715 ,n2700);
    nor g2835(n2756 ,n2710 ,n2753);
    xnor g2836(n2755 ,n2718 ,n2656);
    xnor g2837(n2754 ,n2720 ,n2613);
    xnor g2838(n2763 ,n2716 ,n2686);
    nor g2839(n2761 ,n2725 ,n2746);
    xnor g2840(n2759 ,n2712 ,n2666);
    nor g2841(n2757 ,n2727 ,n2748);
    not g2842(n2752 ,n2751);
    nor g2843(n2750 ,n2656 ,n2719);
    nor g2844(n2749 ,n2614 ,n2721);
    nor g2845(n2748 ,n2701 ,n2724);
    nor g2846(n2747 ,n2657 ,n2718);
    nor g2847(n2746 ,n2685 ,n2726);
    nor g2848(n2745 ,n2708 ,n2722);
    nor g2849(n2753 ,n2709 ,n2723);
    nor g2850(n2751 ,n2694 ,n2728);
    not g2851(n2744 ,n2743);
    not g2852(n2742 ,n2741);
    not g2853(n2740 ,n2739);
    not g2854(n2738 ,n2737);
    nor g2855(n2736 ,n2613 ,n2720);
    xnor g2856(n2735 ,n2695 ,n2672);
    xnor g2857(n2734 ,n2701 ,n2619);
    xnor g2858(n2733 ,n2699 ,n2617);
    nor g2859(n2743 ,n2705 ,n2717);
    xnor g2860(n2741 ,n2689 ,n2632);
    xnor g2861(n2739 ,n2690 ,n2664);
    xnor g2862(n2737 ,n2691 ,n2676);
    not g2863(n2732 ,n2731);
    not g2864(n2730 ,n2729);
    nor g2865(n2728 ,n2648 ,n2707);
    nor g2866(n2727 ,n2619 ,n2697);
    nor g2867(n2726 ,n2695 ,n2673);
    nor g2868(n2725 ,n2696 ,n2672);
    nor g2869(n2724 ,n2259 ,n2698);
    nor g2870(n2723 ,n2704 ,n2700);
    nor g2871(n2722 ,n2686 ,n2692);
    nor g2872(n2731 ,n2594 ,n2706);
    nor g2873(n2729 ,n2681 ,n2702);
    not g2874(n2721 ,n2720);
    not g2875(n2719 ,n2718);
    nor g2876(n2717 ,n2646 ,n2703);
    xnor g2877(n4607 ,n2662 ,n2645);
    xnor g2878(n2716 ,n2643 ,n2670);
    xnor g2879(n2715 ,n2674 ,n2596);
    xnor g2880(n2714 ,n2663 ,n2620);
    xnor g2881(n2713 ,n2684 ,n2654);
    xnor g2882(n2712 ,n2668 ,n2648);
    xnor g2883(n2720 ,n2661 ,n2598);
    xnor g2884(n2718 ,n2602 ,n2687);
    nor g2885(n2710 ,n2655 ,n2684);
    nor g2886(n2709 ,n2597 ,n2674);
    nor g2887(n2708 ,n2644 ,n2671);
    nor g2888(n2707 ,n2669 ,n2667);
    nor g2889(n2706 ,n2576 ,n2688);
    nor g2890(n2705 ,n2641 ,n2665);
    nor g2891(n2704 ,n2596 ,n2675);
    nor g2892(n2703 ,n2642 ,n2664);
    nor g2893(n2702 ,n2682 ,n2676);
    nor g2894(n2711 ,n2650 ,n2680);
    not g2895(n2698 ,n2697);
    not g2896(n2696 ,n2695);
    nor g2897(n2694 ,n2668 ,n2666);
    nor g2898(n2693 ,n2654 ,n2683);
    nor g2899(n2692 ,n2643 ,n2670);
    xnor g2900(n2691 ,n2658 ,n2261);
    xnor g2901(n2690 ,n2641 ,n2646);
    xnor g2902(n2689 ,n2333 ,n2660);
    xnor g2903(n2701 ,n2637 ,n2578);
    nor g2904(n2700 ,n2652 ,n2677);
    nor g2905(n2699 ,n2507 ,n2678);
    nor g2906(n2697 ,n2649 ,n2679);
    xnor g2907(n2695 ,n2516 ,n2647);
    not g2908(n2688 ,n2687);
    not g2909(n2684 ,n2683);
    nor g2910(n2682 ,n2582 ,n2659);
    nor g2911(n2681 ,n2261 ,n2658);
    nor g2912(n2680 ,n2651 ,n2660);
    nor g2913(n2679 ,n2598 ,n2640);
    nor g2914(n2678 ,n2506 ,n2647);
    nor g2915(n2677 ,n2645 ,n2638);
    xnor g2916(n2687 ,n2612 ,n2533);
    nor g2917(n2686 ,n2624 ,n2653);
    nor g2918(n2685 ,n2571 ,n2639);
    xnor g2919(n2683 ,n2609 ,n2260);
    not g2920(n2675 ,n2674);
    not g2921(n2673 ,n2672);
    not g2922(n2671 ,n2670);
    not g2923(n2669 ,n2668);
    not g2924(n2667 ,n2666);
    not g2925(n2665 ,n2664);
    xnor g2926(n4606 ,n2610 ,n2562);
    xnor g2927(n2663 ,n2566 ,n2621);
    xnor g2928(n2662 ,n2492 ,n2615);
    xnor g2929(n2661 ,n2634 ,n2580);
    xnor g2930(n2676 ,n2611 ,n2561);
    xnor g2931(n2674 ,n2607 ,n2522);
    xnor g2932(n2672 ,n2605 ,n2531);
    xnor g2933(n2670 ,n2606 ,n2462);
    xnor g2934(n2668 ,n2608 ,n2484);
    xnor g2935(n2666 ,n2604 ,n2636);
    xnor g2936(n2664 ,n2603 ,n2564);
    not g2937(n2659 ,n2658);
    not g2938(n2657 ,n2656);
    not g2939(n2655 ,n2654);
    nor g2940(n2653 ,n2601 ,n2625);
    nor g2941(n2652 ,n2492 ,n2616);
    nor g2942(n2651 ,n2332 ,n2633);
    nor g2943(n2650 ,n2333 ,n2632);
    nor g2944(n2649 ,n2581 ,n2635);
    nor g2945(n2660 ,n2577 ,n2631);
    nor g2946(n2658 ,n2593 ,n2627);
    nor g2947(n2656 ,n2574 ,n2623);
    nor g2948(n2654 ,n2583 ,n2626);
    not g2949(n2644 ,n2643);
    not g2950(n2642 ,n2641);
    nor g2951(n2640 ,n2580 ,n2634);
    nor g2952(n2639 ,n2636 ,n2592);
    nor g2953(n2638 ,n2491 ,n2615);
    xnor g2954(n2637 ,n2483 ,n2601);
    nor g2955(n2648 ,n2570 ,n2629);
    nor g2956(n2647 ,n2575 ,n2622);
    nor g2957(n2646 ,n2572 ,n2628);
    nor g2958(n2645 ,n2586 ,n2630);
    xnor g2959(n2643 ,n2483 ,n2599);
    xnor g2960(n2641 ,n2567 ,n2541);
    not g2961(n2635 ,n2634);
    not g2962(n2633 ,n2632);
    nor g2963(n2631 ,n2558 ,n2589);
    nor g2964(n2630 ,n2563 ,n2573);
    nor g2965(n2629 ,n2565 ,n2591);
    nor g2966(n2628 ,n2561 ,n2587);
    nor g2967(n2627 ,n2257 ,n2590);
    nor g2968(n2626 ,n2560 ,n2584);
    nor g2969(n2625 ,n2483 ,n2578);
    nor g2970(n2624 ,n2482 ,n2579);
    nor g2971(n2623 ,n2260 ,n2588);
    nor g2972(n2622 ,n2465 ,n2595);
    nor g2973(n2621 ,n2504 ,n2568);
    nor g2974(n2620 ,n2483 ,n2600);
    nor g2975(n2636 ,n2547 ,n2569);
    xnor g2976(n2634 ,n2346 ,n2542);
    nor g2977(n2632 ,n2585 ,n2598);
    not g2978(n2619 ,n2259);
    not g2979(n2618 ,n2617);
    not g2980(n2616 ,n2615);
    not g2981(n2614 ,n2613);
    xnor g2982(n2612 ,n2540 ,n2257);
    xnor g2983(n2611 ,n2519 ,n2536);
    xnor g2984(n2610 ,n2498 ,n2258);
    xnor g2985(n2609 ,n2529 ,n2528);
    xnor g2986(n2608 ,n2518 ,n2465);
    xnor g2987(n2607 ,n2490 ,n2560);
    xnor g2988(n2606 ,n2344 ,n2559);
    xnor g2989(n2605 ,n2558 ,n2538);
    xnor g2990(n2604 ,n2525 ,n2551);
    xnor g2991(n2603 ,n2523 ,n2549);
    xnor g2992(n2602 ,n2496 ,n2553);
    xnor g2993(n2617 ,n2556 ,n2464);
    xnor g2994(n2615 ,n2543 ,n2510);
    xnor g2995(n2613 ,n2555 ,n2488);
    not g2996(n2600 ,n2599);
    not g2997(n2597 ,n2596);
    nor g2998(n2595 ,n2485 ,n2517);
    nor g2999(n2594 ,n2495 ,n2554);
    nor g3000(n2593 ,n2539 ,n2533);
    nor g3001(n2592 ,n2552 ,n2526);
    nor g3002(n2591 ,n2550 ,n2524);
    nor g3003(n2590 ,n2540 ,n2534);
    nor g3004(n2589 ,n2537 ,n2532);
    nor g3005(n2588 ,n2527 ,n2530);
    nor g3006(n2587 ,n2535 ,n2520);
    nor g3007(n2586 ,n2497 ,n2548);
    nor g3008(n2585 ,n2515 ,n2544);
    nor g3009(n2584 ,n2489 ,n2521);
    nor g3010(n2583 ,n2490 ,n2522);
    or g3011(n2601 ,n2345 ,n2542);
    nor g3012(n2599 ,n2499 ,n2557);
    nor g3013(n2598 ,n2514 ,n2545);
    nor g3014(n2596 ,n2511 ,n2543);
    not g3015(n2582 ,n2261);
    not g3016(n2581 ,n2580);
    not g3017(n2579 ,n2578);
    nor g3018(n2577 ,n2538 ,n2531);
    nor g3019(n2576 ,n2496 ,n2553);
    nor g3020(n2575 ,n2484 ,n2518);
    nor g3021(n2574 ,n2528 ,n2529);
    xnor g3022(n4605 ,n2501 ,n2381);
    nor g3023(n2573 ,n2498 ,n2258);
    nor g3024(n2572 ,n2536 ,n2519);
    nor g3025(n2571 ,n2551 ,n2525);
    nor g3026(n2570 ,n2549 ,n2523);
    nor g3027(n2569 ,n2546 ,n2541);
    nor g3028(n2568 ,n2505 ,n2559);
    xnor g3029(n2567 ,n2494 ,n2406);
    xnor g3030(n2566 ,n2503 ,n2456);
    nor g3031(n2580 ,n2464 ,n2556);
    nor g3032(n2578 ,n2488 ,n2555);
    not g3033(n2565 ,n2564);
    not g3034(n2563 ,n2562);
    not g3035(n2554 ,n2553);
    not g3036(n2552 ,n2551);
    not g3037(n2550 ,n2549);
    not g3038(n2548 ,n2258);
    nor g3039(n2547 ,n2407 ,n2493);
    nor g3040(n2546 ,n2406 ,n2494);
    nor g3041(n2564 ,n2502 ,n2509);
    nor g3042(n2562 ,n2382 ,n2501);
    xnor g3043(n2561 ,n2342 ,n2477);
    xnor g3044(n2560 ,n2344 ,n2468);
    xnor g3045(n2559 ,n2342 ,n2450);
    xnor g3046(n2558 ,n2342 ,n2473);
    xnor g3047(n2557 ,n2342 ,n2481);
    xnor g3048(n2556 ,n2342 ,n2460);
    xnor g3049(n2555 ,n2342 ,n2471);
    nor g3050(n2553 ,n2500 ,n2513);
    xnor g3051(n2551 ,n2342 ,n2452);
    xnor g3052(n2549 ,n2342 ,n2455);
    not g3053(n2545 ,n2544);
    not g3054(n2540 ,n2539);
    not g3055(n2538 ,n2537);
    not g3056(n2536 ,n2535);
    not g3057(n2534 ,n2533);
    not g3058(n2532 ,n2531);
    not g3059(n2530 ,n2529);
    not g3060(n2528 ,n2527);
    not g3061(n2526 ,n2525);
    not g3062(n2524 ,n2523);
    not g3063(n2522 ,n2521);
    not g3064(n2520 ,n2519);
    not g3065(n2518 ,n2517);
    xnor g3066(n2544 ,n2344 ,n2461);
    xnor g3067(n2516 ,n2333 ,n2486);
    xnor g3068(n2543 ,n2346 ,n2472);
    xnor g3069(n2542 ,n2344 ,n2457);
    xnor g3070(n2541 ,n2346 ,n2454);
    xnor g3071(n2539 ,n2346 ,n2479);
    xnor g3072(n2537 ,n2345 ,n2476);
    xnor g3073(n2535 ,n2345 ,n2459);
    xnor g3074(n2533 ,n2475 ,n2344);
    xnor g3075(n2531 ,n2480 ,n2344);
    xnor g3076(n2529 ,n2469 ,n2344);
    xnor g3077(n2527 ,n2345 ,n2470);
    xnor g3078(n2525 ,n2458 ,n2344);
    xnor g3079(n2523 ,n2474 ,n2344);
    xnor g3080(n2521 ,n2345 ,n2478);
    xnor g3081(n2519 ,n2453 ,n2344);
    xnor g3082(n2517 ,n2345 ,n2451);
    not g3083(n2515 ,n2514);
    not g3084(n2513 ,n2512);
    not g3085(n2511 ,n2510);
    not g3086(n2509 ,n2508);
    nor g3087(n2507 ,n2332 ,n2486);
    nor g3088(n2506 ,n2333 ,n2487);
    nor g3089(n2505 ,n2344 ,n2463);
    nor g3090(n2504 ,n2343 ,n2462);
    xnor g3091(n2514 ,n2346 ,n2430);
    xnor g3092(n2503 ,n2342 ,n2431);
    nor g3093(n2512 ,n2344 ,n2468);
    nor g3094(n2510 ,n2346 ,n2467);
    nor g3095(n2508 ,n2342 ,n2466);
    not g3096(n2498 ,n2497);
    not g3097(n2496 ,n2495);
    not g3098(n2494 ,n2493);
    not g3099(n2492 ,n2491);
    not g3100(n2490 ,n2489);
    xnor g3101(n2502 ,n2332 ,n2415);
    xnor g3102(n2501 ,n2332 ,n2410);
    xnor g3103(n2500 ,n2332 ,n2409);
    xnor g3104(n2499 ,n2343 ,n2429);
    xnor g3105(n2497 ,n2332 ,n2412);
    xnor g3106(n2495 ,n2332 ,n2411);
    xnor g3107(n2493 ,n2332 ,n2408);
    xnor g3108(n2491 ,n2333 ,n2413);
    xnor g3109(n2489 ,n2333 ,n2414);
    not g3110(n2487 ,n2486);
    not g3111(n2485 ,n2484);
    not g3112(n2482 ,n2483);
    nor g3113(n2481 ,n2397 ,n2417);
    nor g3114(n2480 ,n2366 ,n2435);
    nor g3115(n2479 ,n2370 ,n2433);
    nor g3116(n2478 ,n2364 ,n2447);
    nor g3117(n2477 ,n2361 ,n2416);
    nor g3118(n2476 ,n2403 ,n2446);
    nor g3119(n2475 ,n2374 ,n2434);
    nor g3120(n2474 ,n2372 ,n2420);
    nor g3121(n2473 ,n2373 ,n2449);
    nor g3122(n2472 ,n2375 ,n2432);
    nor g3123(n2471 ,n2377 ,n2427);
    nor g3124(n2470 ,n2369 ,n2448);
    nor g3125(n2469 ,n2362 ,n2428);
    nor g3126(n2488 ,n2384 ,n2441);
    nor g3127(n2486 ,n2390 ,n2443);
    nor g3128(n2484 ,n2396 ,n2439);
    nor g3129(n2483 ,n2389 ,n2438);
    not g3130(n2463 ,n2462);
    nor g3131(n2461 ,n2399 ,n2419);
    nor g3132(n2460 ,n2368 ,n2436);
    nor g3133(n2459 ,n2371 ,n2424);
    nor g3134(n2458 ,n2360 ,n2426);
    nor g3135(n2457 ,n2393 ,n2444);
    nor g3136(n2456 ,n2400 ,n2442);
    nor g3137(n2455 ,n2367 ,n2421);
    nor g3138(n2454 ,n2363 ,n2423);
    nor g3139(n2453 ,n2376 ,n2422);
    nor g3140(n2452 ,n2365 ,n2418);
    nor g3141(n2451 ,n2398 ,n2425);
    nor g3142(n2450 ,n2402 ,n2445);
    xnor g3143(n2468 ,n2343 ,n2358);
    xnor g3144(n2467 ,n2345 ,n2359);
    xnor g3145(n2466 ,n2341 ,n2357);
    xnor g3146(n2465 ,n2333 ,n2383);
    nor g3147(n2464 ,n2386 ,n2440);
    nor g3148(n2462 ,n2395 ,n2437);
    nor g3149(n2449 ,n2272 ,n2378);
    nor g3150(n2448 ,n2265 ,n2380);
    nor g3151(n2447 ,n2262 ,n2380);
    nor g3152(n2446 ,n2275 ,n2380);
    nor g3153(n2445 ,n2275 ,n2378);
    nor g3154(n2444 ,n2275 ,n2379);
    nor g3155(n2443 ,n2262 ,n2405);
    nor g3156(n2442 ,n2264 ,n2405);
    nor g3157(n2441 ,n2272 ,n2405);
    nor g3158(n2440 ,n2265 ,n2405);
    nor g3159(n2439 ,n2274 ,n2405);
    nor g3160(n2438 ,n2263 ,n2405);
    nor g3161(n2437 ,n2273 ,n2405);
    nor g3162(n2436 ,n2263 ,n2378);
    nor g3163(n2435 ,n2273 ,n2379);
    nor g3164(n2434 ,n2262 ,n2379);
    nor g3165(n2433 ,n2272 ,n2380);
    nor g3166(n2432 ,n2274 ,n2380);
    nor g3167(n2431 ,n2276 ,n2378);
    nor g3168(n2430 ,n2276 ,n2380);
    nor g3169(n2429 ,n2276 ,n2379);
    nor g3170(n2428 ,n2274 ,n2379);
    nor g3171(n2427 ,n2273 ,n2378);
    nor g3172(n2426 ,n2263 ,n2379);
    nor g3173(n2425 ,n2264 ,n2380);
    nor g3174(n2424 ,n2263 ,n2380);
    nor g3175(n2423 ,n2273 ,n2380);
    nor g3176(n2422 ,n2265 ,n2379);
    nor g3177(n2421 ,n2262 ,n2378);
    nor g3178(n2420 ,n2272 ,n2379);
    nor g3179(n2419 ,n2264 ,n2379);
    nor g3180(n2418 ,n2265 ,n2378);
    nor g3181(n2417 ,n2264 ,n2378);
    nor g3182(n2416 ,n2274 ,n2378);
    xnor g3183(n4604 ,n2333 ,n2355);
    nor g3184(n2415 ,n2331 ,n2387);
    nor g3185(n2414 ,n2329 ,n2392);
    nor g3186(n2413 ,n2320 ,n2391);
    nor g3187(n2412 ,n2317 ,n2404);
    nor g3188(n2411 ,n2328 ,n2385);
    nor g3189(n2410 ,n2318 ,n2394);
    nor g3190(n2409 ,n2319 ,n2388);
    nor g3191(n2408 ,n2330 ,n2401);
    not g3192(n2407 ,n2406);
    nor g3193(n2404 ,n2262 ,n2356);
    nor g3194(n2403 ,n2276 ,n2352);
    nor g3195(n2402 ,n2276 ,n2354);
    nor g3196(n2401 ,n2275 ,n2356);
    nor g3197(n2400 ,n2275 ,n2348);
    nor g3198(n2399 ,n2275 ,n2350);
    nor g3199(n2398 ,n2275 ,n2352);
    nor g3200(n2397 ,n2275 ,n2354);
    nor g3201(n2396 ,n2262 ,n2348);
    nor g3202(n2395 ,n2264 ,n2348);
    nor g3203(n2394 ,n2274 ,n2356);
    nor g3204(n2393 ,n2276 ,n2350);
    nor g3205(n2392 ,n2272 ,n2356);
    nor g3206(n2391 ,n2265 ,n2356);
    nor g3207(n2390 ,n2265 ,n2348);
    nor g3208(n2389 ,n2273 ,n2348);
    nor g3209(n2388 ,n2263 ,n2356);
    nor g3210(n2387 ,n2264 ,n2356);
    nor g3211(n2386 ,n2272 ,n2348);
    nor g3212(n2385 ,n2273 ,n2356);
    nor g3213(n2384 ,n2263 ,n2348);
    nor g3214(n2383 ,n2276 ,n2356);
    nor g3215(n2406 ,n2274 ,n2348);
    or g3216(n2405 ,n2269 ,n2347);
    not g3217(n2382 ,n2381);
    nor g3218(n2377 ,n2264 ,n2354);
    nor g3219(n2376 ,n2272 ,n2350);
    nor g3220(n2375 ,n2262 ,n2352);
    nor g3221(n2374 ,n2265 ,n2350);
    nor g3222(n2373 ,n2263 ,n2354);
    nor g3223(n2372 ,n2263 ,n2350);
    nor g3224(n2371 ,n2273 ,n2352);
    nor g3225(n2370 ,n2263 ,n2352);
    nor g3226(n2369 ,n2272 ,n2352);
    nor g3227(n2368 ,n2273 ,n2354);
    nor g3228(n2367 ,n2265 ,n2354);
    nor g3229(n2366 ,n2264 ,n2350);
    nor g3230(n2365 ,n2272 ,n2354);
    nor g3231(n2364 ,n2265 ,n2352);
    nor g3232(n2363 ,n2264 ,n2352);
    nor g3233(n2362 ,n2262 ,n2350);
    nor g3234(n2361 ,n2262 ,n2354);
    nor g3235(n2360 ,n2273 ,n2350);
    nor g3236(n2359 ,n2274 ,n2352);
    nor g3237(n2358 ,n2274 ,n2350);
    nor g3238(n2357 ,n2274 ,n2354);
    nor g3239(n2381 ,n2332 ,n2355);
    or g3240(n2380 ,n2337 ,n2351);
    or g3241(n2379 ,n2340 ,n2349);
    or g3242(n2378 ,n2339 ,n2353);
    or g3243(n2356 ,n2307 ,n2338);
    xnor g3244(n2355 ,n2333 ,n2315);
    not g3245(n2354 ,n2353);
    xnor g3246(n2353 ,n2255 ,n2336);
    not g3247(n2352 ,n2351);
    xnor g3248(n2351 ,n2254 ,n2324);
    not g3249(n2350 ,n2349);
    xnor g3250(n2349 ,n2256 ,n2334);
    not g3251(n2348 ,n2347);
    xnor g3252(n2347 ,n2285 ,n2335);
    not g3253(n2345 ,n2346);
    xnor g3254(n2346 ,n2323 ,n2311);
    not g3255(n2343 ,n2344);
    xnor g3256(n2344 ,n2322 ,n2309);
    not g3257(n2341 ,n2342);
    xnor g3258(n2342 ,n2321 ,n2300);
    xnor g3259(n2340 ,n2326 ,n2309);
    xnor g3260(n2339 ,n2325 ,n2300);
    xnor g3261(n2338 ,n2316 ,n2313);
    xnor g3262(n2337 ,n2327 ,n2311);
    nor g3263(n2336 ,n2310 ,n2322);
    nor g3264(n2335 ,n2299 ,n2321);
    nor g3265(n2334 ,n2312 ,n2323);
    not g3266(n2332 ,n2333);
    xnor g3267(n2333 ,n2313 ,n2294);
    nor g3268(n2331 ,n2275 ,n2308);
    nor g3269(n2330 ,n2276 ,n2308);
    nor g3270(n2329 ,n2263 ,n2308);
    nor g3271(n2328 ,n2264 ,n2308);
    nor g3272(n2327 ,n2301 ,n2297);
    nor g3273(n2326 ,n2303 ,n2296);
    nor g3274(n2325 ,n2302 ,n2298);
    nor g3275(n2324 ,n2295 ,n2314);
    nor g3276(n2320 ,n2272 ,n2308);
    nor g3277(n2319 ,n2273 ,n2308);
    nor g3278(n2318 ,n2262 ,n2308);
    nor g3279(n2317 ,n2265 ,n2308);
    nor g3280(n2323 ,n2292 ,n2304);
    nor g3281(n2322 ,n2293 ,n2305);
    nor g3282(n2321 ,n2291 ,n2306);
    nor g3283(n2315 ,n2274 ,n2308);
    not g3284(n2314 ,n2313);
    not g3285(n2312 ,n2311);
    not g3286(n2310 ,n2309);
    not g3287(n2307 ,n2308);
    nor g3288(n2306 ,n2279 ,n2290);
    nor g3289(n2305 ,n2277 ,n2287);
    nor g3290(n2304 ,n2267 ,n2286);
    xnor g3291(n2313 ,n28[1] ,n27[1]);
    xnor g3292(n2311 ,n28[3] ,n27[3]);
    xnor g3293(n2309 ,n28[5] ,n27[5]);
    or g3294(n2308 ,n2294 ,n2288);
    not g3295(n2300 ,n2299);
    xnor g3296(n2298 ,n2279 ,n27[5]);
    xnor g3297(n2297 ,n2267 ,n27[1]);
    xnor g3298(n2296 ,n2277 ,n27[3]);
    xnor g3299(n2303 ,n2277 ,n28[4]);
    xnor g3300(n2302 ,n2279 ,n28[6]);
    xnor g3301(n2301 ,n2267 ,n28[2]);
    xnor g3302(n2299 ,n2269 ,n28[7]);
    not g3303(n2295 ,n2294);
    nor g3304(n2293 ,n2281 ,n2280);
    nor g3305(n2292 ,n2282 ,n2266);
    nor g3306(n2291 ,n2268 ,n2278);
    nor g3307(n2290 ,n28[6] ,n28[5]);
    nor g3308(n2289 ,n28[1] ,n27[1]);
    nor g3309(n2294 ,n2271 ,n2270);
    nor g3310(n2288 ,n28[0] ,n27[0]);
    nor g3311(n2287 ,n28[4] ,n28[3]);
    nor g3312(n2286 ,n28[2] ,n28[1]);
    nor g3313(n2285 ,n28[7] ,n27[7]);
    nor g3314(n2284 ,n28[5] ,n27[5]);
    nor g3315(n2283 ,n28[3] ,n27[3]);
    not g3316(n2282 ,n28[2]);
    not g3317(n2281 ,n28[4]);
    not g3318(n2280 ,n28[3]);
    not g3319(n2279 ,n27[6]);
    not g3320(n2278 ,n28[5]);
    not g3321(n2277 ,n27[4]);
    not g3322(n2276 ,n4628);
    not g3323(n2275 ,n4627);
    not g3324(n2274 ,n4620);
    not g3325(n2273 ,n4625);
    not g3326(n2272 ,n4623);
    not g3327(n2271 ,n28[0]);
    not g3328(n2270 ,n27[0]);
    not g3329(n2269 ,n27[7]);
    not g3330(n2268 ,n28[6]);
    not g3331(n2267 ,n27[2]);
    not g3332(n2266 ,n28[1]);
    not g3333(n2265 ,n4622);
    not g3334(n2264 ,n4626);
    not g3335(n2263 ,n4624);
    not g3336(n2262 ,n4621);
    xor g3337(n2261 ,n2502 ,n2508);
    xor g3338(n2260 ,n2512 ,n2500);
    xor g3339(n2259 ,n2499 ,n2557);
    xor g3340(n2258 ,n2346 ,n2467);
    xor g3341(n2257 ,n2341 ,n2466);
    xor g3342(n2256 ,n2283 ,n2303);
    xor g3343(n2255 ,n2284 ,n2302);
    xor g3344(n2254 ,n2289 ,n2301);
    or g3345(n30[12] ,n3115 ,n3176);
    xnor g3346(n30[11] ,n3121 ,n3175);
    nor g3347(n3176 ,n3117 ,n3175);
    nor g3348(n3175 ,n3147 ,n3174);
    xnor g3349(n30[10] ,n3153 ,n3173);
    nor g3350(n3174 ,n3146 ,n3173);
    nor g3351(n3173 ,n3155 ,n3172);
    xor g3352(n30[9] ,n3163 ,n3171);
    nor g3353(n3172 ,n3160 ,n3171);
    nor g3354(n3171 ,n3158 ,n3170);
    xnor g3355(n30[8] ,n3162 ,n3169);
    nor g3356(n3170 ,n3157 ,n3169);
    nor g3357(n3169 ,n3154 ,n3168);
    xor g3358(n30[7] ,n3161 ,n3167);
    nor g3359(n3168 ,n3159 ,n3167);
    nor g3360(n3167 ,n3138 ,n3166);
    xor g3361(n30[6] ,n3152 ,n3165);
    nor g3362(n3166 ,n3150 ,n3165);
    nor g3363(n3165 ,n3149 ,n3164);
    xnor g3364(n30[5] ,n3151 ,n3156);
    nor g3365(n3164 ,n3148 ,n3156);
    xnor g3366(n3163 ,n3139 ,n3130);
    xnor g3367(n3162 ,n3143 ,n3133);
    xnor g3368(n3161 ,n3141 ,n3128);
    xnor g3369(n30[4] ,n3137 ,n3132);
    nor g3370(n3160 ,n3131 ,n3140);
    nor g3371(n3159 ,n3129 ,n3142);
    nor g3372(n3158 ,n3133 ,n3144);
    nor g3373(n3157 ,n3134 ,n3143);
    nor g3374(n3156 ,n3136 ,n3145);
    nor g3375(n3155 ,n3130 ,n3139);
    nor g3376(n3154 ,n3128 ,n3141);
    xnor g3377(n3153 ,n3092 ,n3126);
    xnor g3378(n3152 ,n3124 ,n3109);
    xnor g3379(n3151 ,n3122 ,n3119);
    nor g3380(n3150 ,n3110 ,n3125);
    nor g3381(n3149 ,n3119 ,n3123);
    nor g3382(n3148 ,n3120 ,n3122);
    nor g3383(n3147 ,n3093 ,n3126);
    nor g3384(n3146 ,n3092 ,n3127);
    nor g3385(n3145 ,n3135 ,n3132);
    not g3386(n3144 ,n3143);
    not g3387(n3142 ,n3141);
    not g3388(n3140 ,n3139);
    nor g3389(n3138 ,n3109 ,n3124);
    xor g3390(n30[3] ,n3104 ,n3094);
    xnor g3391(n3137 ,n3111 ,n3080);
    xnor g3392(n3143 ,n3106 ,n3082);
    xnor g3393(n3141 ,n3105 ,n3083);
    xnor g3394(n3139 ,n3107 ,n3084);
    nor g3395(n3136 ,n3080 ,n3112);
    nor g3396(n3135 ,n3081 ,n3111);
    not g3397(n3134 ,n3133);
    nor g3398(n3133 ,n3087 ,n3114);
    nor g3399(n3132 ,n3097 ,n3113);
    not g3400(n3131 ,n3130);
    nor g3401(n3130 ,n3095 ,n3118);
    not g3402(n3129 ,n3128);
    nor g3403(n3128 ,n3091 ,n3108);
    not g3404(n3127 ,n3126);
    nor g3405(n3126 ,n3099 ,n3116);
    not g3406(n3125 ,n3124);
    xnor g3407(n3124 ,n3085 ,n3069);
    not g3408(n3123 ,n3122);
    xnor g3409(n3122 ,n3086 ,n3073);
    xnor g3410(n3121 ,n3102 ,n2897);
    not g3411(n3120 ,n3119);
    nor g3412(n3118 ,n3082 ,n3096);
    nor g3413(n3117 ,n2897 ,n3103);
    nor g3414(n3116 ,n3084 ,n3090);
    nor g3415(n3115 ,n2898 ,n3102);
    nor g3416(n3114 ,n3083 ,n3100);
    nor g3417(n3113 ,n3094 ,n3088);
    nor g3418(n3119 ,n3040 ,n3089);
    not g3419(n3112 ,n3111);
    not g3420(n3110 ,n3109);
    xor g3421(n30[2] ,n3062 ,n3018);
    nor g3422(n3108 ,n3055 ,n3098);
    xnor g3423(n3107 ,n3071 ,n3014);
    xnor g3424(n3106 ,n3067 ,n3041);
    xnor g3425(n3105 ,n3065 ,n3051);
    xnor g3426(n3104 ,n3063 ,n3016);
    xnor g3427(n3111 ,n3045 ,n3075);
    nor g3428(n3109 ,n3078 ,n3101);
    not g3429(n3103 ,n3102);
    nor g3430(n3101 ,n3074 ,n3079);
    nor g3431(n3100 ,n3052 ,n3066);
    nor g3432(n3099 ,n3015 ,n3072);
    nor g3433(n3098 ,n3054 ,n3070);
    nor g3434(n3097 ,n3017 ,n3064);
    nor g3435(n3096 ,n3042 ,n3067);
    nor g3436(n3095 ,n3041 ,n3068);
    nor g3437(n3102 ,n3005 ,n3076);
    not g3438(n3093 ,n3092);
    nor g3439(n3091 ,n3053 ,n3069);
    nor g3440(n3090 ,n3014 ,n3071);
    nor g3441(n3089 ,n3039 ,n3075);
    nor g3442(n3088 ,n3016 ,n3063);
    nor g3443(n3087 ,n3051 ,n3065);
    xnor g3444(n3086 ,n3049 ,n3047);
    xor g3445(n3085 ,n3054 ,n3055);
    nor g3446(n3094 ,n3058 ,n3077);
    xnor g3447(n3092 ,n3023 ,n3061);
    not g3448(n3081 ,n3080);
    nor g3449(n3079 ,n3048 ,n3050);
    nor g3450(n3078 ,n3047 ,n3049);
    nor g3451(n3077 ,n3019 ,n3057);
    nor g3452(n3076 ,n3006 ,n3061);
    nor g3453(n3084 ,n3001 ,n3060);
    nor g3454(n3083 ,n2998 ,n3056);
    nor g3455(n3082 ,n2995 ,n3046);
    nor g3456(n3080 ,n3000 ,n3059);
    not g3457(n3074 ,n3073);
    not g3458(n3072 ,n3071);
    not g3459(n3070 ,n3069);
    not g3460(n3068 ,n3067);
    not g3461(n3066 ,n3065);
    not g3462(n3064 ,n3063);
    xnor g3463(n3062 ,n3029 ,n2971);
    xnor g3464(n3075 ,n3025 ,n2962);
    xnor g3465(n3073 ,n3035 ,n2981);
    xnor g3466(n3071 ,n3026 ,n2983);
    xnor g3467(n3069 ,n3028 ,n3043);
    xnor g3468(n3067 ,n3022 ,n3031);
    xnor g3469(n3065 ,n3027 ,n3044);
    xnor g3470(n3063 ,n3024 ,n3033);
    nor g3471(n3060 ,n3011 ,n3032);
    nor g3472(n3059 ,n3007 ,n3034);
    nor g3473(n3058 ,n2971 ,n3030);
    nor g3474(n3057 ,n2972 ,n3029);
    nor g3475(n3056 ,n3012 ,n3043);
    nor g3476(n3061 ,n3013 ,n3037);
    not g3477(n3054 ,n3053);
    not g3478(n3052 ,n3051);
    not g3479(n3050 ,n3049);
    not g3480(n3048 ,n3047);
    nor g3481(n3046 ,n3009 ,n3044);
    xnor g3482(n3045 ,n3002 ,n3020);
    nor g3483(n3055 ,n2996 ,n3038);
    xnor g3484(n3053 ,n2990 ,n2984);
    xnor g3485(n3051 ,n2989 ,n2985);
    xnor g3486(n3049 ,n2991 ,n2964);
    nor g3487(n3047 ,n2994 ,n3036);
    not g3488(n3042 ,n3041);
    nor g3489(n3040 ,n3021 ,n3002);
    nor g3490(n3039 ,n3020 ,n3003);
    nor g3491(n3038 ,n2982 ,n3010);
    nor g3492(n3037 ,n2983 ,n3004);
    nor g3493(n4574 ,n3018 ,n2992);
    nor g3494(n3036 ,n2962 ,n3008);
    xnor g3495(n3035 ,n2958 ,n2944);
    nor g3496(n3044 ,n2967 ,n2993);
    nor g3497(n3043 ,n2968 ,n2999);
    nor g3498(n3041 ,n2966 ,n2997);
    not g3499(n3034 ,n3033);
    not g3500(n3032 ,n3031);
    not g3501(n3030 ,n3029);
    xnor g3502(n3028 ,n2946 ,n2979);
    xnor g3503(n3027 ,n2954 ,n2956);
    xnor g3504(n3026 ,n2899 ,n2950);
    xnor g3505(n3025 ,n2948 ,n2973);
    xnor g3506(n3024 ,n2960 ,n2952);
    xnor g3507(n3023 ,n2865 ,n2969);
    xnor g3508(n3022 ,n2975 ,n2977);
    xnor g3509(n3033 ,n2963 ,n2939);
    xnor g3510(n3031 ,n2901 ,n2965);
    xnor g3511(n3029 ,n2986 ,n2917);
    not g3512(n3021 ,n3020);
    not g3513(n3019 ,n3018);
    not g3514(n3017 ,n3016);
    not g3515(n3015 ,n3014);
    nor g3516(n3013 ,n2900 ,n2950);
    nor g3517(n3012 ,n2980 ,n2947);
    nor g3518(n3011 ,n2978 ,n2976);
    nor g3519(n3010 ,n2945 ,n2959);
    nor g3520(n3009 ,n2957 ,n2955);
    nor g3521(n3008 ,n2974 ,n2949);
    nor g3522(n3007 ,n2953 ,n2961);
    nor g3523(n3006 ,n2865 ,n2970);
    nor g3524(n3005 ,n2866 ,n2969);
    nor g3525(n3004 ,n2899 ,n2951);
    nor g3526(n3020 ,n2940 ,n2963);
    nor g3527(n3018 ,n2922 ,n2987);
    nor g3528(n3016 ,n2918 ,n2986);
    nor g3529(n3014 ,n2902 ,n2965);
    not g3530(n3003 ,n3002);
    nor g3531(n3001 ,n2977 ,n2975);
    nor g3532(n3000 ,n2952 ,n2960);
    nor g3533(n2999 ,n2943 ,n2964);
    nor g3534(n2998 ,n2979 ,n2946);
    nor g3535(n2997 ,n2942 ,n2985);
    nor g3536(n2996 ,n2944 ,n2958);
    nor g3537(n2995 ,n2956 ,n2954);
    nor g3538(n2994 ,n2973 ,n2948);
    nor g3539(n2993 ,n2941 ,n2984);
    nor g3540(n2992 ,n2921 ,n2988);
    xnor g3541(n2991 ,n2937 ,n2893);
    xnor g3542(n2990 ,n2913 ,n2891);
    xnor g3543(n2989 ,n2915 ,n2895);
    xnor g3544(n3002 ,n2875 ,n2919);
    not g3545(n2988 ,n2987);
    not g3546(n2982 ,n2981);
    not g3547(n2980 ,n2979);
    not g3548(n2978 ,n2977);
    not g3549(n2976 ,n2975);
    not g3550(n2974 ,n2973);
    not g3551(n2972 ,n2971);
    not g3552(n2970 ,n2969);
    nor g3553(n2968 ,n2894 ,n2938);
    nor g3554(n2967 ,n2892 ,n2914);
    nor g3555(n2966 ,n2896 ,n2916);
    nor g3556(n2987 ,n2877 ,n2929);
    nor g3557(n2986 ,n2880 ,n2927);
    nor g3558(n2985 ,n2857 ,n2923);
    nor g3559(n2984 ,n2885 ,n2934);
    nor g3560(n2983 ,n2888 ,n2925);
    nor g3561(n2981 ,n2876 ,n2920);
    nor g3562(n2979 ,n2882 ,n2909);
    nor g3563(n2977 ,n2878 ,n2928);
    nor g3564(n2975 ,n2861 ,n2907);
    nor g3565(n2973 ,n2890 ,n2926);
    nor g3566(n2971 ,n2859 ,n2911);
    nor g3567(n2969 ,n2889 ,n2935);
    not g3568(n2961 ,n2960);
    not g3569(n2959 ,n2958);
    not g3570(n2957 ,n2956);
    not g3571(n2955 ,n2954);
    not g3572(n2953 ,n2952);
    not g3573(n2951 ,n2950);
    not g3574(n2949 ,n2948);
    not g3575(n2947 ,n2946);
    not g3576(n2945 ,n2944);
    nor g3577(n2943 ,n2893 ,n2937);
    nor g3578(n2942 ,n2895 ,n2915);
    nor g3579(n2941 ,n2891 ,n2913);
    nor g3580(n2965 ,n2884 ,n2906);
    nor g3581(n2964 ,n2887 ,n2933);
    nor g3582(n2963 ,n2883 ,n2936);
    nor g3583(n2962 ,n2862 ,n2932);
    nor g3584(n2960 ,n2863 ,n2931);
    nor g3585(n2958 ,n2864 ,n2905);
    nor g3586(n2956 ,n2855 ,n2904);
    nor g3587(n2954 ,n2858 ,n2910);
    nor g3588(n2952 ,n2886 ,n2924);
    nor g3589(n2950 ,n2860 ,n2903);
    nor g3590(n2948 ,n2879 ,n2908);
    nor g3591(n2946 ,n2856 ,n2930);
    nor g3592(n2944 ,n2881 ,n2912);
    not g3593(n2940 ,n2939);
    not g3594(n2938 ,n2937);
    nor g3595(n2936 ,n2836 ,n2869);
    nor g3596(n2935 ,n2836 ,n2870);
    nor g3597(n2934 ,n2836 ,n2867);
    nor g3598(n2933 ,n2836 ,n2868);
    nor g3599(n2932 ,n2838 ,n2867);
    nor g3600(n2931 ,n2837 ,n2873);
    nor g3601(n2930 ,n2837 ,n2874);
    nor g3602(n2929 ,n2838 ,n2869);
    nor g3603(n2928 ,n2838 ,n2870);
    nor g3604(n2927 ,n2838 ,n2873);
    nor g3605(n2926 ,n2837 ,n2868);
    nor g3606(n2925 ,n2837 ,n2870);
    nor g3607(n2924 ,n2838 ,n2868);
    nor g3608(n2923 ,n2836 ,n2874);
    nor g3609(n2939 ,n2835 ,n2867);
    nor g3610(n2937 ,n2835 ,n2871);
    not g3611(n2922 ,n2921);
    not g3612(n2920 ,n2919);
    not g3613(n2918 ,n2917);
    not g3614(n2916 ,n2915);
    not g3615(n2914 ,n2913);
    nor g3616(n2912 ,n2838 ,n2874);
    nor g3617(n2911 ,n2837 ,n2869);
    nor g3618(n4573 ,n2835 ,n2869);
    nor g3619(n2910 ,n2837 ,n2871);
    nor g3620(n2909 ,n2838 ,n2871);
    nor g3621(n2908 ,n2836 ,n2873);
    nor g3622(n2907 ,n2837 ,n2872);
    nor g3623(n2906 ,n2836 ,n2871);
    nor g3624(n2905 ,n2837 ,n2867);
    nor g3625(n2904 ,n2838 ,n2872);
    nor g3626(n2903 ,n2836 ,n2872);
    nor g3627(n2921 ,n2835 ,n2873);
    nor g3628(n2919 ,n2835 ,n2874);
    nor g3629(n2917 ,n2835 ,n2868);
    nor g3630(n2915 ,n2835 ,n2870);
    nor g3631(n2913 ,n2835 ,n2872);
    not g3632(n2902 ,n2901);
    not g3633(n2900 ,n2899);
    not g3634(n2898 ,n2897);
    not g3635(n2896 ,n2895);
    not g3636(n2894 ,n2893);
    not g3637(n2892 ,n2891);
    nor g3638(n2890 ,n2838 ,n2848);
    nor g3639(n2889 ,n2837 ,n2851);
    nor g3640(n2888 ,n2838 ,n2851);
    nor g3641(n2887 ,n2837 ,n2848);
    nor g3642(n2886 ,n2835 ,n2848);
    nor g3643(n2885 ,n2837 ,n2847);
    nor g3644(n2884 ,n2837 ,n2850);
    nor g3645(n2883 ,n2837 ,n2852);
    nor g3646(n2882 ,n2835 ,n2850);
    nor g3647(n2881 ,n2835 ,n2849);
    nor g3648(n2880 ,n2835 ,n2846);
    nor g3649(n2879 ,n2837 ,n2846);
    nor g3650(n2878 ,n2835 ,n2851);
    nor g3651(n2877 ,n2835 ,n2852);
    nor g3652(n2901 ,n2836 ,n2849);
    nor g3653(n2899 ,n2836 ,n2850);
    nor g3654(n2897 ,n2836 ,n2851);
    nor g3655(n2895 ,n2836 ,n2847);
    nor g3656(n2893 ,n2836 ,n2846);
    nor g3657(n2891 ,n2836 ,n2848);
    not g3658(n2876 ,n2875);
    not g3659(n2866 ,n2865);
    nor g3660(n2864 ,n2838 ,n2847);
    nor g3661(n2863 ,n2838 ,n2846);
    nor g3662(n2862 ,n2835 ,n2847);
    nor g3663(n2861 ,n2838 ,n2854);
    nor g3664(n2860 ,n2837 ,n2854);
    nor g3665(n2859 ,n2838 ,n2852);
    nor g3666(n2858 ,n2838 ,n2850);
    nor g3667(n2857 ,n2837 ,n2849);
    nor g3668(n2856 ,n2838 ,n2849);
    nor g3669(n2855 ,n2835 ,n2854);
    nor g3670(n2875 ,n2836 ,n2852);
    xnor g3671(n2874 ,n4584 ,n4[4]);
    xnor g3672(n2873 ,n4581 ,n4[1]);
    or g3673(n2872 ,n2853 ,n2845);
    xnor g3674(n2871 ,n4585 ,n4[5]);
    xnor g3675(n2870 ,n4587 ,n4[7]);
    xnor g3676(n2869 ,n4580 ,n4[0]);
    xnor g3677(n2868 ,n4582 ,n4[2]);
    xnor g3678(n2867 ,n4583 ,n4[3]);
    nor g3679(n2865 ,n2836 ,n2854);
    not g3680(n2854 ,n2853);
    nor g3681(n2853 ,n2839 ,n2828);
    or g3682(n2852 ,n2832 ,n2834);
    or g3683(n2851 ,n2826 ,n2833);
    or g3684(n2850 ,n2842 ,n2827);
    or g3685(n2849 ,n2844 ,n2840);
    or g3686(n2848 ,n2830 ,n2831);
    or g3687(n2847 ,n2829 ,n2843);
    or g3688(n2846 ,n2825 ,n2841);
    nor g3689(n2845 ,n4586 ,n4[6]);
    not g3690(n2844 ,n4584);
    not g3691(n2843 ,n4[3]);
    not g3692(n2842 ,n4585);
    not g3693(n2841 ,n4[1]);
    not g3694(n2840 ,n4[4]);
    not g3695(n2839 ,n4586);
    not g3696(n2838 ,n5[1]);
    not g3697(n2837 ,n5[2]);
    not g3698(n2836 ,n5[3]);
    not g3699(n2835 ,n5[0]);
    not g3700(n2834 ,n4[0]);
    not g3701(n2833 ,n4[7]);
    not g3702(n2832 ,n4580);
    not g3703(n2831 ,n4[2]);
    not g3704(n2830 ,n4582);
    not g3705(n2829 ,n4583);
    not g3706(n2828 ,n4[6]);
    not g3707(n2827 ,n4[5]);
    not g3708(n2826 ,n4587);
    not g3709(n2825 ,n4581);
    xor g3710(n4603 ,n4156 ,n4271);
    nor g3711(n4271 ,n4177 ,n4270);
    xor g3712(n4602 ,n4198 ,n4269);
    nor g3713(n4270 ,n4195 ,n4269);
    nor g3714(n4269 ,n4217 ,n4268);
    xor g3715(n4601 ,n4232 ,n4267);
    nor g3716(n4268 ,n4267 ,n4231);
    nor g3717(n4267 ,n4240 ,n4266);
    xor g3718(n4600 ,n4246 ,n4265);
    nor g3719(n4266 ,n4265 ,n4241);
    nor g3720(n4265 ,n4264 ,n4248);
    xor g3721(n4599 ,n4256 ,n4263);
    nor g3722(n4264 ,n4263 ,n4253);
    nor g3723(n4263 ,n4252 ,n4262);
    xnor g3724(n4598 ,n4255 ,n4261);
    nor g3725(n4262 ,n4261 ,n4250);
    nor g3726(n4261 ,n4260 ,n4251);
    xnor g3727(n4597 ,n4254 ,n4259);
    nor g3728(n4260 ,n4249 ,n4259);
    nor g3729(n4259 ,n4258 ,n4242);
    xnor g3730(n4596 ,n4245 ,n4257);
    nor g3731(n4258 ,n4243 ,n4257);
    nor g3732(n4257 ,n4230 ,n4247);
    xnor g3733(n4256 ,n4238 ,n4224);
    xnor g3734(n4255 ,n4236 ,n4227);
    xnor g3735(n4254 ,n4234 ,n4220);
    xnor g3736(n4595 ,n4233 ,n4244);
    nor g3737(n4253 ,n4225 ,n4239);
    nor g3738(n4252 ,n4227 ,n4237);
    nor g3739(n4251 ,n4220 ,n4235);
    nor g3740(n4250 ,n4228 ,n4236);
    nor g3741(n4249 ,n4221 ,n4234);
    nor g3742(n4248 ,n4224 ,n4238);
    nor g3743(n4247 ,n4229 ,n4244);
    xnor g3744(n4246 ,n4222 ,n4202);
    xnor g3745(n4245 ,n4206 ,n4218);
    nor g3746(n4243 ,n4219 ,n4206);
    nor g3747(n4242 ,n4218 ,n4207);
    nor g3748(n4241 ,n4203 ,n4223);
    nor g3749(n4240 ,n4202 ,n4222);
    nor g3750(n4244 ,n4182 ,n4226);
    not g3751(n4239 ,n4238);
    not g3752(n4237 ,n4236);
    not g3753(n4235 ,n4234);
    xnor g3754(n4594 ,n4201 ,n4216);
    xnor g3755(n4233 ,n4204 ,n4168);
    xnor g3756(n4232 ,n4183 ,n4214);
    xnor g3757(n4238 ,n4208 ,n4185);
    xnor g3758(n4236 ,n4200 ,n4176);
    xnor g3759(n4234 ,n4199 ,n4186);
    nor g3760(n4231 ,n4184 ,n4215);
    nor g3761(n4230 ,n4168 ,n4205);
    nor g3762(n4229 ,n4169 ,n4204);
    not g3763(n4228 ,n4227);
    nor g3764(n4227 ,n4180 ,n4209);
    nor g3765(n4226 ,n4194 ,n4216);
    not g3766(n4225 ,n4224);
    nor g3767(n4224 ,n4193 ,n4211);
    not g3768(n4223 ,n4222);
    nor g3769(n4222 ,n4178 ,n4212);
    not g3770(n4221 ,n4220);
    nor g3771(n4220 ,n4191 ,n4210);
    not g3772(n4219 ,n4218);
    nor g3773(n4218 ,n4189 ,n4213);
    nor g3774(n4217 ,n4183 ,n4214);
    not g3775(n4215 ,n4214);
    nor g3776(n4213 ,n4091 ,n4188);
    nor g3777(n4212 ,n4185 ,n4197);
    nor g3778(n4211 ,n4176 ,n4192);
    nor g3779(n4210 ,n4135 ,n4190);
    nor g3780(n4209 ,n4196 ,n4187);
    xnor g3781(n4208 ,n4159 ,n4097);
    nor g3782(n4216 ,n4150 ,n4179);
    nor g3783(n4214 ,n4144 ,n4181);
    not g3784(n4207 ,n4206);
    not g3785(n4205 ,n4204);
    not g3786(n4203 ,n4202);
    xnor g3787(n4593 ,n4155 ,n4174);
    xnor g3788(n4201 ,n4166 ,n4108);
    xnor g3789(n4200 ,n4161 ,n4133);
    xnor g3790(n4199 ,n4118 ,n4172);
    xnor g3791(n4198 ,n4116 ,n4170);
    xnor g3792(n4206 ,n4153 ,n4157);
    xnor g3793(n4204 ,n4137 ,n4163);
    xnor g3794(n4202 ,n4154 ,n4175);
    nor g3795(n4197 ,n4098 ,n4160);
    nor g3796(n4196 ,n4119 ,n4173);
    nor g3797(n4195 ,n4117 ,n4171);
    nor g3798(n4194 ,n4109 ,n4166);
    nor g3799(n4193 ,n4133 ,n4162);
    nor g3800(n4192 ,n4134 ,n4161);
    nor g3801(n4191 ,n4107 ,n4157);
    nor g3802(n4190 ,n4106 ,n4158);
    nor g3803(n4189 ,n4080 ,n4163);
    nor g3804(n4188 ,n4079 ,n4164);
    not g3805(n4187 ,n4186);
    not g3806(n4184 ,n4183);
    nor g3807(n4182 ,n4108 ,n4167);
    nor g3808(n4181 ,n4148 ,n4175);
    nor g3809(n4180 ,n4118 ,n4172);
    nor g3810(n4179 ,n4149 ,n4174);
    nor g3811(n4178 ,n4097 ,n4159);
    nor g3812(n4177 ,n4116 ,n4170);
    xnor g3813(n4592 ,n4140 ,n4100);
    xnor g3814(n4186 ,n4139 ,n4099);
    nor g3815(n4185 ,n4152 ,n4165);
    xnor g3816(n4183 ,n4138 ,n4136);
    not g3817(n4173 ,n4172);
    not g3818(n4171 ,n4170);
    not g3819(n4169 ,n4168);
    not g3820(n4167 ,n4166);
    nor g3821(n4165 ,n4058 ,n4151);
    nor g3822(n4176 ,n4127 ,n4142);
    nor g3823(n4175 ,n4131 ,n4141);
    nor g3824(n4174 ,n4129 ,n4146);
    nor g3825(n4172 ,n4124 ,n4145);
    nor g3826(n4170 ,n4132 ,n4143);
    nor g3827(n4168 ,n4077 ,n4147);
    xnor g3828(n4166 ,n4102 ,n4120);
    not g3829(n4164 ,n4163);
    not g3830(n4162 ,n4161);
    not g3831(n4160 ,n4159);
    not g3832(n4158 ,n4157);
    xnor g3833(n4156 ,n4122 ,n3797);
    xnor g3834(n4155 ,n4112 ,n4071);
    xnor g3835(n4154 ,n4114 ,n4046);
    xnor g3836(n4153 ,n4106 ,n4135);
    xnor g3837(n4163 ,n4104 ,n4020);
    xnor g3838(n4161 ,n4101 ,n4110);
    xnor g3839(n4159 ,n4105 ,n4087);
    xnor g3840(n4157 ,n4103 ,n4083);
    nor g3841(n4152 ,n4050 ,n4111);
    nor g3842(n4151 ,n4051 ,n4110);
    nor g3843(n4150 ,n4071 ,n4113);
    nor g3844(n4149 ,n4072 ,n4112);
    nor g3845(n4148 ,n4047 ,n4115);
    nor g3846(n4147 ,n4096 ,n4121);
    nor g3847(n4146 ,n4100 ,n4128);
    nor g3848(n4145 ,n4022 ,n4130);
    nor g3849(n4144 ,n4046 ,n4114);
    nor g3850(n4143 ,n4125 ,n4136);
    nor g3851(n4142 ,n4099 ,n4126);
    nor g3852(n4141 ,n4076 ,n4123);
    xnor g3853(n4140 ,n4089 ,n3999);
    xnor g3854(n4139 ,n4048 ,n4081);
    xnor g3855(n4138 ,n4085 ,n4069);
    xnor g3856(n4137 ,n4079 ,n4091);
    not g3857(n4134 ,n4133);
    nor g3858(n4132 ,n4069 ,n4085);
    nor g3859(n4131 ,n4019 ,n4088);
    nor g3860(n4130 ,n4068 ,n4084);
    nor g3861(n4129 ,n3999 ,n4090);
    nor g3862(n4128 ,n4000 ,n4089);
    nor g3863(n4127 ,n4049 ,n4081);
    nor g3864(n4126 ,n4048 ,n4082);
    nor g3865(n4125 ,n4070 ,n4086);
    nor g3866(n4124 ,n4067 ,n4083);
    nor g3867(n4123 ,n4018 ,n4087);
    nor g3868(n4122 ,n3934 ,n4078);
    nor g3869(n4136 ,n4063 ,n4095);
    nor g3870(n4135 ,n4061 ,n4093);
    nor g3871(n4133 ,n4012 ,n4092);
    not g3872(n4121 ,n4120);
    not g3873(n4119 ,n4118);
    not g3874(n4117 ,n4116);
    not g3875(n4115 ,n4114);
    not g3876(n4113 ,n4112);
    not g3877(n4111 ,n4110);
    not g3878(n4109 ,n4108);
    not g3879(n4107 ,n4106);
    xnor g3880(n4591 ,n4039 ,n4038);
    xnor g3881(n4105 ,n4018 ,n4076);
    xnor g3882(n4104 ,n3964 ,n4074);
    xnor g3883(n4103 ,n4067 ,n4022);
    xnor g3884(n4102 ,n4052 ,n4054);
    xnor g3885(n4101 ,n4050 ,n4058);
    xnor g3886(n4120 ,n4045 ,n3922);
    xnor g3887(n4118 ,n4040 ,n4073);
    xnor g3888(n4116 ,n3956 ,n4075);
    xnor g3889(n4114 ,n4041 ,n4016);
    xnor g3890(n4112 ,n4042 ,n4056);
    xnor g3891(n4110 ,n4044 ,n3976);
    nor g3892(n4108 ,n4014 ,n4094);
    xnor g3893(n4106 ,n4043 ,n3977);
    not g3894(n4098 ,n4097);
    nor g3895(n4096 ,n4055 ,n4053);
    nor g3896(n4095 ,n3979 ,n4060);
    nor g3897(n4094 ,n4023 ,n4057);
    nor g3898(n4093 ,n4074 ,n4062);
    nor g3899(n4092 ,n4036 ,n4073);
    nor g3900(n4100 ,n4028 ,n4064);
    nor g3901(n4099 ,n4034 ,n4066);
    nor g3902(n4097 ,n4032 ,n4059);
    not g3903(n4090 ,n4089);
    not g3904(n4088 ,n4087);
    not g3905(n4086 ,n4085);
    not g3906(n4084 ,n4083);
    not g3907(n4082 ,n4081);
    not g3908(n4080 ,n4079);
    nor g3909(n4078 ,n3938 ,n4075);
    nor g3910(n4077 ,n4054 ,n4052);
    nor g3911(n4091 ,n4030 ,n4065);
    xnor g3912(n4089 ,n4008 ,n3978);
    xnor g3913(n4087 ,n4005 ,n3949);
    xnor g3914(n4085 ,n4007 ,n3952);
    xnor g3915(n4083 ,n4004 ,n3948);
    xnor g3916(n4081 ,n4003 ,n3906);
    xnor g3917(n4079 ,n4006 ,n3924);
    not g3918(n4072 ,n4071);
    not g3919(n4070 ,n4069);
    not g3920(n4068 ,n4067);
    nor g3921(n4066 ,n3977 ,n4033);
    nor g3922(n4065 ,n3930 ,n4029);
    nor g3923(n4064 ,n4038 ,n4035);
    nor g3924(n4063 ,n3940 ,n4016);
    nor g3925(n4062 ,n3964 ,n4020);
    nor g3926(n4061 ,n3965 ,n4021);
    nor g3927(n4060 ,n3941 ,n4017);
    nor g3928(n4059 ,n3976 ,n4031);
    nor g3929(n4076 ,n3980 ,n4013);
    nor g3930(n4075 ,n3993 ,n4024);
    nor g3931(n4074 ,n3995 ,n4011);
    nor g3932(n4073 ,n3984 ,n4037);
    nor g3933(n4071 ,n3992 ,n4025);
    nor g3934(n4069 ,n3994 ,n4027);
    nor g3935(n4067 ,n3989 ,n4015);
    not g3936(n4057 ,n4056);
    not g3937(n4055 ,n4054);
    not g3938(n4053 ,n4052);
    not g3939(n4051 ,n4050);
    not g3940(n4049 ,n4048);
    not g3941(n4047 ,n4046);
    xor g3942(n4590 ,n3953 ,n3900);
    xnor g3943(n4045 ,n3966 ,n3930);
    xnor g3944(n4044 ,n3926 ,n3974);
    xnor g3945(n4043 ,n3920 ,n3970);
    xnor g3946(n4042 ,n3968 ,n3942);
    xnor g3947(n4041 ,n3979 ,n3940);
    xnor g3948(n4040 ,n3972 ,n4001);
    xnor g3949(n4039 ,n3962 ,n3814);
    nor g3950(n4058 ,n3961 ,n4010);
    xnor g3951(n4056 ,n3955 ,n3908);
    nor g3952(n4054 ,n3986 ,n4009);
    xnor g3953(n4052 ,n3958 ,n3912);
    xnor g3954(n4050 ,n3957 ,n3946);
    xnor g3955(n4048 ,n3954 ,n3816);
    nor g3956(n4046 ,n3987 ,n4026);
    nor g3957(n4037 ,n3948 ,n3997);
    nor g3958(n4036 ,n4002 ,n3973);
    nor g3959(n4035 ,n3815 ,n3962);
    nor g3960(n4034 ,n3920 ,n3971);
    nor g3961(n4033 ,n3921 ,n3970);
    nor g3962(n4032 ,n3927 ,n3974);
    nor g3963(n4031 ,n3926 ,n3975);
    nor g3964(n4030 ,n3922 ,n3967);
    nor g3965(n4029 ,n3923 ,n3966);
    nor g3966(n4028 ,n3814 ,n3963);
    nor g3967(n4027 ,n3851 ,n3983);
    nor g3968(n4026 ,n3949 ,n3990);
    nor g3969(n4025 ,n3991 ,n3978);
    nor g3970(n4024 ,n3952 ,n3959);
    nor g3971(n4023 ,n3943 ,n3969);
    nor g3972(n4038 ,n3939 ,n3981);
    not g3973(n4021 ,n4020);
    not g3974(n4019 ,n4018);
    not g3975(n4017 ,n4016);
    nor g3976(n4015 ,n3950 ,n3988);
    nor g3977(n4014 ,n3942 ,n3968);
    nor g3978(n4013 ,n3899 ,n3996);
    nor g3979(n4012 ,n4001 ,n3972);
    nor g3980(n4011 ,n3784 ,n3960);
    nor g3981(n4010 ,n3931 ,n3982);
    nor g3982(n4009 ,n3876 ,n3985);
    xnor g3983(n4008 ,n3904 ,n3849);
    xnor g3984(n4007 ,n3706 ,n3918);
    xnor g3985(n4006 ,n3928 ,n3950);
    xnor g3986(n4005 ,n3916 ,n3914);
    xnor g3987(n4004 ,n3944 ,n3895);
    xnor g3988(n4003 ,n3931 ,n3871);
    nor g3989(n4022 ,n3891 ,n3998);
    xnor g3990(n4020 ,n3902 ,n3951);
    xnor g3991(n4018 ,n3901 ,n3822);
    xnor g3992(n4016 ,n3903 ,n3910);
    not g3993(n4002 ,n4001);
    not g3994(n4000 ,n3999);
    nor g3995(n3998 ,n3890 ,n3951);
    nor g3996(n3997 ,n3896 ,n3945);
    nor g3997(n3996 ,n3811 ,n3947);
    nor g3998(n3995 ,n3870 ,n3913);
    nor g3999(n3994 ,n3715 ,n3911);
    nor g4000(n3993 ,n3707 ,n3919);
    nor g4001(n3992 ,n3849 ,n3905);
    nor g4002(n3991 ,n3850 ,n3904);
    nor g4003(n3990 ,n3915 ,n3916);
    nor g4004(n3989 ,n3928 ,n3925);
    nor g4005(n3988 ,n3929 ,n3924);
    nor g4006(n3987 ,n3914 ,n3917);
    nor g4007(n3986 ,n3867 ,n3909);
    nor g4008(n3985 ,n3868 ,n3908);
    nor g4009(n3984 ,n3895 ,n3944);
    nor g4010(n3983 ,n3714 ,n3910);
    nor g4011(n3982 ,n3872 ,n3907);
    nor g4012(n3981 ,n3900 ,n3932);
    nor g4013(n3980 ,n3810 ,n3946);
    nor g4014(n4001 ,n3837 ,n3936);
    nor g4015(n3999 ,n3846 ,n3937);
    not g4016(n3975 ,n3974);
    not g4017(n3973 ,n3972);
    not g4018(n3971 ,n3970);
    not g4019(n3969 ,n3968);
    not g4020(n3967 ,n3966);
    not g4021(n3965 ,n3964);
    not g4022(n3963 ,n3962);
    nor g4023(n3961 ,n3871 ,n3906);
    nor g4024(n3960 ,n3869 ,n3912);
    nor g4025(n3959 ,n3706 ,n3918);
    xnor g4026(n4589 ,n3533 ,n3853);
    xor g4027(n3958 ,n3870 ,n3784);
    xnor g4028(n3957 ,n3899 ,n3810);
    xnor g4029(n3956 ,n3820 ,n3897);
    xnor g4030(n3955 ,n3867 ,n3876);
    xnor g4031(n3954 ,n3724 ,n3873);
    xnor g4032(n3953 ,n3704 ,n3865);
    nor g4033(n3979 ,n3888 ,n3933);
    xnor g4034(n3978 ,n3860 ,n3787);
    xnor g4035(n3977 ,n3855 ,n3874);
    nor g4036(n3976 ,n3887 ,n3935);
    xnor g4037(n3974 ,n3856 ,n3783);
    xnor g4038(n3972 ,n3854 ,n3718);
    xnor g4039(n3970 ,n3852 ,n3775);
    xnor g4040(n3968 ,n3859 ,n3785);
    xnor g4041(n3966 ,n3861 ,n3740);
    xnor g4042(n3964 ,n3858 ,n3746);
    xnor g4043(n3962 ,n3857 ,n3877);
    not g4044(n3947 ,n3946);
    not g4045(n3945 ,n3944);
    not g4046(n3943 ,n3942);
    not g4047(n3941 ,n3940);
    nor g4048(n3939 ,n3705 ,n3866);
    nor g4049(n3938 ,n3898 ,n3821);
    nor g4050(n3937 ,n3848 ,n3878);
    nor g4051(n3936 ,n3830 ,n3875);
    nor g4052(n3935 ,n3873 ,n3885);
    nor g4053(n3934 ,n3897 ,n3820);
    nor g4054(n3933 ,n3822 ,n3886);
    nor g4055(n3932 ,n3704 ,n3865);
    nor g4056(n3952 ,n3825 ,n3882);
    nor g4057(n3951 ,n3844 ,n3889);
    nor g4058(n3950 ,n3834 ,n3880);
    nor g4059(n3949 ,n3847 ,n3881);
    nor g4060(n3948 ,n3845 ,n3893);
    nor g4061(n3946 ,n3835 ,n3892);
    nor g4062(n3944 ,n3840 ,n3883);
    nor g4063(n3942 ,n3824 ,n3884);
    nor g4064(n3940 ,n3836 ,n3879);
    not g4065(n3929 ,n3928);
    not g4066(n3927 ,n3926);
    not g4067(n3925 ,n3924);
    not g4068(n3923 ,n3922);
    not g4069(n3921 ,n3920);
    not g4070(n3919 ,n3918);
    not g4071(n3917 ,n3916);
    not g4072(n3915 ,n3914);
    not g4073(n3913 ,n3912);
    not g4074(n3911 ,n3910);
    not g4075(n3909 ,n3908);
    not g4076(n3907 ,n3906);
    not g4077(n3905 ,n3904);
    xnor g4078(n3903 ,n3714 ,n3851);
    xnor g4079(n3902 ,n3742 ,n3812);
    xnor g4080(n3901 ,n3732 ,n3818);
    nor g4081(n3931 ,n3842 ,n3894);
    nor g4082(n3930 ,n3828 ,n3863);
    xnor g4083(n3928 ,n3792 ,n3669);
    xnor g4084(n3926 ,n3789 ,n3708);
    xnor g4085(n3924 ,n3791 ,n3781);
    nor g4086(n3922 ,n3843 ,n3864);
    xnor g4087(n3920 ,n3799 ,n3692);
    xnor g4088(n3918 ,n3794 ,n3696);
    xnor g4089(n3916 ,n3795 ,n3734);
    nor g4090(n3914 ,n3827 ,n3862);
    xnor g4091(n3912 ,n3790 ,n3728);
    xnor g4092(n3910 ,n3798 ,n3722);
    xnor g4093(n3908 ,n3788 ,n3712);
    xnor g4094(n3906 ,n3796 ,n3670);
    xnor g4095(n3904 ,n3793 ,n3645);
    not g4096(n3898 ,n3897);
    not g4097(n3896 ,n3895);
    nor g4098(n3894 ,n3786 ,n3807);
    nor g4099(n3893 ,n3747 ,n3802);
    nor g4100(n3892 ,n3749 ,n3832);
    nor g4101(n3891 ,n3743 ,n3812);
    nor g4102(n3890 ,n3742 ,n3813);
    nor g4103(n3889 ,n3748 ,n3801);
    nor g4104(n3888 ,n3733 ,n3818);
    nor g4105(n3887 ,n3725 ,n3816);
    nor g4106(n3886 ,n3732 ,n3819);
    nor g4107(n3885 ,n3724 ,n3817);
    nor g4108(n3884 ,n3787 ,n3805);
    nor g4109(n3883 ,n3693 ,n3839);
    nor g4110(n3882 ,n3663 ,n3829);
    nor g4111(n3881 ,n3783 ,n3808);
    nor g4112(n3880 ,n3664 ,n3833);
    nor g4113(n3879 ,n3671 ,n3831);
    nor g4114(n3900 ,n3634 ,n3838);
    nor g4115(n3899 ,n3766 ,n3800);
    nor g4116(n3897 ,n3762 ,n3804);
    nor g4117(n3895 ,n3760 ,n3823);
    not g4118(n3878 ,n3877);
    not g4119(n3875 ,n3874);
    not g4120(n3872 ,n3871);
    not g4121(n3870 ,n3869);
    not g4122(n3868 ,n3867);
    not g4123(n3866 ,n3865);
    nor g4124(n3864 ,n3785 ,n3803);
    nor g4125(n3863 ,n3691 ,n3826);
    nor g4126(n3862 ,n3690 ,n3841);
    xor g4127(n3861 ,n3748 ,n3738);
    xnor g4128(n3860 ,n3779 ,n3767);
    xnor g4129(n3859 ,n3726 ,n3716);
    xnor g4130(n3858 ,n3720 ,n3736);
    xnor g4131(n3857 ,n3771 ,n3769);
    xnor g4132(n3856 ,n3777 ,n3773);
    xnor g4133(n3855 ,n3730 ,n3685);
    xor g4134(n3854 ,n3749 ,n3687);
    xnor g4135(n3853 ,n3744 ,n3401);
    xor g4136(n3852 ,n3710 ,n3786);
    xnor g4137(n3877 ,n3698 ,n3694);
    nor g4138(n3876 ,n3761 ,n3809);
    xnor g4139(n3874 ,n3701 ,n3667);
    xnor g4140(n3873 ,n3700 ,n3534);
    nor g4141(n3871 ,n3750 ,n3806);
    xnor g4142(n3869 ,n3699 ,n3666);
    xnor g4143(n3867 ,n3702 ,n3538);
    xnor g4144(n3865 ,n3703 ,n3689);
    not g4145(n3850 ,n3849);
    nor g4146(n3848 ,n3771 ,n3769);
    nor g4147(n3847 ,n3778 ,n3774);
    nor g4148(n3846 ,n3772 ,n3770);
    nor g4149(n3845 ,n3721 ,n3737);
    nor g4150(n3844 ,n3741 ,n3739);
    nor g4151(n3843 ,n3727 ,n3717);
    nor g4152(n3842 ,n3776 ,n3711);
    nor g4153(n3841 ,n3650 ,n3708);
    nor g4154(n3840 ,n3657 ,n3782);
    nor g4155(n3839 ,n3658 ,n3781);
    nor g4156(n3838 ,n3598 ,n3745);
    nor g4157(n3837 ,n3685 ,n3731);
    nor g4158(n3836 ,n3659 ,n3735);
    nor g4159(n3835 ,n3687 ,n3719);
    nor g4160(n3834 ,n3653 ,n3729);
    nor g4161(n3833 ,n3654 ,n3728);
    nor g4162(n3832 ,n3688 ,n3718);
    nor g4163(n3831 ,n3660 ,n3734);
    nor g4164(n3830 ,n3686 ,n3730);
    nor g4165(n3829 ,n3656 ,n3722);
    nor g4166(n3828 ,n3683 ,n3713);
    nor g4167(n3827 ,n3649 ,n3709);
    nor g4168(n3826 ,n3684 ,n3712);
    nor g4169(n3825 ,n3655 ,n3723);
    nor g4170(n3824 ,n3780 ,n3768);
    nor g4171(n3823 ,n3669 ,n3758);
    nor g4172(n3851 ,n3530 ,n3752);
    nor g4173(n3849 ,n3673 ,n3759);
    not g4174(n3821 ,n3820);
    not g4175(n3819 ,n3818);
    not g4176(n3817 ,n3816);
    not g4177(n3815 ,n3814);
    not g4178(n3813 ,n3812);
    not g4179(n3811 ,n3810);
    nor g4180(n3809 ,n3695 ,n3763);
    nor g4181(n3808 ,n3777 ,n3773);
    nor g4182(n3807 ,n3775 ,n3710);
    nor g4183(n3806 ,n3692 ,n3765);
    nor g4184(n3805 ,n3779 ,n3767);
    nor g4185(n3804 ,n3696 ,n3764);
    nor g4186(n3803 ,n3726 ,n3716);
    nor g4187(n3802 ,n3720 ,n3736);
    nor g4188(n3801 ,n3740 ,n3738);
    nor g4189(n3800 ,n3670 ,n3755);
    xnor g4190(n3799 ,n3647 ,n3651);
    xnor g4191(n3798 ,n3655 ,n3663);
    nor g4192(n3797 ,n3502 ,n3753);
    xnor g4193(n3796 ,n3641 ,n3643);
    xnor g4194(n3795 ,n3671 ,n3659);
    xnor g4195(n3794 ,n3247 ,n3661);
    xnor g4196(n3793 ,n3497 ,n3695);
    xnor g4197(n3792 ,n3585 ,n3681);
    xnor g4198(n3791 ,n3657 ,n3693);
    xnor g4199(n3790 ,n3653 ,n3664);
    xnor g4200(n3789 ,n3649 ,n3690);
    xnor g4201(n3788 ,n3683 ,n3691);
    nor g4202(n3822 ,n3636 ,n3756);
    xnor g4203(n3820 ,n3561 ,n3665);
    xnor g4204(n3818 ,n3549 ,n3697);
    nor g4205(n3816 ,n3675 ,n3751);
    nor g4206(n3814 ,n3672 ,n3757);
    nor g4207(n3812 ,n3678 ,n3754);
    xnor g4208(n3810 ,n3638 ,n3668);
    not g4209(n3782 ,n3781);
    not g4210(n3780 ,n3779);
    not g4211(n3778 ,n3777);
    not g4212(n3776 ,n3775);
    not g4213(n3774 ,n3773);
    not g4214(n3772 ,n3771);
    not g4215(n3770 ,n3769);
    not g4216(n3768 ,n3767);
    nor g4217(n3766 ,n3643 ,n3641);
    nor g4218(n3765 ,n3652 ,n3648);
    nor g4219(n3764 ,n3247 ,n3662);
    nor g4220(n3763 ,n3497 ,n3646);
    nor g4221(n3762 ,n3248 ,n3661);
    nor g4222(n3761 ,n3498 ,n3645);
    nor g4223(n3760 ,n3585 ,n3681);
    nor g4224(n3759 ,n3694 ,n3676);
    nor g4225(n3758 ,n3586 ,n3682);
    nor g4226(n3757 ,n3689 ,n3679);
    nor g4227(n3756 ,n3600 ,n3668);
    nor g4228(n3755 ,n3644 ,n3642);
    nor g4229(n3754 ,n3666 ,n3677);
    nor g4230(n3753 ,n3496 ,n3665);
    nor g4231(n3752 ,n3493 ,n3697);
    nor g4232(n3751 ,n3667 ,n3674);
    nor g4233(n3750 ,n3651 ,n3647);
    xnor g4234(n3787 ,n3551 ,n3595);
    xor g4235(n3786 ,n3580 ,n3431);
    nor g4236(n3785 ,n3509 ,n3640);
    nor g4237(n3784 ,n3635 ,n3639);
    nor g4238(n3783 ,n3616 ,n3680);
    xnor g4239(n3781 ,n3577 ,n3239);
    xnor g4240(n3779 ,n3596 ,n3217);
    xnor g4241(n3777 ,n3556 ,n3453);
    xnor g4242(n3775 ,n3555 ,n3299);
    xnor g4243(n3773 ,n3578 ,n3387);
    xnor g4244(n3771 ,n3582 ,n3265);
    xnor g4245(n3769 ,n3554 ,n3415);
    xnor g4246(n3767 ,n3581 ,n3413);
    not g4247(n3747 ,n3746);
    not g4248(n3745 ,n3744);
    not g4249(n3743 ,n3742);
    not g4250(n3741 ,n3740);
    not g4251(n3739 ,n3738);
    not g4252(n3737 ,n3736);
    not g4253(n3735 ,n3734);
    not g4254(n3733 ,n3732);
    not g4255(n3731 ,n3730);
    not g4256(n3729 ,n3728);
    not g4257(n3727 ,n3726);
    not g4258(n3725 ,n3724);
    not g4259(n3723 ,n3722);
    not g4260(n3721 ,n3720);
    not g4261(n3719 ,n3718);
    not g4262(n3717 ,n3716);
    not g4263(n3715 ,n3714);
    not g4264(n3713 ,n3712);
    not g4265(n3711 ,n3710);
    not g4266(n3709 ,n3708);
    not g4267(n3707 ,n3706);
    not g4268(n3705 ,n3704);
    xnor g4269(n3703 ,n3587 ,n3269);
    xnor g4270(n3702 ,n3594 ,n3347);
    xnor g4271(n3701 ,n3589 ,n3542);
    xnor g4272(n3700 ,n3593 ,n3253);
    xnor g4273(n3699 ,n3583 ,n3540);
    xnor g4274(n3698 ,n3591 ,n3544);
    xor g4275(n3749 ,n3557 ,n3451);
    xor g4276(n3748 ,n3558 ,n3311);
    xnor g4277(n3746 ,n3571 ,n3237);
    xnor g4278(n3744 ,n3570 ,n3219);
    xnor g4279(n3742 ,n3564 ,n3546);
    xnor g4280(n3740 ,n3548 ,n3449);
    xnor g4281(n3738 ,n3560 ,n3317);
    xnor g4282(n3736 ,n3567 ,n3307);
    xnor g4283(n3734 ,n3566 ,n3428);
    xnor g4284(n3732 ,n3552 ,n3209);
    xnor g4285(n3730 ,n3550 ,n3417);
    xnor g4286(n3728 ,n3573 ,n3434);
    xnor g4287(n3726 ,n3575 ,n3326);
    xnor g4288(n3724 ,n3559 ,n3309);
    xnor g4289(n3722 ,n3563 ,n3322);
    xnor g4290(n3720 ,n3569 ,n3291);
    xnor g4291(n3718 ,n3565 ,n3409);
    xnor g4292(n3716 ,n3562 ,n3438);
    xnor g4293(n3714 ,n3574 ,n3420);
    xnor g4294(n3712 ,n3553 ,n3320);
    xnor g4295(n3710 ,n3576 ,n3313);
    xnor g4296(n3708 ,n3579 ,n3407);
    xnor g4297(n3706 ,n3568 ,n3436);
    xnor g4298(n3704 ,n3572 ,n3341);
    not g4299(n3688 ,n3687);
    not g4300(n3686 ,n3685);
    not g4301(n3684 ,n3683);
    not g4302(n3682 ,n3681);
    nor g4303(n3680 ,n3599 ,n3593);
    nor g4304(n3679 ,n3269 ,n3588);
    nor g4305(n3678 ,n3541 ,n3583);
    nor g4306(n3677 ,n3540 ,n3584);
    nor g4307(n3676 ,n3544 ,n3592);
    nor g4308(n3675 ,n3543 ,n3589);
    nor g4309(n3674 ,n3542 ,n3590);
    nor g4310(n3673 ,n3545 ,n3591);
    nor g4311(n3672 ,n3270 ,n3587);
    nor g4312(n3697 ,n3517 ,n3629);
    nor g4313(n3696 ,n3515 ,n3614);
    nor g4314(n3695 ,n3527 ,n3601);
    nor g4315(n3694 ,n3518 ,n3630);
    nor g4316(n3693 ,n3526 ,n3631);
    nor g4317(n3692 ,n3523 ,n3603);
    nor g4318(n3691 ,n3528 ,n3605);
    nor g4319(n3690 ,n3508 ,n3610);
    nor g4320(n3689 ,n3525 ,n3627);
    nor g4321(n3687 ,n3516 ,n3619);
    nor g4322(n3685 ,n3531 ,n3622);
    nor g4323(n3683 ,n3520 ,n3606);
    nor g4324(n3681 ,n3499 ,n3611);
    not g4325(n3662 ,n3661);
    not g4326(n3660 ,n3659);
    not g4327(n3658 ,n3657);
    not g4328(n3656 ,n3655);
    not g4329(n3654 ,n3653);
    not g4330(n3652 ,n3651);
    not g4331(n3650 ,n3649);
    not g4332(n3648 ,n3647);
    not g4333(n3646 ,n3645);
    not g4334(n3644 ,n3643);
    not g4335(n3642 ,n3641);
    nor g4336(n3640 ,n3489 ,n3595);
    nor g4337(n3639 ,n3597 ,n3594);
    xnor g4338(n3638 ,n3536 ,n3357);
    nor g4339(n3671 ,n3514 ,n3617);
    nor g4340(n3670 ,n3510 ,n3613);
    nor g4341(n3669 ,n3476 ,n3628);
    nor g4342(n3668 ,n3512 ,n3608);
    nor g4343(n3667 ,n3500 ,n3607);
    nor g4344(n3666 ,n3503 ,n3637);
    nor g4345(n3665 ,n3519 ,n3621);
    nor g4346(n3664 ,n3501 ,n3618);
    nor g4347(n3663 ,n3495 ,n3612);
    nor g4348(n3661 ,n3505 ,n3609);
    nor g4349(n3659 ,n3521 ,n3624);
    nor g4350(n3657 ,n3513 ,n3626);
    nor g4351(n3655 ,n3494 ,n3623);
    nor g4352(n3653 ,n3504 ,n3620);
    nor g4353(n3651 ,n3529 ,n3625);
    nor g4354(n3649 ,n3522 ,n3604);
    nor g4355(n3647 ,n3507 ,n3632);
    nor g4356(n3645 ,n3524 ,n3602);
    nor g4357(n3643 ,n3511 ,n3615);
    nor g4358(n3641 ,n3506 ,n3633);
    nor g4359(n3637 ,n3439 ,n3472);
    nor g4360(n3636 ,n3358 ,n3537);
    nor g4361(n3635 ,n3348 ,n3539);
    nor g4362(n3634 ,n3402 ,n3532);
    nor g4363(n3633 ,n3418 ,n3487);
    nor g4364(n3632 ,n3308 ,n3466);
    nor g4365(n3631 ,n3312 ,n3464);
    nor g4366(n3630 ,n3330 ,n3488);
    nor g4367(n3629 ,n3454 ,n3468);
    nor g4368(n3628 ,n3450 ,n3457);
    nor g4369(n3627 ,n3319 ,n3484);
    nor g4370(n3626 ,n3318 ,n3481);
    nor g4371(n3625 ,n3448 ,n3471);
    nor g4372(n3624 ,n3433 ,n3459);
    nor g4373(n3623 ,n3430 ,n3480);
    nor g4374(n3622 ,n3485 ,n3547);
    nor g4375(n3621 ,n3437 ,n3467);
    nor g4376(n3620 ,n3327 ,n3490);
    nor g4377(n3619 ,n3300 ,n3475);
    nor g4378(n3618 ,n3321 ,n3479);
    nor g4379(n3617 ,n3301 ,n3473);
    nor g4380(n3616 ,n3254 ,n3535);
    nor g4381(n3615 ,n3432 ,n3491);
    nor g4382(n3614 ,n3323 ,n3470);
    nor g4383(n3613 ,n3314 ,n3462);
    nor g4384(n3612 ,n3429 ,n3486);
    nor g4385(n3611 ,n3435 ,n3469);
    nor g4386(n3610 ,n3452 ,n3474);
    nor g4387(n3609 ,n3421 ,n3482);
    nor g4388(n3608 ,n3410 ,n3478);
    nor g4389(n3607 ,n3292 ,n3465);
    nor g4390(n3606 ,n3414 ,n3461);
    nor g4391(n3605 ,n3412 ,n3492);
    nor g4392(n3604 ,n3310 ,n3477);
    nor g4393(n3603 ,n3419 ,n3483);
    nor g4394(n3602 ,n3416 ,n3458);
    nor g4395(n3601 ,n3304 ,n3460);
    nor g4396(n3600 ,n3357 ,n3536);
    nor g4397(n3599 ,n3253 ,n3534);
    nor g4398(n3598 ,n3401 ,n3533);
    nor g4399(n3597 ,n3347 ,n3538);
    nor g4400(n4588 ,n3463 ,n3533);
    xnor g4401(n3596 ,n3411 ,n3257);
    not g4402(n3592 ,n3591);
    not g4403(n3590 ,n3589);
    not g4404(n3588 ,n3587);
    not g4405(n3586 ,n3585);
    not g4406(n3584 ,n3583);
    xor g4407(n3582 ,n3304 ,n3213);
    xnor g4408(n3581 ,n3227 ,n3381);
    xnor g4409(n3580 ,n3337 ,n3215);
    xor g4410(n3579 ,n3433 ,n3225);
    xor g4411(n3578 ,n3301 ,n3385);
    xor g4412(n3577 ,n3448 ,n3373);
    xnor g4413(n3576 ,n3229 ,n3345);
    xnor g4414(n3575 ,n3349 ,n3369);
    xnor g4415(n3574 ,n3255 ,n3353);
    xnor g4416(n3573 ,n3245 ,n3221);
    xor g4417(n3572 ,n3330 ,n3393);
    xor g4418(n3571 ,n3419 ,n3267);
    xor g4419(n3570 ,n3319 ,n3389);
    xnor g4420(n3569 ,n3281 ,n3339);
    xnor g4421(n3568 ,n3391 ,n3259);
    xnor g4422(n3567 ,n3375 ,n3333);
    xnor g4423(n3566 ,n3241 ,n3233);
    xnor g4424(n3565 ,n3371 ,n3395);
    xnor g4425(n3564 ,n3235 ,n3275);
    xnor g4426(n3563 ,n3249 ,n3383);
    xnor g4427(n3562 ,n3285 ,n3283);
    xnor g4428(n3561 ,n3377 ,n3359);
    xnor g4429(n3560 ,n3365 ,n3231);
    xnor g4430(n3559 ,n3403 ,n3397);
    xnor g4431(n3558 ,n3343 ,n3211);
    xnor g4432(n3557 ,n3399 ,n3335);
    xnor g4433(n3556 ,n3351 ,n3263);
    xnor g4434(n3555 ,n3405 ,n3363);
    xnor g4435(n3554 ,n3367 ,n3277);
    xnor g4436(n3553 ,n3379 ,n3223);
    xor g4437(n3552 ,n3430 ,n3361);
    xnor g4438(n3551 ,n3261 ,n3251);
    xnor g4439(n3550 ,n3273 ,n3287);
    xnor g4440(n3549 ,n3279 ,n3271);
    xnor g4441(n3548 ,n3355 ,n3243);
    xnor g4442(n3595 ,n3442 ,n3315);
    xnor g4443(n3594 ,n3424 ,n3297);
    xnor g4444(n3593 ,n3328 ,n3422);
    xnor g4445(n3591 ,n3426 ,n3289);
    xnor g4446(n3589 ,n3295 ,n3444);
    xnor g4447(n3587 ,n3324 ,n3293);
    xnor g4448(n3585 ,n3446 ,n3440);
    xnor g4449(n3583 ,n3302 ,n3305);
    not g4450(n3547 ,n3546);
    not g4451(n3545 ,n3544);
    not g4452(n3543 ,n3542);
    not g4453(n3541 ,n3540);
    not g4454(n3539 ,n3538);
    not g4455(n3537 ,n3536);
    not g4456(n3535 ,n3534);
    not g4457(n3532 ,n3533);
    nor g4458(n3531 ,n3276 ,n3236);
    nor g4459(n3530 ,n3272 ,n3280);
    nor g4460(n3529 ,n3240 ,n3374);
    nor g4461(n3528 ,n3258 ,n3218);
    nor g4462(n3527 ,n3214 ,n3266);
    nor g4463(n3526 ,n3212 ,n3344);
    nor g4464(n3525 ,n3390 ,n3220);
    nor g4465(n3524 ,n3278 ,n3368);
    nor g4466(n3523 ,n3238 ,n3268);
    nor g4467(n3522 ,n3398 ,n3404);
    nor g4468(n3521 ,n3408 ,n3226);
    nor g4469(n3520 ,n3382 ,n3228);
    nor g4470(n3519 ,n3260 ,n3392);
    nor g4471(n3518 ,n3342 ,n3394);
    nor g4472(n3517 ,n3264 ,n3352);
    nor g4473(n3516 ,n3364 ,n3406);
    nor g4474(n3515 ,n3384 ,n3250);
    nor g4475(n3514 ,n3386 ,n3388);
    nor g4476(n3513 ,n3232 ,n3366);
    nor g4477(n3512 ,n3396 ,n3372);
    nor g4478(n3511 ,n3216 ,n3338);
    nor g4479(n3510 ,n3346 ,n3230);
    nor g4480(n3509 ,n3252 ,n3262);
    nor g4481(n3508 ,n3336 ,n3400);
    nor g4482(n3507 ,n3334 ,n3376);
    nor g4483(n3506 ,n3288 ,n3274);
    nor g4484(n3505 ,n3354 ,n3256);
    nor g4485(n3504 ,n3370 ,n3350);
    nor g4486(n3503 ,n3284 ,n3286);
    nor g4487(n3502 ,n3360 ,n3378);
    nor g4488(n3501 ,n3224 ,n3380);
    nor g4489(n3500 ,n3340 ,n3282);
    nor g4490(n3499 ,n3222 ,n3246);
    nor g4491(n3546 ,n3306 ,n3303);
    nor g4492(n3544 ,n3294 ,n3325);
    nor g4493(n3542 ,n3441 ,n3447);
    nor g4494(n3540 ,n3298 ,n3425);
    nor g4495(n3538 ,n3316 ,n3443);
    nor g4496(n3536 ,n3423 ,n3329);
    nor g4497(n3534 ,n3445 ,n3296);
    nor g4498(n3533 ,n3332 ,n3456);
    not g4499(n3498 ,n3497);
    nor g4500(n3496 ,n3359 ,n3377);
    nor g4501(n3495 ,n3234 ,n3242);
    nor g4502(n3494 ,n3210 ,n3362);
    nor g4503(n3493 ,n3271 ,n3279);
    nor g4504(n3492 ,n3257 ,n3217);
    nor g4505(n3491 ,n3215 ,n3337);
    nor g4506(n3490 ,n3369 ,n3349);
    nor g4507(n3489 ,n3251 ,n3261);
    nor g4508(n3488 ,n3341 ,n3393);
    nor g4509(n3487 ,n3287 ,n3273);
    nor g4510(n3486 ,n3233 ,n3241);
    nor g4511(n3485 ,n3275 ,n3235);
    nor g4512(n3484 ,n3389 ,n3219);
    nor g4513(n3483 ,n3237 ,n3267);
    nor g4514(n3482 ,n3353 ,n3255);
    nor g4515(n3481 ,n3231 ,n3365);
    nor g4516(n3480 ,n3209 ,n3361);
    nor g4517(n3479 ,n3223 ,n3379);
    nor g4518(n3478 ,n3395 ,n3371);
    nor g4519(n3477 ,n3397 ,n3403);
    nor g4520(n3476 ,n3244 ,n3356);
    nor g4521(n3475 ,n3363 ,n3405);
    nor g4522(n3474 ,n3335 ,n3399);
    nor g4523(n3473 ,n3385 ,n3387);
    nor g4524(n3472 ,n3283 ,n3285);
    nor g4525(n3471 ,n3239 ,n3373);
    nor g4526(n3470 ,n3383 ,n3249);
    nor g4527(n3469 ,n3221 ,n3245);
    nor g4528(n3468 ,n3263 ,n3351);
    nor g4529(n3467 ,n3259 ,n3391);
    nor g4530(n3466 ,n3333 ,n3375);
    nor g4531(n3465 ,n3339 ,n3281);
    nor g4532(n3464 ,n3211 ,n3343);
    nor g4533(n3463 ,n3331 ,n3455);
    nor g4534(n3462 ,n3345 ,n3229);
    nor g4535(n3461 ,n3381 ,n3227);
    nor g4536(n3460 ,n3213 ,n3265);
    nor g4537(n3459 ,n3407 ,n3225);
    nor g4538(n3458 ,n3277 ,n3367);
    nor g4539(n3457 ,n3243 ,n3355);
    nor g4540(n3497 ,n3290 ,n3427);
    not g4541(n3456 ,n3455);
    not g4542(n3454 ,n3453);
    not g4543(n3452 ,n3451);
    not g4544(n3450 ,n3449);
    not g4545(n3447 ,n3446);
    not g4546(n3445 ,n3444);
    not g4547(n3443 ,n3442);
    not g4548(n3441 ,n3440);
    not g4549(n3439 ,n3438);
    not g4550(n3437 ,n3436);
    not g4551(n3435 ,n3434);
    not g4552(n3432 ,n3431);
    not g4553(n3429 ,n3428);
    not g4554(n3427 ,n3426);
    not g4555(n3425 ,n3424);
    not g4556(n3423 ,n3422);
    not g4557(n3421 ,n3420);
    not g4558(n3418 ,n3417);
    not g4559(n3416 ,n3415);
    not g4560(n3414 ,n3413);
    not g4561(n3412 ,n3411);
    not g4562(n3410 ,n3409);
    not g4563(n3408 ,n3407);
    not g4564(n3406 ,n3405);
    not g4565(n3404 ,n3403);
    not g4566(n3402 ,n3401);
    not g4567(n3400 ,n3399);
    not g4568(n3398 ,n3397);
    not g4569(n3396 ,n3395);
    not g4570(n3394 ,n3393);
    not g4571(n3392 ,n3391);
    not g4572(n3390 ,n3389);
    not g4573(n3388 ,n3387);
    not g4574(n3386 ,n3385);
    not g4575(n3384 ,n3383);
    not g4576(n3382 ,n3381);
    not g4577(n3380 ,n3379);
    not g4578(n3378 ,n3377);
    not g4579(n3376 ,n3375);
    not g4580(n3374 ,n3373);
    not g4581(n3372 ,n3371);
    not g4582(n3370 ,n3369);
    not g4583(n3368 ,n3367);
    not g4584(n3366 ,n3365);
    not g4585(n3364 ,n3363);
    not g4586(n3362 ,n3361);
    not g4587(n3360 ,n3359);
    not g4588(n3358 ,n3357);
    not g4589(n3356 ,n3355);
    not g4590(n3354 ,n3353);
    not g4591(n3352 ,n3351);
    not g4592(n3350 ,n3349);
    not g4593(n3348 ,n3347);
    not g4594(n3346 ,n3345);
    not g4595(n3344 ,n3343);
    not g4596(n3342 ,n3341);
    not g4597(n3340 ,n3339);
    not g4598(n3338 ,n3337);
    not g4599(n3336 ,n3335);
    not g4600(n3334 ,n3333);
    nor g4601(n3455 ,n3198 ,n3182);
    nor g4602(n3453 ,n3187 ,n3188);
    nor g4603(n3451 ,n3201 ,n3178);
    nor g4604(n3449 ,n3201 ,n3207);
    or g4605(n3448 ,n3195 ,n3204);
    nor g4606(n3446 ,n3183 ,n3191);
    nor g4607(n3444 ,n3196 ,n3190);
    nor g4608(n3442 ,n3187 ,n3191);
    nor g4609(n3440 ,n3196 ,n3192);
    nor g4610(n3438 ,n3200 ,n3204);
    nor g4611(n3436 ,n3179 ,n3178);
    nor g4612(n3434 ,n3195 ,n3194);
    or g4613(n3433 ,n3206 ,n3184);
    nor g4614(n3431 ,n3200 ,n3205);
    or g4615(n3430 ,n3206 ,n3178);
    nor g4616(n3428 ,n3187 ,n3177);
    nor g4617(n3426 ,n3202 ,n3191);
    nor g4618(n3424 ,n3180 ,n3191);
    nor g4619(n3422 ,n3196 ,n3193);
    nor g4620(n3420 ,n3208 ,n3205);
    or g4621(n3419 ,n3200 ,n3207);
    nor g4622(n3417 ,n3185 ,n3178);
    nor g4623(n3415 ,n3185 ,n3204);
    nor g4624(n3413 ,n3185 ,n3186);
    nor g4625(n3411 ,n3198 ,n3207);
    nor g4626(n3409 ,n3195 ,n3207);
    nor g4627(n3407 ,n3202 ,n3177);
    nor g4628(n3405 ,n3195 ,n3186);
    nor g4629(n3403 ,n3206 ,n3205);
    nor g4630(n3401 ,n3199 ,n3192);
    nor g4631(n3399 ,n3180 ,n3197);
    nor g4632(n3397 ,n3202 ,n3188);
    nor g4633(n3395 ,n3187 ,n3189);
    nor g4634(n3393 ,n3201 ,n3182);
    nor g4635(n3391 ,n3183 ,n3188);
    nor g4636(n3389 ,n3181 ,n3191);
    nor g4637(n3387 ,n3208 ,n3186);
    nor g4638(n3385 ,n3180 ,n3189);
    nor g4639(n3383 ,n3180 ,n3177);
    nor g4640(n3381 ,n3181 ,n3193);
    nor g4641(n3379 ,n3202 ,n3190);
    nor g4642(n3377 ,n3208 ,n3178);
    nor g4643(n3375 ,n3208 ,n3182);
    nor g4644(n3373 ,n3180 ,n3190);
    nor g4645(n3371 ,n3179 ,n3186);
    nor g4646(n3369 ,n3181 ,n3197);
    nor g4647(n3367 ,n3201 ,n3194);
    nor g4648(n3365 ,n3206 ,n3204);
    nor g4649(n3363 ,n3202 ,n3189);
    nor g4650(n3361 ,n3208 ,n3207);
    nor g4651(n3359 ,n3183 ,n3177);
    nor g4652(n3357 ,n3179 ,n3207);
    nor g4653(n3355 ,n3187 ,n3190);
    nor g4654(n3353 ,n3196 ,n3188);
    nor g4655(n3351 ,n3183 ,n3193);
    nor g4656(n3349 ,n3201 ,n3186);
    nor g4657(n3347 ,n3195 ,n3182);
    nor g4658(n3345 ,n3187 ,n3197);
    nor g4659(n3343 ,n3185 ,n3205);
    nor g4660(n3341 ,n3185 ,n3194);
    nor g4661(n3339 ,n3199 ,n3177);
    nor g4662(n3337 ,n3180 ,n3193);
    nor g4663(n3335 ,n3203 ,n3177);
    nor g4664(n3333 ,n3202 ,n3197);
    not g4665(n3332 ,n3331);
    not g4666(n3329 ,n3328);
    not g4667(n3327 ,n3326);
    not g4668(n3325 ,n3324);
    not g4669(n3323 ,n3322);
    not g4670(n3321 ,n3320);
    not g4671(n3318 ,n3317);
    not g4672(n3316 ,n3315);
    not g4673(n3314 ,n3313);
    not g4674(n3312 ,n3311);
    not g4675(n3310 ,n3309);
    not g4676(n3308 ,n3307);
    not g4677(n3306 ,n3305);
    not g4678(n3303 ,n3302);
    not g4679(n3300 ,n3299);
    not g4680(n3298 ,n3297);
    not g4681(n3296 ,n3295);
    not g4682(n3294 ,n3293);
    not g4683(n3292 ,n3291);
    not g4684(n3290 ,n3289);
    not g4685(n3288 ,n3287);
    not g4686(n3286 ,n3285);
    not g4687(n3284 ,n3283);
    not g4688(n3282 ,n3281);
    not g4689(n3280 ,n3279);
    not g4690(n3278 ,n3277);
    not g4691(n3276 ,n3275);
    not g4692(n3274 ,n3273);
    not g4693(n3272 ,n3271);
    not g4694(n3270 ,n3269);
    not g4695(n3268 ,n3267);
    not g4696(n3266 ,n3265);
    not g4697(n3264 ,n3263);
    not g4698(n3262 ,n3261);
    not g4699(n3260 ,n3259);
    not g4700(n3258 ,n3257);
    not g4701(n3256 ,n3255);
    not g4702(n3254 ,n3253);
    not g4703(n3252 ,n3251);
    not g4704(n3250 ,n3249);
    not g4705(n3248 ,n3247);
    not g4706(n3246 ,n3245);
    not g4707(n3244 ,n3243);
    not g4708(n3242 ,n3241);
    not g4709(n3240 ,n3239);
    not g4710(n3238 ,n3237);
    not g4711(n3236 ,n3235);
    not g4712(n3234 ,n3233);
    not g4713(n3232 ,n3231);
    not g4714(n3230 ,n3229);
    not g4715(n3228 ,n3227);
    not g4716(n3226 ,n3225);
    not g4717(n3224 ,n3223);
    not g4718(n3222 ,n3221);
    not g4719(n3220 ,n3219);
    not g4720(n3218 ,n3217);
    not g4721(n3216 ,n3215);
    not g4722(n3214 ,n3213);
    not g4723(n3212 ,n3211);
    not g4724(n3210 ,n3209);
    nor g4725(n3331 ,n3199 ,n3191);
    or g4726(n3330 ,n3198 ,n3204);
    nor g4727(n3328 ,n3183 ,n3190);
    nor g4728(n3326 ,n3185 ,n3207);
    nor g4729(n3324 ,n3203 ,n3191);
    nor g4730(n3322 ,n3195 ,n3178);
    nor g4731(n3320 ,n3198 ,n3205);
    or g4732(n3319 ,n3198 ,n3194);
    nor g4733(n3317 ,n3200 ,n3186);
    nor g4734(n3315 ,n3202 ,n3192);
    nor g4735(n3313 ,n3179 ,n3204);
    nor g4736(n3311 ,n3198 ,n3184);
    nor g4737(n3309 ,n3200 ,n3184);
    nor g4738(n3307 ,n3179 ,n3194);
    nor g4739(n3305 ,n3180 ,n3192);
    or g4740(n3304 ,n3198 ,n3186);
    nor g4741(n3302 ,n3196 ,n3191);
    or g4742(n3301 ,n3200 ,n3178);
    nor g4743(n3299 ,n3206 ,n3207);
    nor g4744(n3297 ,n3187 ,n3192);
    nor g4745(n3295 ,n3183 ,n3192);
    nor g4746(n3293 ,n3181 ,n3192);
    nor g4747(n3291 ,n3198 ,n3178);
    nor g4748(n3289 ,n3203 ,n3192);
    nor g4749(n3287 ,n3181 ,n3177);
    nor g4750(n3285 ,n3206 ,n3194);
    nor g4751(n3283 ,n3203 ,n3193);
    nor g4752(n3281 ,n3187 ,n3193);
    nor g4753(n3279 ,n3179 ,n3205);
    nor g4754(n3277 ,n3181 ,n3190);
    nor g4755(n3275 ,n3185 ,n3184);
    nor g4756(n3273 ,n3201 ,n3184);
    nor g4757(n3271 ,n3195 ,n3184);
    nor g4758(n3269 ,n3199 ,n3190);
    nor g4759(n3267 ,n3206 ,n3186);
    nor g4760(n3265 ,n3200 ,n3182);
    nor g4761(n3263 ,n3196 ,n3197);
    nor g4762(n3261 ,n3206 ,n3182);
    nor g4763(n3259 ,n3196 ,n3177);
    nor g4764(n3257 ,n3199 ,n3197);
    nor g4765(n3255 ,n3183 ,n3189);
    nor g4766(n3253 ,n3208 ,n3204);
    nor g4767(n3251 ,n3200 ,n3194);
    nor g4768(n3249 ,n3179 ,n3184);
    nor g4769(n3247 ,n3208 ,n3184);
    nor g4770(n3245 ,n3179 ,n3182);
    nor g4771(n3243 ,n3181 ,n3189);
    nor g4772(n3241 ,n3183 ,n3197);
    nor g4773(n3239 ,n3203 ,n3189);
    nor g4774(n3237 ,n3181 ,n3188);
    nor g4775(n3235 ,n3201 ,n3205);
    nor g4776(n3233 ,n3196 ,n3189);
    nor g4777(n3231 ,n3203 ,n3197);
    nor g4778(n3229 ,n3208 ,n3194);
    nor g4779(n3227 ,n3201 ,n3204);
    nor g4780(n3225 ,n3195 ,n3205);
    nor g4781(n3223 ,n3199 ,n3189);
    nor g4782(n3221 ,n3202 ,n3193);
    nor g4783(n3219 ,n3185 ,n3182);
    nor g4784(n3217 ,n3203 ,n3190);
    nor g4785(n3215 ,n3203 ,n3188);
    nor g4786(n3213 ,n3199 ,n3193);
    nor g4787(n3211 ,n3199 ,n3188);
    nor g4788(n3209 ,n3180 ,n3188);
    not g4789(n3208 ,n27[7]);
    not g4790(n3207 ,n4[4]);
    not g4791(n3206 ,n27[4]);
    not g4792(n3205 ,n4[5]);
    not g4793(n3204 ,n4[2]);
    not g4794(n3203 ,n28[2]);
    not g4795(n3202 ,n28[3]);
    not g4796(n3201 ,n27[2]);
    not g4797(n3200 ,n27[3]);
    not g4798(n3199 ,n28[0]);
    not g4799(n3198 ,n27[0]);
    not g4800(n3197 ,n26[4]);
    not g4801(n3196 ,n28[6]);
    not g4802(n3195 ,n27[5]);
    not g4803(n3194 ,n4[1]);
    not g4804(n3193 ,n26[3]);
    not g4805(n3192 ,n26[1]);
    not g4806(n3191 ,n26[0]);
    not g4807(n3190 ,n26[2]);
    not g4808(n3189 ,n26[5]);
    not g4809(n3188 ,n26[6]);
    not g4810(n3187 ,n28[4]);
    not g4811(n3186 ,n4[3]);
    not g4812(n3185 ,n27[1]);
    not g4813(n3184 ,n4[6]);
    not g4814(n3183 ,n28[7]);
    not g4815(n3182 ,n4[0]);
    not g4816(n3181 ,n28[1]);
    not g4817(n3180 ,n28[5]);
    not g4818(n3179 ,n27[6]);
    not g4819(n3178 ,n4[7]);
    not g4820(n3177 ,n26[7]);
    nor g4821(n4628 ,n4283 ,n4312);
    xnor g4822(n4627 ,n4291 ,n4311);
    nor g4823(n4312 ,n4291 ,n4311);
    nor g4824(n4311 ,n4284 ,n4310);
    xor g4825(n4626 ,n4292 ,n4308);
    nor g4826(n4310 ,n4292 ,n4309);
    not g4827(n4309 ,n4308);
    nor g4828(n4308 ,n4290 ,n4307);
    xor g4829(n4625 ,n4295 ,n4306);
    nor g4830(n4307 ,n4295 ,n4306);
    nor g4831(n4306 ,n4288 ,n4305);
    xor g4832(n4624 ,n4294 ,n4304);
    nor g4833(n4305 ,n4294 ,n4304);
    nor g4834(n4304 ,n4286 ,n4303);
    xor g4835(n4623 ,n4297 ,n4302);
    nor g4836(n4303 ,n4297 ,n4302);
    nor g4837(n4302 ,n4289 ,n4301);
    xnor g4838(n4622 ,n4296 ,n4299);
    nor g4839(n4301 ,n4296 ,n4300);
    not g4840(n4300 ,n4299);
    nor g4841(n4299 ,n4282 ,n4298);
    xnor g4842(n4621 ,n4293 ,n4287);
    nor g4843(n4298 ,n4287 ,n4293);
    xnor g4844(n4297 ,n4[3] ,n26[3]);
    nor g4845(n4620 ,n4287 ,n4285);
    xnor g4846(n4296 ,n4[2] ,n26[2]);
    xnor g4847(n4295 ,n4[5] ,n26[5]);
    xnor g4848(n4294 ,n4[4] ,n26[4]);
    xnor g4849(n4293 ,n4[1] ,n26[1]);
    xnor g4850(n4292 ,n4[6] ,n26[6]);
    xnor g4851(n4291 ,n4[7] ,n26[7]);
    nor g4852(n4290 ,n4274 ,n4278);
    nor g4853(n4289 ,n4275 ,n4272);
    nor g4854(n4288 ,n4273 ,n4281);
    nor g4855(n4287 ,n4276 ,n4277);
    nor g4856(n4286 ,n4279 ,n4280);
    nor g4857(n4285 ,n26[0] ,n4[0]);
    nor g4858(n4284 ,n26[6] ,n4[6]);
    nor g4859(n4283 ,n26[7] ,n4[7]);
    nor g4860(n4282 ,n26[1] ,n4[1]);
    not g4861(n4281 ,n4[4]);
    not g4862(n4280 ,n4[3]);
    not g4863(n4279 ,n26[3]);
    not g4864(n4278 ,n4[5]);
    not g4865(n4277 ,n4[0]);
    not g4866(n4276 ,n26[0]);
    not g4867(n4275 ,n26[2]);
    not g4868(n4274 ,n26[5]);
    not g4869(n4273 ,n26[4]);
    not g4870(n4272 ,n4[2]);
    xor g4871(n4579 ,n4339 ,n4382);
    nor g4872(n4382 ,n4333 ,n4381);
    xor g4873(n4578 ,n4352 ,n4380);
    nor g4874(n4381 ,n4352 ,n4380);
    nor g4875(n4380 ,n4334 ,n4379);
    xor g4876(n4577 ,n4353 ,n4378);
    nor g4877(n4379 ,n4353 ,n4378);
    nor g4878(n4378 ,n4336 ,n4377);
    xor g4879(n4576 ,n4351 ,n4376);
    nor g4880(n4377 ,n4351 ,n4376);
    nor g4881(n4376 ,n4337 ,n4375);
    xnor g4882(n4575 ,n4350 ,n4373);
    nor g4883(n4375 ,n4350 ,n4374);
    not g4884(n4374 ,n4373);
    nor g4885(n4373 ,n4326 ,n4372);
    xnor g4886(n4629 ,n4347 ,n4371);
    nor g4887(n4372 ,n4347 ,n4371);
    nor g4888(n4371 ,n4327 ,n4370);
    xnor g4889(n4630 ,n4343 ,n4369);
    nor g4890(n4370 ,n4343 ,n4369);
    nor g4891(n4369 ,n4332 ,n4368);
    xnor g4892(n4631 ,n4340 ,n4367);
    nor g4893(n4368 ,n4340 ,n4367);
    nor g4894(n4367 ,n4323 ,n4366);
    xnor g4895(n4632 ,n4341 ,n4365);
    nor g4896(n4366 ,n4341 ,n4365);
    nor g4897(n4365 ,n4331 ,n4364);
    xnor g4898(n4633 ,n4349 ,n4363);
    nor g4899(n4364 ,n4349 ,n4363);
    nor g4900(n4363 ,n4335 ,n4362);
    xnor g4901(n4634 ,n4348 ,n4361);
    nor g4902(n4362 ,n4348 ,n4361);
    nor g4903(n4361 ,n4329 ,n4360);
    xnor g4904(n4635 ,n4342 ,n4359);
    nor g4905(n4360 ,n4342 ,n4359);
    nor g4906(n4359 ,n4324 ,n4358);
    xnor g4907(n4636 ,n4345 ,n4357);
    nor g4908(n4358 ,n4345 ,n4357);
    nor g4909(n4357 ,n4328 ,n4356);
    xnor g4910(n4637 ,n4344 ,n4355);
    nor g4911(n4356 ,n4344 ,n4355);
    nor g4912(n4355 ,n4325 ,n4354);
    xnor g4913(n4638 ,n4346 ,n4338);
    nor g4914(n4354 ,n4338 ,n4346);
    nor g4915(n4639 ,n4338 ,n4330);
    xnor g4916(n4353 ,n4617 ,n4601);
    xnor g4917(n4352 ,n4618 ,n4602);
    xnor g4918(n4351 ,n4616 ,n4600);
    xnor g4919(n4350 ,n4615 ,n4599);
    xnor g4920(n4349 ,n4610 ,n4594);
    xnor g4921(n4348 ,n4609 ,n4593);
    xnor g4922(n4347 ,n4614 ,n4598);
    xnor g4923(n4346 ,n4589 ,n4605);
    xnor g4924(n4345 ,n4607 ,n4591);
    xnor g4925(n4344 ,n4606 ,n4590);
    xnor g4926(n4343 ,n4613 ,n4597);
    xnor g4927(n4342 ,n4608 ,n4592);
    xnor g4928(n4341 ,n4611 ,n4595);
    xnor g4929(n4340 ,n4612 ,n4596);
    xnor g4930(n4339 ,n4619 ,n4603);
    nor g4931(n4337 ,n4319 ,n4318);
    nor g4932(n4336 ,n4316 ,n4322);
    nor g4933(n4335 ,n4609 ,n4593);
    nor g4934(n4334 ,n4314 ,n4321);
    nor g4935(n4333 ,n4313 ,n4315);
    nor g4936(n4332 ,n4612 ,n4596);
    nor g4937(n4331 ,n4610 ,n4594);
    nor g4938(n4338 ,n4320 ,n4317);
    nor g4939(n4330 ,n4604 ,n4588);
    nor g4940(n4329 ,n4608 ,n4592);
    nor g4941(n4328 ,n4606 ,n4590);
    nor g4942(n4327 ,n4613 ,n4597);
    nor g4943(n4326 ,n4614 ,n4598);
    nor g4944(n4325 ,n4605 ,n4589);
    nor g4945(n4324 ,n4607 ,n4591);
    nor g4946(n4323 ,n4611 ,n4595);
    not g4947(n4322 ,n4600);
    not g4948(n4321 ,n4601);
    not g4949(n4320 ,n4604);
    not g4950(n4319 ,n4615);
    not g4951(n4318 ,n4599);
    not g4952(n4317 ,n4588);
    not g4953(n4316 ,n4616);
    not g4954(n4315 ,n4602);
    not g4955(n4314 ,n4617);
    not g4956(n4313 ,n4618);
    not g4957(n2316 ,n27[0]);
endmodule
