module top (n0, n1, n2, n3, n4, n5, n6, n8, n9, n7, n10, n11, n12, n13, n14, n15);
    input n0, n1;
    input [7:0] n2, n3, n4, n5, n6, n7;
    input [2:0] n8;
    input [3:0] n9;
    output [15:0] n10, n11, n12, n13, n14;
    output [7:0] n15;
    wire n0, n1;
    wire [7:0] n2, n3, n4, n5, n6, n7;
    wire [2:0] n8;
    wire [3:0] n9;
    wire [15:0] n10, n11, n12, n13, n14;
    wire [7:0] n15;
    wire [15:0] n16;
    wire [15:0] n17;
    wire [3:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [15:0] n23;
    wire [15:0] n24;
    wire [7:0] n25;
    wire [2:0] n26;
    wire [15:0] n27;
    wire [15:0] n28;
    wire [15:0] n29;
    wire [15:0] n30;
    wire [15:0] n31;
    wire [15:0] n32;
    wire [7:0] n33;
    wire [15:0] n34;
    wire [15:0] n35;
    wire [15:0] n36;
    wire [7:0] n37;
    wire [15:0] n38;
    wire [15:0] n39;
    wire [15:0] n40;
    wire [15:0] n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310, n311, n312, n313;
    wire n314, n315, n316, n317, n318, n319, n320, n321;
    wire n322, n323, n324, n325, n326, n327, n328, n329;
    wire n330, n331, n332, n333, n334, n335, n336, n337;
    wire n338, n339, n340, n341, n342, n343, n344, n345;
    wire n346, n347, n348, n349, n350, n351, n352, n353;
    wire n354, n355, n356, n357, n358, n359, n360, n361;
    wire n362, n363, n364, n365, n366, n367, n368, n369;
    wire n370, n371, n372, n373, n374, n375, n376, n377;
    wire n378, n379, n380, n381, n382, n383, n384, n385;
    wire n386, n387, n388, n389, n390, n391, n392, n393;
    wire n394, n395, n396, n397, n398, n399, n400, n401;
    wire n402, n403, n404, n405, n406, n407, n408, n409;
    wire n410, n411, n412, n413, n414, n415, n416, n417;
    wire n418, n419, n420, n421, n422, n423, n424, n425;
    wire n426, n427, n428, n429, n430, n431, n432, n433;
    wire n434, n435, n436, n437, n438, n439, n440, n441;
    wire n442, n443, n444, n445, n446, n447, n448, n449;
    wire n450, n451, n452, n453, n454, n455, n456, n457;
    wire n458, n459, n460, n461, n462, n463, n464, n465;
    wire n466, n467, n468, n469, n470, n471, n472, n473;
    wire n474, n475, n476, n477, n478, n479, n480, n481;
    wire n482, n483, n484, n485, n486, n487, n488, n489;
    wire n490, n491, n492, n493, n494, n495, n496, n497;
    wire n498, n499, n500, n501, n502, n503, n504, n505;
    wire n506, n507, n508, n509, n510, n511, n512, n513;
    wire n514, n515, n516, n517, n518, n519, n520, n521;
    wire n522, n523, n524, n525, n526, n527, n528, n529;
    wire n530, n531, n532, n533, n534, n535, n536, n537;
    wire n538, n539, n540, n541, n542, n543, n544, n545;
    wire n546, n547, n548, n549, n550, n551, n552, n553;
    wire n554, n555, n556, n557, n558, n559, n560, n561;
    wire n562, n563, n564, n565, n566, n567, n568, n569;
    wire n570, n571, n572, n573, n574, n575, n576, n577;
    wire n578, n579, n580, n581, n582, n583, n584, n585;
    wire n586, n587, n588, n589, n590, n591, n592, n593;
    wire n594, n595, n596, n597, n598, n599, n600, n601;
    wire n602, n603, n604, n605, n606, n607, n608, n609;
    wire n610, n611, n612, n613, n614, n615, n616, n617;
    wire n618, n619, n620, n621, n622, n623, n624, n625;
    wire n626, n627, n628, n629, n630, n631, n632, n633;
    wire n634, n635, n636, n637, n638, n639, n640, n641;
    wire n642, n643, n644, n645, n646, n647, n648, n649;
    wire n650, n651, n652, n653, n654, n655, n656, n657;
    wire n658, n659, n660, n661, n662, n663, n664, n665;
    wire n666, n667, n668, n669, n670, n671, n672, n673;
    wire n674, n675, n676, n677, n678, n679, n680, n681;
    wire n682, n683, n684, n685, n686, n687, n688, n689;
    wire n690, n691, n692, n693, n694, n695, n696, n697;
    wire n698, n699, n700, n701, n702, n703, n704, n705;
    wire n706, n707, n708, n709, n710, n711, n712, n713;
    wire n714, n715, n716, n717, n718, n719, n720, n721;
    wire n722, n723, n724, n725, n726, n727, n728, n729;
    wire n730, n731, n732, n733, n734, n735, n736, n737;
    wire n738, n739, n740, n741, n742, n743, n744, n745;
    wire n746, n747, n748, n749, n750, n751, n752, n753;
    wire n754, n755, n756, n757, n758, n759, n760, n761;
    wire n762, n763, n764, n765, n766, n767, n768, n769;
    wire n770, n771, n772, n773, n774, n775, n776, n777;
    wire n778, n779, n780, n781, n782, n783, n784, n785;
    wire n786, n787, n788, n789, n790, n791, n792, n793;
    wire n794, n795, n796, n797, n798, n799, n800, n801;
    wire n802, n803, n804, n805, n806, n807, n808, n809;
    wire n810, n811, n812, n813, n814, n815, n816, n817;
    wire n818, n819, n820, n821, n822, n823, n824, n825;
    wire n826, n827, n828, n829, n830, n831, n832, n833;
    wire n834, n835, n836, n837, n838, n839, n840, n841;
    wire n842, n843, n844, n845, n846, n847, n848, n849;
    wire n850, n851, n852, n853, n854, n855, n856, n857;
    wire n858, n859, n860, n861, n862, n863, n864, n865;
    wire n866, n867, n868, n869, n870, n871, n872, n873;
    wire n874, n875, n876, n877, n878, n879, n880, n881;
    wire n882, n883, n884, n885, n886, n887, n888, n889;
    wire n890, n891, n892, n893, n894, n895, n896, n897;
    wire n898, n899, n900, n901, n902, n903, n904, n905;
    wire n906, n907, n908, n909, n910, n911, n912, n913;
    wire n914, n915, n916, n917, n918, n919, n920, n921;
    wire n922, n923, n924, n925, n926, n927, n928, n929;
    wire n930, n931, n932, n933, n934, n935, n936, n937;
    wire n938, n939, n940, n941, n942, n943, n944, n945;
    wire n946, n947, n948, n949, n950, n951, n952, n953;
    wire n954, n955, n956, n957, n958, n959, n960, n961;
    wire n962, n963, n964, n965, n966, n967, n968, n969;
    wire n970, n971, n972, n973, n974, n975, n976, n977;
    wire n978, n979, n980, n981, n982, n983, n984, n985;
    wire n986, n987, n988, n989, n990, n991, n992, n993;
    wire n994, n995, n996, n997, n998, n999, n1000, n1001;
    wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
    wire n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
    wire n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
    wire n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
    wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
    wire n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049;
    wire n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
    wire n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065;
    wire n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
    wire n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081;
    wire n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089;
    wire n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097;
    wire n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105;
    wire n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113;
    wire n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121;
    wire n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129;
    wire n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137;
    wire n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145;
    wire n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153;
    wire n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161;
    wire n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169;
    wire n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177;
    wire n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185;
    wire n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193;
    wire n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201;
    wire n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209;
    wire n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217;
    wire n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225;
    wire n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;
    wire n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241;
    wire n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249;
    wire n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257;
    wire n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265;
    wire n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273;
    wire n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281;
    wire n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289;
    wire n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297;
    wire n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305;
    wire n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313;
    wire n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321;
    wire n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329;
    wire n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337;
    wire n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345;
    wire n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353;
    wire n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;
    wire n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369;
    wire n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377;
    wire n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385;
    wire n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393;
    wire n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401;
    wire n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409;
    wire n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417;
    wire n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425;
    wire n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433;
    wire n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441;
    wire n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449;
    wire n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457;
    wire n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465;
    wire n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473;
    wire n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481;
    wire n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
    wire n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497;
    wire n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505;
    wire n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513;
    wire n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
    wire n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529;
    wire n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537;
    wire n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545;
    wire n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553;
    wire n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561;
    wire n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569;
    wire n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577;
    wire n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585;
    wire n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593;
    wire n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601;
    wire n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609;
    wire n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617;
    wire n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625;
    wire n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633;
    wire n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641;
    wire n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649;
    wire n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657;
    wire n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665;
    wire n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673;
    wire n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681;
    wire n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689;
    wire n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
    wire n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705;
    wire n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713;
    wire n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721;
    wire n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729;
    wire n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737;
    wire n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745;
    wire n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753;
    wire n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761;
    wire n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769;
    wire n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777;
    wire n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785;
    wire n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793;
    wire n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801;
    wire n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809;
    wire n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817;
    wire n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825;
    wire n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833;
    wire n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;
    wire n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849;
    wire n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857;
    wire n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865;
    wire n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873;
    wire n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881;
    wire n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889;
    wire n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897;
    wire n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905;
    wire n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913;
    wire n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921;
    wire n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929;
    wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
    wire n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945;
    wire n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953;
    wire n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961;
    wire n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969;
    wire n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977;
    wire n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985;
    wire n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993;
    wire n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001;
    wire n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009;
    wire n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017;
    wire n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025;
    wire n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033;
    wire n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041;
    wire n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049;
    wire n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057;
    wire n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065;
    wire n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073;
    wire n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081;
    wire n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089;
    wire n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097;
    wire n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105;
    wire n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113;
    wire n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121;
    wire n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129;
    wire n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137;
    wire n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145;
    wire n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153;
    wire n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161;
    wire n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169;
    wire n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177;
    wire n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185;
    wire n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193;
    wire n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201;
    wire n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209;
    wire n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217;
    wire n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225;
    wire n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233;
    wire n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241;
    wire n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
    wire n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257;
    wire n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265;
    wire n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273;
    wire n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281;
    wire n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289;
    wire n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297;
    wire n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305;
    wire n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313;
    wire n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321;
    wire n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329;
    wire n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337;
    wire n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345;
    wire n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353;
    wire n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361;
    wire n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369;
    wire n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377;
    wire n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385;
    wire n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
    wire n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401;
    wire n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409;
    wire n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417;
    wire n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425;
    wire n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433;
    wire n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441;
    wire n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449;
    wire n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457;
    wire n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465;
    wire n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473;
    wire n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481;
    wire n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489;
    wire n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497;
    wire n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505;
    wire n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513;
    wire n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521;
    wire n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529;
    wire n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537;
    wire n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545;
    wire n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553;
    wire n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561;
    wire n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569;
    wire n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577;
    wire n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585;
    wire n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593;
    wire n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601;
    wire n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609;
    wire n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617;
    wire n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625;
    wire n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633;
    wire n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641;
    wire n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649;
    wire n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657;
    wire n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665;
    wire n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673;
    wire n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681;
    wire n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689;
    wire n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697;
    wire n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705;
    wire n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713;
    wire n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721;
    wire n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729;
    wire n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737;
    wire n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745;
    wire n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753;
    wire n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761;
    wire n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769;
    wire n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777;
    wire n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785;
    wire n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793;
    wire n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
    wire n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809;
    wire n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817;
    wire n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825;
    wire n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833;
    wire n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841;
    wire n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849;
    wire n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857;
    wire n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865;
    wire n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873;
    wire n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881;
    wire n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889;
    wire n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897;
    wire n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905;
    wire n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913;
    wire n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921;
    wire n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929;
    wire n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937;
    wire n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945;
    wire n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953;
    wire n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961;
    wire n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969;
    wire n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977;
    wire n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985;
    wire n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993;
    wire n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001;
    wire n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009;
    wire n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017;
    wire n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025;
    wire n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033;
    wire n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041;
    wire n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049;
    wire n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057;
    wire n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065;
    wire n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073;
    wire n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081;
    wire n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089;
    wire n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097;
    wire n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105;
    wire n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113;
    wire n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121;
    wire n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129;
    wire n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137;
    wire n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145;
    wire n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153;
    wire n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161;
    wire n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169;
    wire n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177;
    wire n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185;
    wire n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193;
    wire n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201;
    wire n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209;
    wire n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217;
    wire n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225;
    wire n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233;
    wire n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241;
    wire n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249;
    wire n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257;
    wire n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265;
    wire n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273;
    wire n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281;
    wire n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289;
    wire n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297;
    wire n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305;
    wire n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313;
    wire n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321;
    wire n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329;
    wire n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337;
    wire n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345;
    wire n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353;
    wire n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361;
    wire n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369;
    wire n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377;
    wire n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385;
    wire n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393;
    wire n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401;
    wire n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409;
    wire n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417;
    wire n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425;
    wire n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433;
    wire n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441;
    wire n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449;
    wire n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457;
    wire n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465;
    wire n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473;
    wire n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481;
    wire n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489;
    wire n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497;
    wire n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505;
    wire n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513;
    wire n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521;
    wire n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529;
    wire n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537;
    wire n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545;
    wire n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553;
    wire n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561;
    wire n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569;
    wire n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577;
    wire n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585;
    wire n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593;
    wire n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601;
    wire n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609;
    wire n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617;
    wire n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625;
    wire n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633;
    wire n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641;
    wire n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649;
    wire n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657;
    wire n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665;
    wire n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673;
    wire n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681;
    wire n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689;
    wire n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697;
    wire n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705;
    wire n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713;
    wire n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721;
    wire n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729;
    wire n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737;
    wire n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745;
    wire n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753;
    wire n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761;
    wire n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769;
    wire n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777;
    wire n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785;
    wire n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793;
    wire n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801;
    wire n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809;
    wire n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817;
    wire n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825;
    wire n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833;
    wire n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841;
    wire n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849;
    wire n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857;
    wire n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865;
    wire n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873;
    wire n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881;
    wire n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889;
    wire n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897;
    wire n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905;
    wire n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913;
    wire n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921;
    wire n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929;
    wire n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937;
    wire n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945;
    wire n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953;
    wire n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961;
    wire n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969;
    wire n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977;
    wire n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985;
    wire n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993;
    wire n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001;
    wire n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009;
    wire n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017;
    wire n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025;
    wire n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033;
    wire n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041;
    wire n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049;
    wire n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057;
    wire n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065;
    wire n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073;
    wire n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081;
    wire n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089;
    wire n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097;
    wire n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105;
    wire n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113;
    wire n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121;
    wire n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129;
    wire n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137;
    wire n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145;
    wire n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153;
    wire n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161;
    wire n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169;
    wire n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177;
    wire n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185;
    wire n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193;
    wire n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201;
    wire n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209;
    wire n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217;
    wire n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225;
    wire n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233;
    wire n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241;
    wire n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249;
    wire n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257;
    wire n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265;
    wire n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273;
    wire n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281;
    wire n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289;
    wire n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297;
    wire n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305;
    wire n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313;
    wire n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321;
    wire n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329;
    wire n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337;
    wire n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345;
    wire n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353;
    wire n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361;
    wire n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369;
    wire n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377;
    wire n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385;
    wire n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393;
    wire n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401;
    wire n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409;
    wire n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417;
    wire n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425;
    wire n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433;
    wire n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441;
    wire n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449;
    wire n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457;
    wire n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465;
    wire n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473;
    wire n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481;
    wire n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489;
    wire n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497;
    wire n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505;
    wire n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513;
    wire n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521;
    wire n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529;
    wire n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537;
    wire n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545;
    wire n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553;
    wire n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561;
    wire n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569;
    wire n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577;
    wire n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585;
    wire n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593;
    wire n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601;
    wire n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609;
    wire n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617;
    wire n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625;
    wire n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633;
    wire n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641;
    wire n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649;
    wire n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657;
    wire n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665;
    wire n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673;
    wire n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681;
    wire n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689;
    wire n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697;
    wire n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705;
    wire n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713;
    wire n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721;
    wire n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729;
    wire n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737;
    wire n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745;
    wire n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753;
    wire n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761;
    wire n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769;
    wire n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777;
    wire n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785;
    wire n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793;
    wire n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801;
    wire n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809;
    wire n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817;
    wire n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825;
    wire n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833;
    wire n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841;
    wire n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849;
    wire n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857;
    wire n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865;
    wire n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873;
    wire n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881;
    wire n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889;
    wire n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897;
    wire n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905;
    wire n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913;
    wire n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921;
    wire n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929;
    wire n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937;
    wire n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945;
    wire n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953;
    wire n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961;
    wire n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969;
    wire n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977;
    wire n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985;
    wire n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993;
    wire n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001;
    wire n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009;
    wire n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017;
    wire n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025;
    wire n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033;
    wire n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041;
    wire n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049;
    wire n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057;
    wire n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065;
    wire n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073;
    wire n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081;
    wire n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089;
    wire n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097;
    wire n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105;
    wire n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113;
    wire n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121;
    wire n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129;
    wire n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137;
    wire n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145;
    wire n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153;
    wire n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161;
    wire n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169;
    wire n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177;
    wire n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185;
    wire n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193;
    wire n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201;
    wire n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209;
    wire n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217;
    wire n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225;
    wire n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233;
    wire n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241;
    wire n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249;
    wire n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257;
    wire n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265;
    wire n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273;
    wire n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281;
    wire n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289;
    wire n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297;
    wire n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305;
    wire n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313;
    wire n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321;
    wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
    wire n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337;
    wire n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345;
    wire n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353;
    wire n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361;
    wire n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369;
    wire n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377;
    wire n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385;
    wire n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393;
    wire n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401;
    wire n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409;
    wire n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417;
    wire n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425;
    wire n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433;
    wire n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441;
    wire n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449;
    wire n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457;
    wire n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465;
    wire n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473;
    wire n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481;
    wire n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489;
    wire n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497;
    wire n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505;
    wire n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513;
    wire n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521;
    wire n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529;
    wire n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537;
    wire n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545;
    wire n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553;
    wire n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561;
    wire n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569;
    wire n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577;
    wire n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585;
    wire n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593;
    wire n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601;
    wire n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609;
    wire n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617;
    wire n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625;
    wire n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633;
    wire n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641;
    wire n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649;
    wire n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657;
    wire n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665;
    wire n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673;
    wire n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681;
    wire n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689;
    wire n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697;
    wire n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705;
    wire n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713;
    wire n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721;
    wire n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729;
    wire n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737;
    wire n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745;
    wire n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753;
    wire n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761;
    wire n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769;
    wire n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777;
    wire n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785;
    wire n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793;
    wire n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801;
    wire n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809;
    wire n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817;
    wire n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825;
    wire n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833;
    wire n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841;
    wire n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849;
    wire n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857;
    wire n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865;
    wire n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873;
    wire n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881;
    wire n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889;
    wire n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897;
    wire n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905;
    wire n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913;
    wire n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921;
    wire n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929;
    wire n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937;
    wire n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945;
    wire n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953;
    wire n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961;
    wire n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969;
    wire n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977;
    wire n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985;
    wire n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993;
    wire n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001;
    wire n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009;
    wire n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017;
    wire n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025;
    wire n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033;
    wire n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041;
    wire n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049;
    wire n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057;
    wire n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065;
    wire n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073;
    wire n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081;
    wire n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089;
    wire n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097;
    wire n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105;
    wire n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113;
    wire n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121;
    wire n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129;
    wire n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137;
    wire n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145;
    wire n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153;
    wire n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161;
    wire n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169;
    wire n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177;
    wire n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185;
    wire n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193;
    wire n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201;
    wire n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209;
    wire n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217;
    wire n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225;
    wire n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233;
    wire n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241;
    wire n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249;
    wire n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257;
    wire n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265;
    wire n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273;
    wire n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281;
    wire n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289;
    wire n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297;
    wire n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305;
    wire n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313;
    wire n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321;
    wire n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329;
    wire n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337;
    wire n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345;
    wire n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353;
    wire n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361;
    wire n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369;
    wire n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377;
    wire n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385;
    wire n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393;
    wire n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401;
    wire n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409;
    wire n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417;
    wire n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425;
    wire n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433;
    wire n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441;
    wire n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449;
    wire n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457;
    wire n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465;
    wire n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473;
    wire n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481;
    wire n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489;
    wire n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497;
    wire n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505;
    wire n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513;
    wire n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521;
    wire n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529;
    wire n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537;
    wire n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545;
    wire n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553;
    wire n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561;
    wire n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569;
    wire n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577;
    wire n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585;
    wire n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593;
    wire n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601;
    wire n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609;
    wire n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617;
    wire n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625;
    wire n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633;
    wire n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641;
    wire n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649;
    wire n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657;
    wire n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665;
    wire n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673;
    wire n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681;
    wire n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689;
    wire n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697;
    wire n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705;
    wire n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713;
    wire n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721;
    wire n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729;
    wire n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737;
    wire n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745;
    wire n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753;
    wire n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761;
    wire n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769;
    wire n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777;
    wire n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785;
    wire n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793;
    wire n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801;
    wire n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809;
    wire n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817;
    wire n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825;
    wire n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833;
    wire n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841;
    wire n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849;
    wire n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857;
    wire n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865;
    wire n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873;
    wire n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881;
    wire n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889;
    wire n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897;
    wire n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905;
    wire n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913;
    wire n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921;
    wire n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929;
    wire n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937;
    wire n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945;
    wire n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953;
    wire n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961;
    wire n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969;
    wire n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977;
    wire n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985;
    wire n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993;
    wire n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001;
    wire n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009;
    wire n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017;
    wire n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025;
    wire n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033;
    wire n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041;
    wire n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049;
    wire n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057;
    wire n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065;
    wire n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073;
    wire n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081;
    wire n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089;
    wire n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097;
    wire n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105;
    wire n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113;
    wire n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121;
    wire n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129;
    wire n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137;
    wire n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145;
    wire n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153;
    wire n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161;
    wire n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169;
    wire n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177;
    wire n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185;
    wire n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193;
    wire n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201;
    wire n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209;
    wire n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217;
    wire n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225;
    wire n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233;
    wire n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241;
    wire n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249;
    wire n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257;
    wire n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265;
    wire n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273;
    wire n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281;
    wire n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289;
    wire n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297;
    wire n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305;
    wire n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313;
    wire n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321;
    wire n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329;
    wire n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337;
    wire n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345;
    wire n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353;
    wire n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361;
    wire n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369;
    wire n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377;
    wire n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385;
    wire n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393;
    wire n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401;
    wire n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409;
    wire n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417;
    wire n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425;
    wire n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433;
    wire n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441;
    wire n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449;
    wire n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457;
    wire n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465;
    wire n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473;
    wire n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481;
    wire n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489;
    wire n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497;
    wire n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505;
    wire n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513;
    wire n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521;
    wire n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529;
    wire n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537;
    wire n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545;
    wire n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553;
    wire n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561;
    wire n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569;
    wire n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577;
    wire n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585;
    wire n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593;
    wire n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601;
    wire n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609;
    wire n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617;
    wire n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625;
    wire n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633;
    wire n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641;
    wire n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649;
    wire n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657;
    wire n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665;
    wire n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673;
    wire n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681;
    wire n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689;
    wire n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697;
    wire n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705;
    wire n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713;
    wire n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721;
    wire n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729;
    wire n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737;
    wire n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745;
    wire n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753;
    wire n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761;
    wire n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769;
    wire n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777;
    wire n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785;
    wire n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793;
    wire n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801;
    wire n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809;
    wire n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817;
    wire n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825;
    wire n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833;
    wire n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841;
    wire n7842, n7843, n7844, n7845, n7846;
    not g0(n3436 ,n3435);
    nor g1(n4486 ,n4349 ,n4407);
    nor g2(n6550 ,n6372 ,n6448);
    nor g3(n2622 ,n2545 ,n2591);
    not g4(n6641 ,n6640);
    nor g5(n4143 ,n4007 ,n4024);
    nor g6(n4174 ,n4013 ,n4007);
    xnor g7(n5003 ,n4957 ,n4918);
    not g8(n1969 ,n1970);
    xnor g9(n6283 ,n5974 ,n5994);
    nor g10(n4657 ,n4469 ,n4544);
    or g11(n1773 ,n1410 ,n1500);
    xnor g12(n3898 ,n41[5] ,n7806);
    nor g13(n3116 ,n3013 ,n3037);
    nor g14(n3915 ,n3883 ,n3914);
    not g15(n502 ,n501);
    dff g16(.RN(n1), .SN(1'b1), .CK(n0), .D(n1742), .Q(n30[1]));
    nor g17(n2353 ,n2261 ,n2325);
    not g18(n884 ,n31[4]);
    or g19(n5539 ,n5098 ,n5109);
    nor g20(n7315 ,n7304 ,n7314);
    nor g21(n6454 ,n6093 ,n6330);
    not g22(n3163 ,n3162);
    nor g23(n4641 ,n4463 ,n4528);
    xnor g24(n6403 ,n6154 ,n6152);
    not g25(n809 ,n27[4]);
    nor g26(n5607 ,n5264 ,n5440);
    xnor g27(n4900 ,n4820 ,n4733);
    nor g28(n5206 ,n5088 ,n5119);
    not g29(n4666 ,n4665);
    nor g30(n511 ,n436 ,n482);
    not g31(n4925 ,n4924);
    not g32(n3215 ,n3214);
    not g33(n7242 ,n7241);
    not g34(n745 ,n1874);
    nor g35(n7459 ,n41[7] ,n7821);
    xnor g36(n7812 ,n2406 ,n2414);
    xnor g37(n6183 ,n5782 ,n5530);
    or g38(n7638 ,n7534 ,n7543);
    not g39(n2248 ,n2247);
    nor g40(n4329 ,n4167 ,n4069);
    nor g41(n3560 ,n3526 ,n3532);
    not g42(n4219 ,n4218);
    xnor g43(n3076 ,n40[13] ,n7752);
    or g44(n3038 ,n3000 ,n3001);
    nor g45(n5573 ,n5108 ,n5106);
    xnor g46(n4606 ,n4474 ,n4499);
    nor g47(n7013 ,n6924 ,n6941);
    or g48(n1585 ,n1246 ,n1110);
    or g49(n7693 ,n7625 ,n7640);
    nor g50(n7558 ,n7418 ,n7478);
    not g51(n948 ,n29[6]);
    nor g52(n117 ,n102 ,n115);
    xor g53(n4371 ,n4244 ,n4044);
    or g54(n7662 ,n7594 ,n7593);
    xor g55(n5798 ,n5539 ,n5148);
    nor g56(n2743 ,n2697 ,n2698);
    nor g57(n1355 ,n853 ,n636);
    not g58(n3006 ,n7746);
    nor g59(n316 ,n170 ,n240);
    nor g60(n2922 ,n2878 ,n2892);
    not g61(n4195 ,n4194);
    not g62(n406 ,n405);
    or g63(n1728 ,n1369 ,n1178);
    nor g64(n5619 ,n5172 ,n5356);
    nor g65(n7304 ,n7299 ,n7290);
    nor g66(n2755 ,n2666 ,n2717);
    nor g67(n1159 ,n1102 ,n1077);
    nor g68(n2087 ,n2015 ,n2040);
    nor g69(n572 ,n541 ,n553);
    nor g70(n7281 ,n7261 ,n7251);
    xnor g71(n3401 ,n3329 ,n3152);
    nor g72(n5190 ,n5088 ,n5102);
    not g73(n831 ,n23[5]);
    or g74(n7615 ,n7596 ,n7587);
    nor g75(n5297 ,n5103 ,n5094);
    nor g76(n5005 ,n4916 ,n4976);
    not g77(n5103 ,n21[1]);
    not g78(n6107 ,n6106);
    xnor g79(n7106 ,n6998 ,n7046);
    not g80(n7215 ,n7214);
    xnor g81(n2810 ,n2736 ,n2710);
    not g82(n7084 ,n7083);
    not g83(n878 ,n21[5]);
    nor g84(n622 ,n599 ,n621);
    nor g85(n621 ,n606 ,n620);
    nor g86(n557 ,n517 ,n530);
    not g87(n2323 ,n2322);
    nor g88(n4510 ,n4317 ,n4448);
    or g89(n93 ,n33[1] ,n91);
    nor g90(n7008 ,n6869 ,n6939);
    not g91(n6570 ,n6569);
    not g92(n2699 ,n2698);
    nor g93(n571 ,n542 ,n557);
    xnor g94(n2773 ,n2694 ,n2720);
    xnor g95(n2856 ,n2781 ,n2702);
    xnor g96(n3789 ,n3727 ,n3703);
    nor g97(n1955 ,n1902 ,n1937);
    nor g98(n394 ,n298 ,n357);
    nor g99(n3369 ,n3313 ,n3358);
    not g100(n2714 ,n2713);
    nor g101(n624 ,n615 ,n623);
    nor g102(n5651 ,n5414 ,n5130);
    nor g103(n2020 ,n1903 ,n1982);
    or g104(n7633 ,n7600 ,n7513);
    not g105(n773 ,n4[7]);
    not g106(n805 ,n6[1]);
    nor g107(n2952 ,n2927 ,n2933);
    nor g108(n6661 ,n6488 ,n6557);
    not g109(n5277 ,n5276);
    nor g110(n1430 ,n684 ,n638);
    nor g111(n4413 ,n4080 ,n4353);
    not g112(n6639 ,n6638);
    nor g113(n259 ,n156 ,n153);
    not g114(n6793 ,n6792);
    dff g115(.RN(n1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n22[1]));
    not g116(n3209 ,n3208);
    xnor g117(n4785 ,n4673 ,n4691);
    not g118(n149 ,n19[2]);
    nor g119(n561 ,n502 ,n522);
    nor g120(n1551 ,n938 ,n1100);
    xor g121(n7780 ,n4767 ,n4711);
    nor g122(n3683 ,n3627 ,n3636);
    not g123(n3595 ,n7784);
    nor g124(n2370 ,n2312 ,n2358);
    not g125(n885 ,n21[3]);
    nor g126(n2488 ,n2442 ,n2477);
    nor g127(n5670 ,n5265 ,n5441);
    nor g128(n7494 ,n7362 ,n7475);
    nor g129(n6483 ,n6013 ,n6363);
    not g130(n5112 ,n22[2]);
    not g131(n6153 ,n6152);
    not g132(n688 ,n32[7]);
    nor g133(n7551 ,n7435 ,n7481);
    not g134(n5463 ,n5462);
    nor g135(n2615 ,n2444 ,n2549);
    xnor g136(n3843 ,n37[7] ,n19[7]);
    nor g137(n7321 ,n7320 ,n7284);
    nor g138(n1431 ,n932 ,n637);
    xnor g139(n6722 ,n6515 ,n6581);
    xnor g140(n7083 ,n6975 ,n6883);
    not g141(n6826 ,n6825);
    not g142(n2964 ,n2963);
    dff g143(.RN(n1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n23[0]));
    or g144(n7696 ,n7645 ,n7642);
    nor g145(n1328 ,n944 ,n642);
    xnor g146(n3074 ,n40[0] ,n7739);
    not g147(n675 ,n36[9]);
    nor g148(n3575 ,n3530 ,n3574);
    nor g149(n2091 ,n2024 ,n2044);
    nor g150(n7294 ,n7278 ,n7276);
    nor g151(n1484 ,n793 ,n639);
    or g152(n979 ,n18[0] ,n18[1]);
    nor g153(n4188 ,n4020 ,n4028);
    xnor g154(n7030 ,n6913 ,n6835);
    nor g155(n3916 ,n3889 ,n3915);
    nor g156(n1227 ,n827 ,n642);
    nor g157(n1119 ,n635 ,n1053);
    nor g158(n3229 ,n3044 ,n3130);
    nor g159(n6666 ,n6130 ,n6535);
    nor g160(n559 ,n484 ,n526);
    nor g161(n3944 ,n3935 ,n3932);
    nor g162(n6675 ,n6328 ,n6512);
    xnor g163(n2845 ,n2780 ,n2730);
    nor g164(n5142 ,n5095 ,n5110);
    xnor g165(n1981 ,n1959 ,n1951);
    nor g166(n2410 ,n2409 ,n2361);
    not g167(n2296 ,n2295);
    xnor g168(n6856 ,n6720 ,n6548);
    not g169(n4816 ,n4815);
    nor g170(n1998 ,n1890 ,n1978);
    not g171(n2576 ,n2575);
    nor g172(n1128 ,n635 ,n1097);
    nor g173(n2623 ,n2532 ,n2592);
    not g174(n5375 ,n5374);
    buf g175(n13[0], n10[0]);
    not g176(n4360 ,n4359);
    nor g177(n6725 ,n6549 ,n6688);
    xor g178(n5772 ,n5303 ,n5250);
    xnor g179(n1979 ,n1883 ,n1960);
    nor g180(n1312 ,n698 ,n637);
    not g181(n2346 ,n2345);
    nor g182(n5635 ,n5162 ,n5266);
    nor g183(n7196 ,n7132 ,n7171);
    or g184(n1628 ,n1295 ,n1493);
    nor g185(n3261 ,n3094 ,n3175);
    xor g186(n5801 ,n5335 ,n5274);
    xor g187(n6405 ,n6176 ,n6134);
    not g188(n3014 ,n7740);
    nor g189(n6702 ,n6362 ,n6553);
    nor g190(n2879 ,n2824 ,n2853);
    nor g191(n4332 ,n4203 ,n4049);
    not g192(n3602 ,n7810);
    not g193(n4504 ,n4503);
    nor g194(n5440 ,n5098 ,n5110);
    not g195(n5199 ,n5198);
    dff g196(.RN(n1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n17[1]));
    xnor g197(n6154 ,n5798 ,n5280);
    nor g198(n2463 ,n2440 ,n2439);
    nor g199(n2619 ,n2571 ,n2614);
    not g200(n158 ,n19[3]);
    xnor g201(n4869 ,n4772 ,n4758);
    or g202(n7647 ,n7588 ,n7559);
    nor g203(n7532 ,n7365 ,n7477);
    xnor g204(n2222 ,n2155 ,n2123);
    nor g205(n1952 ,n1929 ,n1923);
    not g206(n6615 ,n6614);
    nor g207(n1556 ,n934 ,n1100);
    nor g208(n1298 ,n952 ,n1101);
    xnor g209(n3329 ,n3120 ,n3266);
    nor g210(n1986 ,n1901 ,n1976);
    nor g211(n2185 ,n2106 ,n2164);
    not g212(n7201 ,n7200);
    nor g213(n5923 ,n5346 ,n5588);
    not g214(n3111 ,n3110);
    not g215(n3219 ,n3218);
    or g216(n5534 ,n5097 ,n5110);
    nor g217(n4138 ,n4015 ,n4022);
    xnor g218(n3399 ,n3332 ,n3358);
    nor g219(n2809 ,n2749 ,n2803);
    nor g220(n7312 ,n7280 ,n7311);
    nor g221(n4072 ,n4029 ,n4022);
    not g222(n5949 ,n5948);
    not g223(n7396 ,n7822);
    xor g224(n5795 ,n5310 ,n5414);
    not g225(n749 ,n1847);
    xnor g226(n602 ,n565 ,n510);
    nor g227(n4276 ,n4168 ,n4234);
    or g228(n1708 ,n1353 ,n1161);
    nor g229(n6569 ,n6382 ,n6458);
    nor g230(n4249 ,n4015 ,n4006);
    nor g231(n4346 ,n4047 ,n4195);
    nor g232(n4749 ,n4542 ,n4687);
    nor g233(n4962 ,n4863 ,n4930);
    xnor g234(n3435 ,n3360 ,n3251);
    not g235(n3113 ,n3112);
    nor g236(n4480 ,n4319 ,n4437);
    nor g237(n615 ,n593 ,n603);
    not g238(n5314 ,n5313);
    nor g239(n2626 ,n2562 ,n2613);
    nor g240(n7152 ,n7105 ,n7115);
    xnor g241(n6277 ,n5950 ,n6000);
    nor g242(n3980 ,n3937 ,n3979);
    not g243(n4047 ,n4046);
    not g244(n3382 ,n3381);
    xnor g245(n6979 ,n6862 ,n6910);
    nor g246(n6573 ,n6378 ,n6459);
    nor g247(n3052 ,n2994 ,n3038);
    or g248(n2574 ,n2438 ,n2516);
    nor g249(n2086 ,n2010 ,n2048);
    not g250(n2447 ,n21[5]);
    not g251(n7331 ,n41[15]);
    nor g252(n3645 ,n39[11] ,n7812);
    nor g253(n3085 ,n2995 ,n3029);
    dff g254(.RN(n1), .SN(1'b1), .CK(n0), .D(n1666), .Q(n35[3]));
    nor g255(n2905 ,n2782 ,n2889);
    nor g256(n4694 ,n4476 ,n4647);
    nor g257(n1402 ,n911 ,n642);
    or g258(n1768 ,n1406 ,n1548);
    nor g259(n7571 ,n7445 ,n7481);
    not g260(n4539 ,n4538);
    not g261(n975 ,n1835);
    not g262(n4529 ,n4528);
    xnor g263(n4817 ,n4743 ,n4630);
    xnor g264(n6715 ,n6545 ,n6589);
    xnor g265(n7821 ,n3787 ,n3807);
    nor g266(n3171 ,n2995 ,n3064);
    not g267(n2379 ,n2378);
    xnor g268(n2114 ,n1958 ,n2034);
    not g269(n7394 ,n7821);
    not g270(n3734 ,n3733);
    not g271(n830 ,n20[6]);
    xnor g272(n2316 ,n2286 ,n2263);
    xnor g273(n4676 ,n4534 ,n4532);
    nor g274(n7184 ,n7036 ,n7156);
    xnor g275(n1081 ,n814 ,n652);
    xnor g276(n6533 ,n6288 ,n5999);
    nor g277(n5186 ,n5108 ,n5099);
    not g278(n2221 ,n2220);
    nor g279(n4236 ,n4012 ,n4022);
    not g280(n858 ,n16[2]);
    xor g281(n1885 ,n1967 ,n2083);
    not g282(n7406 ,n7793);
    nor g283(n1545 ,n894 ,n641);
    nor g284(n3204 ,n3088 ,n3189);
    not g285(n6095 ,n6094);
    not g286(n1907 ,n19[3]);
    nor g287(n6772 ,n6651 ,n6649);
    nor g288(n6564 ,n6333 ,n6435);
    not g289(n3696 ,n3695);
    nor g290(n3914 ,n3899 ,n3913);
    nor g291(n2252 ,n2200 ,n2228);
    xnor g292(n6874 ,n6710 ,n6654);
    not g293(n5425 ,n5424);
    not g294(n2444 ,n7768);
    not g295(n3490 ,n3489);
    nor g296(n2535 ,n2433 ,n2519);
    nor g297(n4429 ,n4109 ,n4273);
    nor g298(n7671 ,n7471 ,n7487);
    nor g299(n3992 ,n3941 ,n3991);
    dff g300(.RN(n1), .SN(1'b1), .CK(n0), .D(n1668), .Q(n25[5]));
    nor g301(n6013 ,n5742 ,n5930);
    nor g302(n1177 ,n1106 ,n1068);
    nor g303(n5721 ,n5233 ,n5379);
    nor g304(n5732 ,n5167 ,n5229);
    nor g305(n1152 ,n1100 ,n1072);
    nor g306(n1489 ,n794 ,n639);
    not g307(n3319 ,n3318);
    nor g308(n3061 ,n3012 ,n3032);
    nor g309(n3089 ,n2995 ,n3030);
    or g310(n5521 ,n5091 ,n5109);
    xnor g311(n419 ,n331 ,n171);
    or g312(n2525 ,n2476 ,n2507);
    nor g313(n7608 ,n7401 ,n7476);
    not g314(n303 ,n302);
    nor g315(n5661 ,n5166 ,n5228);
    xnor g316(n2669 ,n2501 ,n2578);
    nor g317(n5646 ,n5124 ,n5474);
    xnor g318(n6413 ,n6243 ,n6038);
    not g319(n6329 ,n6328);
    not g320(n5325 ,n5324);
    nor g321(n3135 ,n3012 ,n3067);
    xnor g322(n7801 ,n1959 ,n1981);
    or g323(n1769 ,n1225 ,n1196);
    or g324(n1199 ,n1093 ,n1092);
    nor g325(n7586 ,n7452 ,n7477);
    not g326(n7353 ,n7810);
    xnor g327(n5818 ,n5284 ,n5508);
    nor g328(n4913 ,n4887 ,n4870);
    xnor g329(n2275 ,n2214 ,n2169);
    xor g330(n4393 ,n4269 ,n4084);
    nor g331(n2569 ,n2444 ,n2517);
    xnor g332(n6138 ,n5834 ,n5198);
    nor g333(n5028 ,n4962 ,n4998);
    xnor g334(n4779 ,n4674 ,n4518);
    nor g335(n6996 ,n6848 ,n6922);
    xnor g336(n6986 ,n6844 ,n6885);
    xnor g337(n7831 ,n3954 ,n3978);
    nor g338(n6475 ,n6194 ,n6350);
    nor g339(n4311 ,n4093 ,n4231);
    nor g340(n7467 ,n7393 ,n7396);
    nor g341(n6671 ,n6503 ,n6574);
    not g342(n2654 ,n2653);
    not g343(n254 ,n253);
    nor g344(n6365 ,n6094 ,n6246);
    not g345(n892 ,n33[5]);
    nor g346(n6334 ,n6015 ,n6207);
    not g347(n4521 ,n4520);
    nor g348(n6447 ,n6169 ,n6303);
    nor g349(n3939 ,n7779 ,n38[2]);
    nor g350(n6551 ,n6391 ,n6461);
    nor g351(n6485 ,n6203 ,n6325);
    not g352(n585 ,n584);
    nor g353(n516 ,n459 ,n490);
    xnor g354(n7070 ,n6878 ,n7021);
    not g355(n7445 ,n7799);
    nor g356(n2329 ,n2224 ,n2313);
    nor g357(n1429 ,n891 ,n640);
    nor g358(n3088 ,n2995 ,n3034);
    nor g359(n1470 ,n729 ,n639);
    xnor g360(n1850 ,n609 ,n612);
    xnor g361(n2279 ,n2160 ,n2239);
    not g362(n7447 ,n7791);
    nor g363(n1154 ,n1100 ,n1075);
    not g364(n6429 ,n6428);
    nor g365(n6887 ,n6839 ,n6773);
    not g366(n5963 ,n5962);
    nor g367(n3247 ,n3043 ,n3181);
    xnor g368(n552 ,n473 ,n505);
    xnor g369(n6243 ,n5815 ,n5550);
    or g370(n1011 ,n874 ,n931);
    nor g371(n6694 ,n6480 ,n6532);
    nor g372(n608 ,n577 ,n583);
    xnor g373(n4673 ,n4540 ,n4583);
    nor g374(n4127 ,n4018 ,n4024);
    nor g375(n4995 ,n4915 ,n4975);
    nor g376(n4824 ,n4690 ,n4799);
    nor g377(n1191 ,n1000 ,n1104);
    not g378(n794 ,n2[4]);
    nor g379(n6917 ,n6804 ,n6854);
    nor g380(n4648 ,n4500 ,n4520);
    xnor g381(n4767 ,n4591 ,n4682);
    nor g382(n4258 ,n4019 ,n4017);
    nor g383(n3589 ,n3559 ,n3588);
    dff g384(.RN(n1), .SN(1'b1), .CK(n0), .D(n1762), .Q(n28[13]));
    nor g385(n7589 ,n7374 ,n7476);
    nor g386(n5885 ,n5549 ,n5653);
    xnor g387(n4515 ,n4406 ,n4349);
    xnor g388(n2506 ,n2496 ,n2480);
    not g389(n4091 ,n4090);
    not g390(n4584 ,n4583);
    xor g391(n1874 ,n25[7] ,n120);
    nor g392(n6464 ,n6272 ,n6353);
    nor g393(n5238 ,n5112 ,n5089);
    nor g394(n1491 ,n790 ,n639);
    nor g395(n6006 ,n5737 ,n5903);
    not g396(n7371 ,n7725);
    or g397(n1615 ,n1272 ,n1483);
    xnor g398(n2145 ,n1971 ,n2093);
    not g399(n2108 ,n2107);
    nor g400(n2629 ,n2537 ,n2605);
    nor g401(n3661 ,n3591 ,n3616);
    nor g402(n6327 ,n6002 ,n6227);
    not g403(n6390 ,n6389);
    or g404(n1675 ,n1355 ,n1568);
    xnor g405(n3537 ,n3484 ,n3450);
    nor g406(n2422 ,n2372 ,n2421);
    nor g407(n2593 ,n2432 ,n2549);
    not g408(n2469 ,n2468);
    not g409(n3398 ,n3397);
    nor g410(n1268 ,n967 ,n638);
    nor g411(n5462 ,n5117 ,n5116);
    nor g412(n5602 ,n5484 ,n5182);
    nor g413(n5601 ,n5224 ,n5380);
    xor g414(n5790 ,n5521 ,n5254);
    nor g415(n6318 ,n6140 ,n6134);
    nor g416(n1442 ,n673 ,n634);
    or g417(n7640 ,n7548 ,n7576);
    nor g418(n5162 ,n5115 ,n5089);
    xor g419(n40[5] ,n39[6] ,n7834);
    or g420(n7651 ,n7569 ,n7568);
    xnor g421(n3433 ,n3331 ,n3364);
    xnor g422(n7758 ,n3999 ,n4005);
    xnor g423(n343 ,n241 ,n179);
    not g424(n4071 ,n4070);
    not g425(n938 ,n28[13]);
    or g426(n1637 ,n1305 ,n1572);
    xor g427(n4674 ,n4562 ,n4495);
    xnor g428(n4977 ,n4922 ,n4834);
    nor g429(n6226 ,n5965 ,n6025);
    nor g430(n5632 ,n5284 ,n5508);
    xnor g431(n3391 ,n3335 ,n3339);
    nor g432(n4100 ,n4020 ,n4026);
    xnor g433(n2712 ,n2515 ,n2641);
    not g434(n4010 ,n20[6]);
    nor g435(n3864 ,n3843 ,n3863);
    nor g436(n6571 ,n6384 ,n6416);
    not g437(n5219 ,n5218);
    not g438(n974 ,n1833);
    nor g439(n6699 ,n6473 ,n6522);
    nor g440(n5623 ,n5480 ,n5150);
    nor g441(n1535 ,n772 ,n641);
    nor g442(n2871 ,n2851 ,n2845);
    nor g443(n3652 ,n3597 ,n3594);
    or g444(n1582 ,n1243 ,n1469);
    nor g445(n3585 ,n3555 ,n3584);
    not g446(n5447 ,n5446);
    nor g447(n1252 ,n703 ,n640);
    xnor g448(n6630 ,n6399 ,n6180);
    nor g449(n1284 ,n975 ,n638);
    xnor g450(n7807 ,n2360 ,n2391);
    xnor g451(n7813 ,n2402 ,n2416);
    nor g452(n2935 ,n2900 ,n2906);
    nor g453(n389 ,n302 ,n345);
    nor g454(n5982 ,n5667 ,n5870);
    xnor g455(n6245 ,n5760 ,n5846);
    nor g456(n2564 ,n2433 ,n2517);
    nor g457(n6827 ,n6667 ,n6749);
    nor g458(n5266 ,n5115 ,n5111);
    xnor g459(n4552 ,n4378 ,n4267);
    nor g460(n4275 ,n4154 ,n4052);
    nor g461(n3810 ,n3780 ,n3809);
    nor g462(n1150 ,n1100 ,n1070);
    nor g463(n5647 ,n5430 ,n5372);
    or g464(n1729 ,n1368 ,n1173);
    not g465(n4683 ,n4682);
    nor g466(n2744 ,n2653 ,n2687);
    nor g467(n3946 ,n7787 ,n7772);
    nor g468(n3185 ,n3013 ,n3065);
    nor g469(n5126 ,n5096 ,n5119);
    nor g470(n1325 ,n959 ,n642);
    or g471(n5322 ,n5112 ,n5092);
    nor g472(n3257 ,n3082 ,n3187);
    nor g473(n4414 ,n4198 ,n4355);
    not g474(n3532 ,n3531);
    nor g475(n5717 ,n5457 ,n5417);
    xnor g476(n415 ,n343 ,n279);
    not g477(n3626 ,n7807);
    nor g478(n5460 ,n5099 ,n5097);
    xnor g479(n2735 ,n2672 ,n2625);
    xnor g480(n4867 ,n4771 ,n4723);
    not g481(n5255 ,n5254);
    xnor g482(n7140 ,n7101 ,n7060);
    nor g483(n1137 ,n641 ,n1048);
    nor g484(n4102 ,n4022 ,n4017);
    nor g485(n7306 ,n7274 ,n7293);
    nor g486(n1101 ,n18[2] ,n1018);
    xnor g487(n39[13] ,n2973 ,n2989);
    nor g488(n219 ,n146 ,n153);
    nor g489(n4838 ,n4763 ,n4797);
    xnor g490(n3959 ,n7791 ,n7776);
    nor g491(n4309 ,n4035 ,n4163);
    not g492(n4239 ,n4238);
    nor g493(n1543 ,n718 ,n641);
    not g494(n834 ,n22[5]);
    not g495(n6824 ,n6823);
    xnor g496(n2730 ,n2511 ,n2646);
    xor g497(n2423 ,n2458 ,n2470);
    xnor g498(n2959 ,n2933 ,n2926);
    xnor g499(n2214 ,n2139 ,n2154);
    nor g500(n5648 ,n5170 ,n5502);
    nor g501(n6484 ,n6206 ,n6321);
    nor g502(n3684 ,n3605 ,n3638);
    xor g503(n5830 ,n5309 ,n5152);
    nor g504(n3114 ,n3013 ,n3033);
    dff g505(.RN(n1), .SN(1'b1), .CK(n0), .D(n1616), .Q(n11[14]));
    nor g506(n7128 ,n7060 ,n7102);
    nor g507(n2768 ,n2668 ,n2726);
    nor g508(n137 ,n33[4] ,n135);
    or g509(n4137 ,n4006 ,n4009);
    not g510(n5121 ,n5120);
    xor g511(n5828 ,n5518 ,n5202);
    nor g512(n7568 ,n7385 ,n7476);
    not g513(n4169 ,n4168);
    xnor g514(n7757 ,n4000 ,n4003);
    xnor g515(n7814 ,n2395 ,n2418);
    xnor g516(n3397 ,n3333 ,n3228);
    not g517(n784 ,n4[6]);
    nor g518(n2847 ,n2675 ,n2816);
    xnor g519(n4873 ,n4770 ,n4717);
    dff g520(.RN(n1), .SN(1'b1), .CK(n0), .D(n1758), .Q(n22[7]));
    not g521(n7366 ,n7807);
    nor g522(n1262 ,n928 ,n640);
    nor g523(n6692 ,n6472 ,n6580);
    nor g524(n5262 ,n5096 ,n5089);
    not g525(n7395 ,n7817);
    not g526(n7336 ,n7824);
    nor g527(n5895 ,n5512 ,n5596);
    nor g528(n1504 ,n799 ,n639);
    nor g529(n5194 ,n5108 ,n5114);
    or g530(n7639 ,n7544 ,n7542);
    xnor g531(n4626 ,n4369 ,n4480);
    nor g532(n2256 ,n2159 ,n2239);
    not g533(n375 ,n374);
    xnor g534(n6612 ,n6415 ,n6168);
    dff g535(.RN(n1), .SN(1'b1), .CK(n0), .D(n1726), .Q(n31[2]));
    xnor g536(n6096 ,n5816 ,n5182);
    nor g537(n3780 ,n3698 ,n3745);
    nor g538(n6762 ,n6578 ,n6626);
    xnor g539(n7773 ,n3894 ,n3923);
    dff g540(.RN(n1), .SN(1'b1), .CK(n0), .D(n1671), .Q(n25[3]));
    not g541(n808 ,n18[0]);
    nor g542(n2980 ,n2939 ,n2979);
    not g543(n4736 ,n4735);
    xnor g544(n7171 ,n7108 ,n7087);
    xnor g545(n4955 ,n4900 ,n4908);
    not g546(n2369 ,n2368);
    xnor g547(n2299 ,n2129 ,n2252);
    nor g548(n1821 ,n1104 ,n1816);
    not g549(n5090 ,n21[0]);
    nor g550(n87 ,n85 ,n84);
    nor g551(n575 ,n536 ,n547);
    nor g552(n1207 ,n810 ,n1107);
    not g553(n2437 ,n21[6]);
    nor g554(n5886 ,n5329 ,n5632);
    not g555(n3869 ,n7805);
    not g556(n3207 ,n3206);
    nor g557(n4998 ,n4963 ,n4992);
    nor g558(n6753 ,n6589 ,n6698);
    nor g559(n2817 ,n2739 ,n2798);
    xnor g560(n3792 ,n3751 ,n3699);
    nor g561(n554 ,n500 ,n521);
    nor g562(n6304 ,n5997 ,n6220);
    not g563(n4358 ,n4357);
    xnor g564(n2885 ,n2812 ,n2839);
    nor g565(n6062 ,n5671 ,n5856);
    nor g566(n4295 ,n4060 ,n4224);
    not g567(n5959 ,n5958);
    not g568(n762 ,n4[3]);
    nor g569(n5408 ,n5115 ,n5099);
    not g570(n6093 ,n6092);
    nor g571(n1244 ,n935 ,n637);
    nor g572(n4994 ,n4934 ,n4988);
    nor g573(n300 ,n180 ,n242);
    not g574(n5098 ,n21[2]);
    nor g575(n57 ,n46 ,n47);
    nor g576(n6379 ,n6155 ,n6153);
    xnor g577(n2781 ,n2709 ,n2426);
    nor g578(n1317 ,n914 ,n642);
    not g579(n967 ,n19[1]);
    not g580(n5331 ,n5330);
    nor g581(n2552 ,n2445 ,n2525);
    nor g582(n2761 ,n2721 ,n2695);
    nor g583(n2613 ,n2444 ,n2548);
    xnor g584(n4716 ,n4548 ,n4628);
    nor g585(n2289 ,n2231 ,n2259);
    nor g586(n3521 ,n3471 ,n3487);
    not g587(n2865 ,n2864);
    or g588(n7707 ,n7616 ,n7680);
    xnor g589(n5061 ,n5019 ,n5033);
    xnor g590(n2683 ,n2515 ,n2599);
    not g591(n6047 ,n6046);
    not g592(n218 ,n217);
    dff g593(.RN(n1), .SN(1'b1), .CK(n0), .D(n1599), .Q(n19[3]));
    nor g594(n5414 ,n5089 ,n5091);
    not g595(n2288 ,n2287);
    nor g596(n7241 ,n7219 ,n7211);
    xnor g597(n6080 ,n5823 ,n5304);
    nor g598(n5188 ,n5103 ,n5109);
    nor g599(n1434 ,n883 ,n1103);
    nor g600(n5637 ,n5374 ,n5126);
    xnor g601(n3333 ,n3106 ,n3257);
    not g602(n5185 ,n5184);
    or g603(n1718 ,n1228 ,n1538);
    nor g604(n3979 ,n3954 ,n3978);
    nor g605(n1559 ,n913 ,n1106);
    not g606(n3723 ,n3722);
    not g607(n636 ,n634);
    not g608(n4105 ,n4104);
    not g609(n4153 ,n4152);
    or g610(n1698 ,n1309 ,n1530);
    dff g611(.RN(n1), .SN(1'b1), .CK(n0), .D(n1712), .Q(n32[2]));
    nor g612(n6757 ,n6478 ,n6630);
    dff g613(.RN(n1), .SN(1'b1), .CK(n0), .D(n1761), .Q(n22[5]));
    or g614(n5303 ,n5100 ,n5105);
    nor g615(n1526 ,n727 ,n641);
    not g616(n6480 ,n6479);
    not g617(n6929 ,n6928);
    dff g618(.RN(n1), .SN(1'b1), .CK(n0), .D(n1626), .Q(n11[8]));
    not g619(n4262 ,n4261);
    not g620(n924 ,n33[1]);
    nor g621(n2504 ,n2468 ,n2490);
    xnor g622(n7262 ,n7216 ,n7235);
    xnor g623(n2971 ,n2948 ,n2920);
    nor g624(n4624 ,n4489 ,n4572);
    xnor g625(n3320 ,n3110 ,n3210);
    or g626(n3035 ,n2996 ,n2999);
    nor g627(n5913 ,n5307 ,n5641);
    nor g628(n6724 ,n6439 ,n6687);
    dff g629(.RN(n1), .SN(1'b1), .CK(n0), .D(n1617), .Q(n11[13]));
    nor g630(n1519 ,n745 ,n641);
    or g631(n1747 ,n1387 ,n1170);
    not g632(n6516 ,n6515);
    nor g633(n2866 ,n2818 ,n2848);
    nor g634(n2798 ,n2734 ,n2760);
    not g635(n907 ,n28[9]);
    or g636(n7701 ,n7673 ,n7655);
    xnor g637(n2085 ,n1969 ,n1984);
    nor g638(n6307 ,n6261 ,n6132);
    nor g639(n1473 ,n751 ,n639);
    nor g640(n357 ,n266 ,n291);
    nor g641(n5728 ,n5195 ,n5241);
    not g642(n5020 ,n5019);
    or g643(n7675 ,n7503 ,n7667);
    xnor g644(n39[8] ,n2942 ,n2979);
    not g645(n5106 ,n19[3]);
    not g646(n951 ,n12[14]);
    xnor g647(n3793 ,n3725 ,n3710);
    nor g648(n1107 ,n18[0] ,n1016);
    nor g649(n2095 ,n1999 ,n2045);
    not g650(n7199 ,n7198);
    not g651(n6617 ,n6616);
    xor g652(n5773 ,n5323 ,n5184);
    not g653(n7086 ,n7085);
    not g654(n3612 ,n7789);
    nor g655(n1872 ,n131 ,n132);
    nor g656(n4220 ,n4011 ,n4006);
    not g657(n3159 ,n3158);
    nor g658(n2855 ,n2793 ,n2822);
    xnor g659(n3751 ,n39[12] ,n3676);
    nor g660(n1296 ,n915 ,n637);
    xnor g661(n1036 ,n881 ,n840);
    not g662(n6433 ,n6432);
    not g663(n44 ,n37[5]);
    not g664(n2705 ,n2704);
    not g665(n721 ,n12[4]);
    xor g666(n340 ,n198 ,n245);
    nor g667(n4437 ,n4239 ,n4282);
    nor g668(n2981 ,n2980 ,n2937);
    nor g669(n7027 ,n7000 ,n7009);
    nor g670(n6439 ,n6201 ,n6337);
    not g671(n6544 ,n6543);
    nor g672(n3279 ,n3208 ,n3200);
    dff g673(.RN(n1), .SN(1'b1), .CK(n0), .D(n1594), .Q(n19[5]));
    nor g674(n1501 ,n737 ,n1099);
    nor g675(n1868 ,n143 ,n144);
    nor g676(n2738 ,n2715 ,n2710);
    xnor g677(n3782 ,n3733 ,n3695);
    nor g678(n4450 ,n4199 ,n4356);
    nor g679(n1332 ,n855 ,n637);
    nor g680(n4487 ,n4350 ,n4406);
    nor g681(n3926 ,n3891 ,n3925);
    xnor g682(n3729 ,n39[14] ,n3670);
    nor g683(n5675 ,n5375 ,n5127);
    or g684(n7481 ,n7326 ,n7325);
    nor g685(n5920 ,n5345 ,n5636);
    nor g686(n537 ,n410 ,n506);
    nor g687(n3885 ,n7801 ,n7793);
    not g688(n5115 ,n22[0]);
    nor g689(n4894 ,n4865 ,n4867);
    not g690(n3024 ,n7752);
    xnor g691(n4714 ,n4550 ,n4624);
    not g692(n4113 ,n4112);
    xnor g693(n7843 ,n3900 ,n3905);
    not g694(n5487 ,n5486);
    nor g695(n4125 ,n4021 ,n4017);
    nor g696(n4172 ,n4011 ,n4018);
    not g697(n194 ,n193);
    not g698(n739 ,n4[2]);
    xnor g699(n6737 ,n6491 ,n6418);
    xnor g700(n5821 ,n5144 ,n5438);
    not g701(n2693 ,n2692);
    nor g702(n6222 ,n6021 ,n5971);
    nor g703(n3523 ,n3476 ,n3494);
    nor g704(n2795 ,n2729 ,n2753);
    nor g705(n1560 ,n962 ,n1106);
    nor g706(n3087 ,n2995 ,n3041);
    not g707(n4097 ,n4096);
    nor g708(n1418 ,n901 ,n637);
    nor g709(n593 ,n555 ,n573);
    nor g710(n3777 ,n3722 ,n3738);
    buf g711(n37[6] ,n1837);
    nor g712(n7657 ,n7472 ,n7488);
    nor g713(n3757 ,n3695 ,n3734);
    nor g714(n2127 ,n1970 ,n2085);
    xnor g715(n6796 ,n6597 ,n6533);
    nor g716(n2120 ,n1970 ,n2099);
    nor g717(n2356 ,n2310 ,n2330);
    nor g718(n2579 ,n2487 ,n2563);
    nor g719(n6587 ,n6381 ,n6456);
    or g720(n1010 ,n878 ,n960);
    nor g721(n2793 ,n2651 ,n2748);
    nor g722(n2374 ,n2346 ,n2344);
    xnor g723(n6913 ,n6792 ,n6833);
    not g724(n5253 ,n5252);
    xnor g725(n1854 ,n475 ,n457);
    not g726(n2112 ,n2111);
    nor g727(n7251 ,n7233 ,n7209);
    not g728(n6619 ,n6618);
    nor g729(n3982 ,n3940 ,n3981);
    xnor g730(n3073 ,n40[7] ,n7746);
    nor g731(n6044 ,n5724 ,n5904);
    xor g732(n6167 ,n5774 ,n5563);
    nor g733(n7577 ,n7357 ,n7480);
    xnor g734(n2713 ,n2513 ,n2630);
    nor g735(n2762 ,n2708 ,n2702);
    nor g736(n536 ,n449 ,n503);
    nor g737(n7493 ,n7352 ,n7475);
    nor g738(n2202 ,n2105 ,n2165);
    xnor g739(n2272 ,n2212 ,n2098);
    xnor g740(n2129 ,n1959 ,n2100);
    xnor g741(n1023 ,n36[9] ,n34[9]);
    xnor g742(n2690 ,n2514 ,n2647);
    not g743(n6172 ,n6171);
    nor g744(n4701 ,n4549 ,n4628);
    not g745(n6869 ,n6868);
    not g746(n529 ,n528);
    nor g747(n1520 ,n796 ,n641);
    nor g748(n4277 ,n4222 ,n4058);
    nor g749(n4222 ,n4023 ,n4022);
    nor g750(n1949 ,n1920 ,n1934);
    nor g751(n5668 ,n5279 ,n5165);
    nor g752(n1373 ,n831 ,n1103);
    nor g753(n1259 ,n910 ,n640);
    nor g754(n3778 ,n3700 ,n3751);
    nor g755(n1565 ,n683 ,n635);
    xnor g756(n4363 ,n4182 ,n4210);
    not g757(n6149 ,n6148);
    nor g758(n1960 ,n1939 ,n1948);
    nor g759(n2280 ,n2244 ,n2255);
    not g760(n4937 ,n4936);
    nor g761(n4440 ,n4120 ,n4286);
    nor g762(n6032 ,n5720 ,n5894);
    not g763(n953 ,n28[14]);
    xnor g764(n4671 ,n4546 ,n4587);
    nor g765(n6539 ,n6371 ,n6447);
    not g766(n5393 ,n5392);
    not g767(n6087 ,n6086);
    nor g768(n2961 ,n2930 ,n2946);
    nor g769(n2916 ,n2826 ,n2887);
    not g770(n4065 ,n4064);
    not g771(n870 ,n28[4]);
    nor g772(n1469 ,n739 ,n639);
    nor g773(n1950 ,n1922 ,n1941);
    xnor g774(n6293 ,n5968 ,n5952);
    not g775(n1897 ,n19[4]);
    nor g776(n1513 ,n784 ,n639);
    nor g777(n1112 ,n635 ,n1022);
    or g778(n7642 ,n7552 ,n7549);
    xnor g779(n355 ,n255 ,n193);
    nor g780(n6816 ,n6618 ,n6737);
    nor g781(n2591 ,n2434 ,n2548);
    not g782(n7334 ,n7820);
    nor g783(n5192 ,n5095 ,n5111);
    nor g784(n3296 ,n3149 ,n3206);
    nor g785(n6055 ,n5669 ,n5882);
    nor g786(n6910 ,n6768 ,n6815);
    nor g787(n5639 ,n5408 ,n5282);
    nor g788(n6560 ,n6241 ,n6427);
    not g789(n2802 ,n2801);
    nor g790(n6362 ,n6239 ,n6121);
    xnor g791(n6872 ,n6711 ,n6519);
    not g792(n3238 ,n3237);
    nor g793(n5952 ,n5699 ,n5862);
    xnor g794(n7777 ,n3887 ,n3931);
    xnor g795(n3951 ,n7792 ,n7777);
    nor g796(n289 ,n221 ,n229);
    not g797(n4974 ,n4973);
    xnor g798(n1032 ,n859 ,n849);
    not g799(n5580 ,n5579);
    not g800(n4250 ,n4249);
    nor g801(n1293 ,n906 ,n636);
    not g802(n4271 ,n4270);
    not g803(n3512 ,n3511);
    dff g804(.RN(n1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n20[2]));
    nor g805(n6199 ,n5972 ,n5938);
    dff g806(.RN(n1), .SN(1'b1), .CK(n0), .D(n1716), .Q(n32[0]));
    nor g807(n2536 ,n2434 ,n2523);
    not g808(n646 ,n24[4]);
    nor g809(n4571 ,n4456 ,n4464);
    xnor g810(n4524 ,n4383 ,n4141);
    xnor g811(n5787 ,n5418 ,n5258);
    xnor g812(n3677 ,n7807 ,n7784);
    not g813(n43 ,n37[4]);
    nor g814(n1921 ,n1900 ,n1899);
    not g815(n6077 ,n6076);
    xnor g816(n6884 ,n6714 ,n6483);
    nor g817(n7131 ,n6971 ,n7080);
    dff g818(.RN(n1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n22[2]));
    not g819(n3700 ,n3699);
    nor g820(n7049 ,n6937 ,n6993);
    xnor g821(n3064 ,n40[5] ,n7744);
    xnor g822(n2522 ,n2424 ,n2505);
    nor g823(n1457 ,n733 ,n634);
    xnor g824(n7236 ,n7198 ,n7147);
    or g825(n1684 ,n1335 ,n1526);
    xor g826(n5804 ,n5321 ,n5252);
    xor g827(n7744 ,n7806 ,n7783);
    nor g828(n3685 ,n3611 ,n3640);
    nor g829(n2010 ,n1890 ,n1974);
    nor g830(n175 ,n154 ,n157);
    nor g831(n1919 ,n1908 ,n1905);
    nor g832(n2453 ,n21[5] ,n22[5]);
    xor g833(n6411 ,n6175 ,n6074);
    xor g834(n7743 ,n7805 ,n7782);
    not g835(n6803 ,n6802);
    xnor g836(n2218 ,n2112 ,n2172);
    nor g837(n5898 ,n5343 ,n5659);
    nor g838(n3937 ,n7785 ,n7770);
    dff g839(.RN(n1), .SN(1'b1), .CK(n0), .D(n1659), .Q(n35[6]));
    dff g840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1635), .Q(n11[0]));
    or g841(n7665 ,n7601 ,n7599);
    nor g842(n4443 ,n4142 ,n4287);
    xnor g843(n7287 ,n7260 ,n7251);
    nor g844(n4056 ,n4029 ,n4018);
    nor g845(n213 ,n150 ,n149);
    nor g846(n4636 ,n4309 ,n4576);
    xnor g847(n3568 ,n3539 ,n3523);
    nor g848(n1475 ,n767 ,n639);
    not g849(n1104 ,n1105);
    nor g850(n3759 ,n3699 ,n3752);
    not g851(n115 ,n114);
    nor g852(n2597 ,n2443 ,n2548);
    nor g853(n1264 ,n712 ,n640);
    nor g854(n1811 ,n1106 ,n1809);
    not g855(n7450 ,n7771);
    xnor g856(n2711 ,n2513 ,n2626);
    xnor g857(n3552 ,n3509 ,n3501);
    xnor g858(n346 ,n207 ,n209);
    dff g859(.RN(n1), .SN(1'b1), .CK(n0), .D(n1706), .Q(n32[5]));
    xnor g860(n4930 ,n4860 ,n4830);
    xnor g861(n5770 ,n5406 ,n5386);
    nor g862(n1201 ,n811 ,n1107);
    nor g863(n6237 ,n6031 ,n6035);
    nor g864(n3488 ,n3417 ,n3461);
    nor g865(n5936 ,n5681 ,n5876);
    xnor g866(n580 ,n546 ,n543);
    not g867(n5217 ,n5216);
    nor g868(n6839 ,n6697 ,n6748);
    xnor g869(n4608 ,n4501 ,n4460);
    nor g870(n2993 ,n2951 ,n2992);
    nor g871(n5665 ,n5369 ,n5221);
    nor g872(n3167 ,n3012 ,n3063);
    xnor g873(n39[7] ,n2941 ,n2975);
    xnor g874(n6106 ,n5768 ,n5142);
    xor g875(n7841 ,n3898 ,n3910);
    xnor g876(n6086 ,n5780 ,n5398);
    not g877(n3621 ,n7785);
    nor g878(n6038 ,n5719 ,n5915);
    nor g879(n1117 ,n634 ,n1051);
    nor g880(n512 ,n465 ,n498);
    nor g881(n4968 ,n4882 ,n4929);
    nor g882(n5940 ,n5662 ,n5889);
    xnor g883(n6140 ,n5830 ,n5486);
    nor g884(n1386 ,n960 ,n1101);
    nor g885(n5998 ,n5726 ,n5917);
    xor g886(n1889 ,n2127 ,n2116);
    nor g887(n444 ,n304 ,n400);
    xor g888(n6166 ,n5794 ,n5212);
    not g889(n4246 ,n4245);
    nor g890(n3475 ,n3386 ,n3424);
    xnor g891(n7845 ,n3893 ,n3886);
    nor g892(n5722 ,n5471 ,n5397);
    nor g893(n2236 ,n2169 ,n2203);
    nor g894(n3189 ,n3013 ,n3066);
    dff g895(.RN(n1), .SN(1'b1), .CK(n0), .D(n1641), .Q(n10[10]));
    not g896(n539 ,n538);
    nor g897(n5396 ,n5115 ,n5105);
    xnor g898(n3414 ,n3341 ,n3230);
    not g899(n5102 ,n37[6]);
    nor g900(n5504 ,n5098 ,n5104);
    nor g901(n1134 ,n641 ,n1027);
    or g902(n1665 ,n1385 ,n1520);
    or g903(n7680 ,n7605 ,n7657);
    nor g904(n2396 ,n2362 ,n2383);
    not g905(n3611 ,n7787);
    nor g906(n3057 ,n3012 ,n3038);
    nor g907(n3968 ,n3936 ,n3967);
    not g908(n846 ,n34[5]);
    not g909(n2106 ,n2105);
    not g910(n4221 ,n4220);
    nor g911(n3460 ,n3383 ,n3427);
    nor g912(n3190 ,n3013 ,n3067);
    not g913(n4625 ,n4624);
    or g914(n7613 ,n7497 ,n7529);
    dff g915(.RN(n1), .SN(1'b1), .CK(n0), .D(n1622), .Q(n11[10]));
    not g916(n5973 ,n5972);
    not g917(n4185 ,n4184);
    buf g918(n14[13], n11[13]);
    nor g919(n4654 ,n4503 ,n4537);
    nor g920(n3353 ,n3222 ,n3286);
    xnor g921(n413 ,n342 ,n211);
    nor g922(n1356 ,n848 ,n636);
    nor g923(n373 ,n284 ,n352);
    nor g924(n5418 ,n5090 ,n5111);
    nor g925(n6733 ,n6636 ,n6634);
    nor g926(n4705 ,n4551 ,n4624);
    nor g927(n5918 ,n5344 ,n5637);
    or g928(n1801 ,n1438 ,n1515);
    nor g929(n7091 ,n7043 ,n7053);
    nor g930(n4048 ,n4014 ,n4020);
    nor g931(n4695 ,n4474 ,n4648);
    nor g932(n6802 ,n6607 ,n6755);
    nor g933(n5699 ,n5239 ,n5405);
    nor g934(n2599 ,n2445 ,n2549);
    xnor g935(n4769 ,n4626 ,n4709);
    nor g936(n2609 ,n2434 ,n2574);
    nor g937(n1395 ,n664 ,n640);
    not g938(n642 ,n641);
    nor g939(n1856 ,n285 ,n328);
    nor g940(n5736 ,n5163 ,n5267);
    nor g941(n5378 ,n5117 ,n5098);
    nor g942(n4476 ,n4346 ,n4436);
    nor g943(n7045 ,n6949 ,n6987);
    nor g944(n7322 ,n7272 ,n7321);
    not g945(n4742 ,n4741);
    xnor g946(n399 ,n333 ,n352);
    not g947(n3620 ,n39[8]);
    or g948(n3029 ,n3016 ,n3009);
    nor g949(n4882 ,n4806 ,n4840);
    nor g950(n4353 ,n4149 ,n4250);
    not g951(n3025 ,n7749);
    nor g952(n2796 ,n2426 ,n2759);
    xnor g953(n1082 ,n812 ,n651);
    xnor g954(n7159 ,n7088 ,n7043);
    nor g955(n1116 ,n634 ,n1050);
    nor g956(n4808 ,n4527 ,n4740);
    nor g957(n7234 ,n7206 ,n7188);
    nor g958(n6455 ,n6164 ,n6316);
    not g959(n305 ,n304);
    not g960(n5193 ,n5192);
    nor g961(n5258 ,n5112 ,n5114);
    nor g962(n3908 ,n3884 ,n3907);
    xnor g963(n6394 ,n6146 ,n6144);
    nor g964(n3588 ,n3562 ,n3587);
    nor g965(n2193 ,n2111 ,n2135);
    not g966(n2689 ,n2688);
    xnor g967(n2169 ,n1968 ,n2068);
    xnor g968(n6878 ,n6713 ,n6493);
    not g969(n5536 ,n5535);
    not g970(n890 ,n31[7]);
    buf g971(n37[0] ,n1831);
    or g972(n1581 ,n1242 ,n1109);
    nor g973(n5226 ,n5093 ,n5105);
    dff g974(.RN(n1), .SN(1'b1), .CK(n0), .D(n1577), .Q(n12[15]));
    or g975(n1767 ,n1407 ,n1498);
    xnor g976(n2366 ,n2315 ,n2299);
    nor g977(n3930 ,n3892 ,n3929);
    nor g978(n3995 ,n37[2] ,n20[2]);
    dff g979(.RN(n1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n21[5]));
    nor g980(n253 ,n150 ,n155);
    nor g981(n4842 ,n4761 ,n4783);
    nor g982(n7280 ,n7259 ,n7241);
    nor g983(n2567 ,n2444 ,n2521);
    xnor g984(n6713 ,n6507 ,n6550);
    nor g985(n1554 ,n714 ,n1100);
    xnor g986(n4411 ,n4038 ,n4178);
    xnor g987(n4739 ,n4612 ,n4482);
    xnor g988(n3550 ,n3507 ,n3499);
    nor g989(n2090 ,n1991 ,n2066);
    nor g990(n2985 ,n2965 ,n2984);
    not g991(n649 ,n35[1]);
    nor g992(n1404 ,n714 ,n642);
    not g993(n5097 ,n21[4]);
    xnor g994(n2364 ,n2318 ,n2289);
    nor g995(n2587 ,n2434 ,n2547);
    dff g996(.RN(n1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n28[3]));
    not g997(n148 ,n19[6]);
    nor g998(n3803 ,n3753 ,n3802);
    nor g999(n6957 ,n6789 ,n6880);
    nor g1000(n6063 ,n5735 ,n5909);
    nor g1001(n2405 ,n2379 ,n2392);
    nor g1002(n3131 ,n3012 ,n3070);
    nor g1003(n6215 ,n5753 ,n6037);
    xnor g1004(n4544 ,n4391 ,n4104);
    or g1005(n7677 ,n7574 ,n7669);
    nor g1006(n2627 ,n2529 ,n2595);
    nor g1007(n628 ,n604 ,n627);
    nor g1008(n3297 ,n3154 ,n3260);
    nor g1009(n6588 ,n6360 ,n6463);
    not g1010(n4724 ,n4723);
    not g1011(n2223 ,n2222);
    nor g1012(n7157 ,n7052 ,n7124);
    xnor g1013(n7786 ,n5061 ,n5073);
    nor g1014(n5633 ,n5180 ,n5428);
    nor g1015(n5588 ,n5358 ,n5248);
    dff g1016(.RN(n1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n16[6]));
    nor g1017(n2912 ,n2874 ,n2886);
    nor g1018(n5899 ,n5531 ,n5654);
    dff g1019(.RN(n1), .SN(1'b1), .CK(n0), .D(n1730), .Q(n31[0]));
    nor g1020(n3494 ,n3416 ,n3468);
    nor g1021(n317 ,n222 ,n230);
    nor g1022(n1364 ,n666 ,n1105);
    not g1023(n6873 ,n6872);
    not g1024(n7434 ,n39[1]);
    not g1025(n2262 ,n2261);
    xnor g1026(n6706 ,n6503 ,n6588);
    not g1027(n837 ,n34[0]);
    not g1028(n3248 ,n3247);
    nor g1029(n3169 ,n2995 ,n3075);
    xor g1030(n7748 ,n7810 ,n7787);
    nor g1031(n3227 ,n3091 ,n3171);
    nor g1032(n1365 ,n689 ,n1103);
    nor g1033(n5684 ,n5153 ,n5487);
    xnor g1034(n6301 ,n5942 ,n6040);
    or g1035(n1600 ,n1266 ,n1480);
    nor g1036(n1474 ,n746 ,n639);
    not g1037(n4237 ,n4236);
    nor g1038(n3374 ,n3305 ,n3347);
    xnor g1039(n7278 ,n7236 ,n7253);
    nor g1040(n4418 ,n4260 ,n4272);
    nor g1041(n3045 ,n2994 ,n3039);
    nor g1042(n5128 ,n5091 ,n5106);
    xnor g1043(n5781 ,n5380 ,n5224);
    nor g1044(n7595 ,n7342 ,n7481);
    nor g1045(n3754 ,n3697 ,n3746);
    nor g1046(n2592 ,n2442 ,n2549);
    nor g1047(n1357 ,n667 ,n637);
    xor g1048(n1883 ,n1910 ,n1931);
    not g1049(n45 ,n37[2]);
    nor g1050(n2243 ,n2079 ,n2208);
    dff g1051(.RN(n1), .SN(1'b1), .CK(n0), .D(n1665), .Q(n25[6]));
    nor g1052(n7541 ,n7376 ,n7478);
    xor g1053(n5807 ,n5561 ,n5478);
    nor g1054(n6375 ,n6137 ,n6123);
    nor g1055(n358 ,n272 ,n301);
    nor g1056(n4308 ,n4206 ,n4204);
    xnor g1057(n3847 ,n37[5] ,n19[5]);
    nor g1058(n7296 ,n7263 ,n7286);
    nor g1059(n3251 ,n3053 ,n3132);
    nor g1060(n3406 ,n3311 ,n3363);
    xnor g1061(n6876 ,n6719 ,n6584);
    not g1062(n5991 ,n5990);
    nor g1063(n2186 ,n1959 ,n2159);
    nor g1064(n7015 ,n6897 ,n6945);
    not g1065(n925 ,n12[10]);
    or g1066(n1777 ,n1414 ,n1502);
    nor g1067(n393 ,n300 ,n367);
    nor g1068(n6326 ,n6061 ,n6215);
    nor g1069(n1934 ,n1906 ,n1915);
    nor g1070(n4965 ,n4911 ,n4937);
    xnor g1071(n6781 ,n6614 ,n6575);
    nor g1072(n2571 ,n2445 ,n2523);
    nor g1073(n1412 ,n872 ,n642);
    or g1074(n7636 ,n7546 ,n7539);
    nor g1075(n2940 ,n2786 ,n2910);
    not g1076(n694 ,n1838);
    nor g1077(n5706 ,n5395 ,n5231);
    xnor g1078(n7036 ,n6914 ,n6880);
    xnor g1079(n4686 ,n4517 ,n4355);
    xnor g1080(n6402 ,n6255 ,n6251);
    nor g1081(n2281 ,n2253 ,n2256);
    not g1082(n7407 ,n7732);
    nor g1083(n5726 ,n5255 ,n5287);
    nor g1084(n4848 ,n4729 ,n4782);
    not g1085(n7016 ,n7015);
    nor g1086(n2915 ,n2854 ,n2895);
    not g1087(n456 ,n455);
    nor g1088(n2741 ,n2705 ,n2688);
    nor g1089(n7097 ,n7012 ,n7059);
    not g1090(n811 ,n27[3]);
    nor g1091(n3281 ,n3160 ,n3246);
    not g1092(n6875 ,n6874);
    or g1093(n1681 ,n1324 ,n1524);
    buf g1094(n37[1] ,n1832);
    nor g1095(n3349 ,n3229 ,n3271);
    nor g1096(n5046 ,n4986 ,n5022);
    not g1097(n3633 ,n39[5]);
    xnor g1098(n4546 ,n4372 ,n4160);
    not g1099(n3593 ,n7779);
    not g1100(n2377 ,n2376);
    xnor g1101(n3667 ,n7812 ,n7789);
    nor g1102(n1477 ,n754 ,n639);
    or g1103(n7682 ,n7611 ,n7665);
    xnor g1104(n429 ,n334 ,n247);
    nor g1105(n297 ,n161 ,n195);
    or g1106(n1611 ,n1275 ,n1120);
    xnor g1107(n4971 ,n4940 ,n4614);
    nor g1108(n4118 ,n4015 ,n4021);
    xnor g1109(n6298 ,n5976 ,n6050);
    nor g1110(n7566 ,n7348 ,n7477);
    nor g1111(n6947 ,n6704 ,n6901);
    not g1112(n5235 ,n5234);
    not g1113(n4543 ,n4542);
    nor g1114(n5122 ,n5101 ,n5114);
    nor g1115(n4580 ,n4176 ,n4471);
    or g1116(n7617 ,n7505 ,n7504);
    not g1117(n2709 ,n2708);
    nor g1118(n4040 ,n4012 ,n4021);
    nor g1119(n2630 ,n2568 ,n2588);
    nor g1120(n5476 ,n5112 ,n5102);
    xnor g1121(n6142 ,n5805 ,n5466);
    xnor g1122(n1028 ,n678 ,n672);
    or g1123(n1799 ,n1206 ,n1341);
    not g1124(n4163 ,n4162);
    xnor g1125(n6777 ,n6624 ,n6704);
    nor g1126(n1463 ,n1839 ,n634);
    nor g1127(n3542 ,n3480 ,n3513);
    not g1128(n6266 ,n6265);
    xnor g1129(n2904 ,n2864 ,n2841);
    nor g1130(n1476 ,n750 ,n639);
    nor g1131(n4283 ,n4036 ,n4156);
    not g1132(n5419 ,n5418);
    not g1133(n1900 ,n19[0]);
    nor g1134(n6364 ,n6088 ,n6085);
    nor g1135(n542 ,n469 ,n515);
    nor g1136(n1465 ,n847 ,n635);
    or g1137(n5562 ,n5089 ,n5116);
    nor g1138(n4337 ,n4233 ,n4033);
    nor g1139(n5652 ,n5450 ,n5270);
    nor g1140(n6948 ,n6763 ,n6884);
    not g1141(n950 ,n10[15]);
    nor g1142(n3804 ,n3768 ,n3803);
    nor g1143(n2034 ,n1957 ,n2016);
    not g1144(n840 ,n22[3]);
    nor g1145(n6219 ,n5743 ,n5957);
    dff g1146(.RN(n1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n17[3]));
    xnor g1147(n6914 ,n6788 ,n6842);
    nor g1148(n5364 ,n5095 ,n5109);
    xnor g1149(n7823 ,n3785 ,n3803);
    not g1150(n136 ,n135);
    nor g1151(n5649 ,n5262 ,n5364);
    xnor g1152(n6982 ,n6852 ,n6811);
    not g1153(n7351 ,n40[3]);
    xor g1154(n5789 ,n5569 ,n5204);
    not g1155(n700 ,n25[6]);
    not g1156(n3994 ,n37[0]);
    nor g1157(n294 ,n235 ,n175);
    or g1158(n1824 ,n1132 ,n1821);
    not g1159(n7348 ,n7814);
    nor g1160(n6273 ,n5929 ,n5933);
    or g1161(n7478 ,n7326 ,n7324);
    xnor g1162(n6415 ,n6247 ,n6080);
    nor g1163(n3362 ,n3282 ,n3354);
    dff g1164(.RN(n1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n21[0]));
    nor g1165(n2255 ,n2242 ,n2189);
    nor g1166(n2457 ,n21[0] ,n22[0]);
    nor g1167(n2868 ,n2676 ,n2847);
    xnor g1168(n2881 ,n2837 ,n2817);
    not g1169(n6534 ,n6533);
    nor g1170(n5701 ,n5145 ,n5439);
    nor g1171(n2540 ,n2442 ,n2521);
    nor g1172(n6059 ,n5709 ,n5896);
    xnor g1173(n3395 ,n3330 ,n3229);
    xor g1174(n442 ,n321 ,n380);
    not g1175(n517 ,n516);
    nor g1176(n4216 ,n4018 ,n4026);
    nor g1177(n2123 ,n1972 ,n2082);
    not g1178(n687 ,n36[14]);
    nor g1179(n3545 ,n3500 ,n3508);
    xnor g1180(n7817 ,n3781 ,n3823);
    nor g1181(n6891 ,n6616 ,n6787);
    not g1182(n4633 ,n4632);
    buf g1183(n13[8], n10[8]);
    nor g1184(n1161 ,n1102 ,n1064);
    or g1185(n1775 ,n1412 ,n1137);
    nor g1186(n5702 ,n5415 ,n5131);
    or g1187(n1604 ,n1265 ,n1131);
    or g1188(n1654 ,n1436 ,n1554);
    nor g1189(n1278 ,n936 ,n638);
    nor g1190(n7190 ,n7041 ,n7143);
    xnor g1191(n5849 ,n5565 ,n5188);
    nor g1192(n3099 ,n3012 ,n3042);
    nor g1193(n2541 ,n2432 ,n2519);
    not g1194(n6657 ,n6656);
    not g1195(n6621 ,n6620);
    not g1196(n755 ,n4[5]);
    not g1197(n125 ,n33[1]);
    nor g1198(n5218 ,n5097 ,n5105);
    nor g1199(n5390 ,n5093 ,n5104);
    nor g1200(n2342 ,n2254 ,n2332);
    or g1201(n7622 ,n7517 ,n7516);
    nor g1202(n2094 ,n2023 ,n2052);
    nor g1203(n5888 ,n5294 ,n5639);
    not g1204(n791 ,n8[0]);
    xnor g1205(n6287 ,n5753 ,n6036);
    nor g1206(n3763 ,n3711 ,n3725);
    nor g1207(n6337 ,n6057 ,n6238);
    not g1208(n918 ,n19[5]);
    not g1209(n1958 ,n1959);
    not g1210(n4590 ,n4589);
    nor g1211(n5301 ,n5089 ,n5090);
    nor g1212(n3753 ,n3701 ,n3736);
    nor g1213(n4823 ,n4636 ,n4796);
    nor g1214(n7005 ,n6868 ,n6938);
    not g1215(n4519 ,n4518);
    nor g1216(n5404 ,n5098 ,n5111);
    not g1217(n5031 ,n5030);
    xnor g1218(n1062 ,n36[15] ,n34[15]);
    xnor g1219(n6503 ,n6284 ,n5980);
    not g1220(n7148 ,n7147);
    not g1221(n6576 ,n6575);
    nor g1222(n2565 ,n2431 ,n2517);
    nor g1223(n1528 ,n761 ,n641);
    nor g1224(n1114 ,n635 ,n1024);
    not g1225(n5289 ,n5288);
    not g1226(n934 ,n28[8]);
    buf g1227(n14[4], n10[4]);
    or g1228(n5344 ,n5101 ,n5109);
    not g1229(n5417 ,n5416);
    nor g1230(n1943 ,n1890 ,n1937);
    or g1231(n86 ,n25[6] ,n25[5]);
    nor g1232(n3985 ,n3963 ,n3984);
    not g1233(n5485 ,n5484);
    xnor g1234(n4789 ,n4667 ,n4599);
    nor g1235(n2197 ,n2133 ,n2148);
    nor g1236(n1215 ,n815 ,n642);
    nor g1237(n3267 ,n3092 ,n3178);
    nor g1238(n3375 ,n3303 ,n3350);
    not g1239(n5501 ,n5500);
    xnor g1240(n4391 ,n4062 ,n4070);
    or g1241(n7706 ,n7610 ,n7681);
    nor g1242(n3096 ,n2994 ,n3035);
    xnor g1243(n3666 ,n7804 ,n7781);
    nor g1244(n2604 ,n2442 ,n2548);
    xnor g1245(n351 ,n215 ,n213);
    not g1246(n732 ,n3[4]);
    nor g1247(n3655 ,n3604 ,n3593);
    not g1248(n7422 ,n7727);
    nor g1249(n3422 ,n3316 ,n3391);
    nor g1250(n6332 ,n5714 ,n6212);
    nor g1251(n2612 ,n2431 ,n2574);
    xnor g1252(n4958 ,n4896 ,n4813);
    nor g1253(n4180 ,n4018 ,n4025);
    nor g1254(n7539 ,n7353 ,n7477);
    nor g1255(n5970 ,n5713 ,n5863);
    nor g1256(n2746 ,n2707 ,n2700);
    nor g1257(n2557 ,n2432 ,n2525);
    xnor g1258(n5019 ,n4970 ,n4973);
    nor g1259(n4038 ,n4014 ,n4007);
    not g1260(n7432 ,n7733);
    not g1261(n4780 ,n4779);
    nor g1262(n2409 ,n2374 ,n2408);
    nor g1263(n4439 ,n4259 ,n4290);
    nor g1264(n2015 ,n1893 ,n1976);
    nor g1265(n5660 ,n5492 ,n5198);
    not g1266(n5377 ,n5376);
    nor g1267(n1455 ,n837 ,n634);
    xnor g1268(n6257 ,n5810 ,n5166);
    nor g1269(n558 ,n483 ,n527);
    nor g1270(n1219 ,n823 ,n642);
    nor g1271(n534 ,n409 ,n505);
    nor g1272(n3462 ,n3437 ,n3420);
    nor g1273(n6728 ,n6583 ,n6692);
    nor g1274(n3407 ,n3307 ,n3374);
    nor g1275(n1240 ,n954 ,n637);
    nor g1276(n623 ,n614 ,n622);
    not g1277(n758 ,n5[1]);
    nor g1278(n3196 ,n3099 ,n3172);
    not g1279(n49 ,n37[3]);
    not g1280(n5203 ,n5202);
    dff g1281(.RN(n1), .SN(1'b1), .CK(n0), .D(n1607), .Q(n19[0]));
    not g1282(n864 ,n16[0]);
    nor g1283(n5883 ,n5558 ,n5601);
    nor g1284(n2608 ,n2443 ,n2574);
    nor g1285(n3515 ,n3467 ,n3496);
    xnor g1286(n2806 ,n2652 ,n2770);
    not g1287(n3632 ,n39[3]);
    dff g1288(.RN(n1), .SN(1'b1), .CK(n0), .D(n1737), .Q(n30[4]));
    xor g1289(n4382 ,n4134 ,n4188);
    nor g1290(n7556 ,n7361 ,n7480);
    not g1291(n4055 ,n4054);
    nor g1292(n6344 ,n6065 ,n6222);
    nor g1293(n7603 ,n7454 ,n7476);
    nor g1294(n437 ,n360 ,n371);
    xnor g1295(n600 ,n567 ,n542);
    dff g1296(.RN(n1), .SN(1'b1), .CK(n0), .D(n1689), .Q(n34[1]));
    or g1297(n7685 ,n7627 ,n7626);
    not g1298(n3434 ,n3433);
    nor g1299(n3718 ,n3658 ,n3680);
    xnor g1300(n4936 ,n4857 ,n4760);
    nor g1301(n6218 ,n5227 ,n6048);
    not g1302(n2163 ,n2162);
    or g1303(n7477 ,n26[1] ,n7457);
    nor g1304(n1468 ,n762 ,n639);
    or g1305(n1635 ,n1303 ,n1235);
    nor g1306(n3095 ,n2995 ,n3035);
    nor g1307(n4843 ,n4760 ,n4784);
    nor g1308(n3809 ,n3779 ,n3808);
    nor g1309(n1313 ,n723 ,n636);
    nor g1310(n4914 ,n4889 ,n4881);
    nor g1311(n7535 ,n7333 ,n7481);
    nor g1312(n2057 ,n1890 ,n2003);
    not g1313(n684 ,n21[1]);
    not g1314(n1980 ,n1979);
    dff g1315(.RN(n1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n26[1]));
    nor g1316(n4154 ,n4014 ,n4021);
    not g1317(n645 ,n27[6]);
    nor g1318(n7040 ,n6952 ,n7014);
    not g1319(n210 ,n209);
    xnor g1320(n6288 ,n5992 ,n5936);
    not g1321(n5022 ,n5021);
    nor g1322(n4331 ,n4041 ,n4083);
    xnor g1323(n7806 ,n2316 ,n2358);
    nor g1324(n6669 ,n6487 ,n6561);
    xnor g1325(n6990 ,n6845 ,n6823);
    or g1326(n89 ,n25[7] ,n88);
    not g1327(n7454 ,n7728);
    nor g1328(n3695 ,n3655 ,n3693);
    not g1329(n4017 ,n20[0]);
    xnor g1330(n6418 ,n6072 ,n5745);
    xnor g1331(n2782 ,n2724 ,n2657);
    nor g1332(n4456 ,n4326 ,n4443);
    not g1333(n434 ,n433);
    nor g1334(n1120 ,n634 ,n1090);
    nor g1335(n7247 ,n7214 ,n7225);
    xnor g1336(n6515 ,n6280 ,n6171);
    or g1337(n1007 ,n860 ,n897);
    xor g1338(n2425 ,n2452 ,n2472);
    not g1339(n766 ,n2[0]);
    nor g1340(n6451 ,n6182 ,n6315);
    nor g1341(n6693 ,n6526 ,n6524);
    not g1342(n792 ,n1856);
    nor g1343(n4573 ,n4399 ,n4506);
    nor g1344(n4184 ,n4013 ,n4018);
    not g1345(n4313 ,n4312);
    nor g1346(n1345 ,n892 ,n637);
    xnor g1347(n4379 ,n4064 ,n4164);
    or g1348(n1629 ,n1293 ,n1230);
    xnor g1349(n7759 ,n3951 ,n3992);
    not g1350(n909 ,n24[13]);
    not g1351(n3830 ,n19[5]);
    not g1352(n150 ,n37[6]);
    nor g1353(n2368 ,n2333 ,n2354);
    nor g1354(n1231 ,n648 ,n634);
    nor g1355(n6441 ,n6197 ,n6310);
    nor g1356(n2033 ,n1944 ,n2017);
    not g1357(n5977 ,n5976);
    nor g1358(n1420 ,n886 ,n642);
    nor g1359(n2936 ,n2880 ,n2918);
    nor g1360(n3160 ,n2994 ,n3065);
    xnor g1361(n7811 ,n2401 ,n2412);
    not g1362(n7333 ,n41[7]);
    nor g1363(n3366 ,n3284 ,n3346);
    nor g1364(n2631 ,n2564 ,n2606);
    not g1365(n816 ,n17[5]);
    xnor g1366(n2972 ,n2947 ,n2930);
    nor g1367(n6678 ,n6425 ,n6500);
    or g1368(n977 ,n23[2] ,n23[3]);
    xnor g1369(n4369 ,n4228 ,n4072);
    not g1370(n3600 ,n7806);
    nor g1371(n6324 ,n5995 ,n6232);
    xor g1372(n6397 ,n6166 ,n6078);
    xor g1373(n1846 ,n611 ,n626);
    not g1374(n4872 ,n4871);
    or g1375(n5570 ,n5090 ,n5104);
    nor g1376(n7604 ,n7388 ,n7476);
    not g1377(n3972 ,n3971);
    not g1378(n4868 ,n4867);
    nor g1379(n3942 ,n7788 ,n7773);
    nor g1380(n2742 ,n2667 ,n2427);
    nor g1381(n6586 ,n6386 ,n6466);
    xnor g1382(n2864 ,n2685 ,n2816);
    nor g1383(n3129 ,n3012 ,n3064);
    not g1384(n182 ,n181);
    or g1385(n7629 ,n7515 ,n7528);
    nor g1386(n6773 ,n6653 ,n6647);
    nor g1387(n5681 ,n5281 ,n5149);
    or g1388(n1710 ,n1354 ,n1162);
    nor g1389(n6321 ,n5999 ,n6231);
    not g1390(n258 ,n257);
    xnor g1391(n2213 ,n2152 ,n1885);
    nor g1392(n6890 ,n6774 ,n6816);
    nor g1393(n3301 ,n3155 ,n3259);
    nor g1394(n6016 ,n5757 ,n5838);
    xor g1395(n7793 ,n6069 ,n5450);
    not g1396(n3117 ,n3116);
    nor g1397(n1242 ,n951 ,n637);
    not g1398(n5229 ,n5228);
    nor g1399(n1258 ,n877 ,n638);
    not g1400(n782 ,n2[3]);
    or g1401(n1589 ,n1251 ,n1112);
    nor g1402(n5634 ,n5276 ,n5128);
    or g1403(n1796 ,n1201 ,n1562);
    xnor g1404(n4735 ,n4610 ,n4508);
    nor g1405(n360 ,n184 ,n327);
    not g1406(n6631 ,n6630);
    dff g1407(.RN(n1), .SN(1'b1), .CK(n0), .D(n1657), .Q(n35[8]));
    xnor g1408(n4374 ,n4098 ,n4094);
    or g1409(n5561 ,n5097 ,n5104);
    nor g1410(n4646 ,n4496 ,n4518);
    or g1411(n5548 ,n5090 ,n5105);
    nor g1412(n4447 ,n4268 ,n4275);
    xnor g1413(n7715 ,n39[0] ,n3679);
    nor g1414(n2077 ,n1995 ,n2057);
    not g1415(n4467 ,n4466);
    not g1416(n5467 ,n5466);
    nor g1417(n4748 ,n4637 ,n4700);
    or g1418(n1663 ,n1325 ,n1519);
    nor g1419(n293 ,n185 ,n181);
    dff g1420(.RN(n1), .SN(1'b1), .CK(n0), .D(n1704), .Q(n32[6]));
    nor g1421(n5914 ,n5566 ,n5630);
    nor g1422(n7230 ,n7134 ,n7208);
    nor g1423(n1233 ,n653 ,n634);
    nor g1424(n4470 ,n4342 ,n4429);
    nor g1425(n1957 ,n1894 ,n1937);
    xnor g1426(n2508 ,n2494 ,n2469);
    nor g1427(n302 ,n260 ,n270);
    nor g1428(n2413 ,n2412 ,n2399);
    nor g1429(n6462 ,n6160 ,n6308);
    nor g1430(n4080 ,n4007 ,n4028);
    nor g1431(n3818 ,n3778 ,n3817);
    nor g1432(n3318 ,n3123 ,n3265);
    or g1433(n1732 ,n1372 ,n1186);
    or g1434(n7634 ,n7533 ,n7532);
    nor g1435(n3175 ,n2995 ,n3065);
    not g1436(n5373 ,n5372);
    nor g1437(n1368 ,n671 ,n1103);
    xnor g1438(n6719 ,n6499 ,n6424);
    xnor g1439(n2634 ,n2502 ,n2552);
    nor g1440(n2560 ,n2434 ,n2525);
    nor g1441(n1536 ,n743 ,n641);
    dff g1442(.RN(n1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n28[11]));
    xnor g1443(n2285 ,n2217 ,n1889);
    or g1444(n1778 ,n1417 ,n1503);
    xnor g1445(n2668 ,n2512 ,n2598);
    nor g1446(n267 ,n160 ,n151);
    nor g1447(n422 ,n189 ,n379);
    not g1448(n2476 ,n2477);
    xnor g1449(n4593 ,n4411 ,n4102);
    nor g1450(n2638 ,n2531 ,n2597);
    not g1451(n2999 ,n7751);
    or g1452(n5343 ,n5117 ,n5091);
    not g1453(n855 ,n34[7]);
    xnor g1454(n39[1] ,n2670 ,n2550);
    xor g1455(n7766 ,n3847 ,n3858);
    nor g1456(n1462 ,n795 ,n634);
    xnor g1457(n2706 ,n2514 ,n2645);
    not g1458(n736 ,n1845);
    not g1459(n965 ,n10[11]);
    nor g1460(n7561 ,n7370 ,n7474);
    xnor g1461(n1098 ,n645 ,n819);
    nor g1462(n3653 ,n3603 ,n3596);
    not g1463(n5096 ,n22[7]);
    nor g1464(n2203 ,n2153 ,n2140);
    not g1465(n4978 ,n4977);
    not g1466(n5451 ,n5450);
    not g1467(n708 ,n33[2]);
    nor g1468(n5508 ,n5100 ,n5113);
    xnor g1469(n2774 ,n2727 ,n2707);
    nor g1470(n7507 ,n7417 ,n7478);
    nor g1471(n1138 ,n641 ,n1046);
    nor g1472(n6905 ,n6758 ,n6817);
    xnor g1473(n6084 ,n5820 ,n5841);
    not g1474(n270 ,n269);
    nor g1475(n1441 ,n839 ,n634);
    nor g1476(n5868 ,n5546 ,n5649);
    or g1477(n1750 ,n1390 ,n1171);
    xnor g1478(n6711 ,n6527 ,n6547);
    nor g1479(n6048 ,n5682 ,n5906);
    nor g1480(n3479 ,n3352 ,n3443);
    xor g1481(n38[5] ,n39[5] ,n7841);
    nor g1482(n3120 ,n3013 ,n3034);
    nor g1483(n4758 ,n4650 ,n4703);
    not g1484(n786 ,n1858);
    nor g1485(n3686 ,n3632 ,n3644);
    nor g1486(n4302 ,n4226 ,n4054);
    nor g1487(n1188 ,n1003 ,n1104);
    xnor g1488(n2381 ,n2322 ,n2356);
    xnor g1489(n7167 ,n7111 ,n7081);
    dff g1490(.RN(n1), .SN(1'b1), .CK(n0), .D(n1649), .Q(n10[4]));
    xnor g1491(n3527 ,n3482 ,n3376);
    nor g1492(n5712 ,n5217 ,n5193);
    nor g1493(n5585 ,n5200 ,n5388);
    xor g1494(n41[15] ,n7237 ,n7322);
    or g1495(n1013 ,n887 ,n916);
    not g1496(n124 ,n33[3]);
    xnor g1497(n3343 ,n3108 ,n3223);
    xnor g1498(n530 ,n478 ,n455);
    not g1499(n3702 ,n3701);
    nor g1500(n2747 ,n2657 ,n2724);
    dff g1501(.RN(n1), .SN(1'b1), .CK(n0), .D(n1620), .Q(n11[11]));
    not g1502(n7031 ,n7030);
    nor g1503(n2119 ,n1959 ,n2101);
    or g1504(n36[8] ,n7688 ,n7686);
    nor g1505(n1299 ,n702 ,n636);
    not g1506(n4790 ,n4789);
    nor g1507(n3643 ,n7807 ,n7784);
    not g1508(n5369 ,n5368);
    not g1509(n6867 ,n6866);
    nor g1510(n6066 ,n5675 ,n5918);
    xnor g1511(n1053 ,n647 ,n832);
    nor g1512(n2753 ,n2658 ,n2690);
    nor g1513(n2544 ,n2431 ,n2521);
    xor g1514(n5806 ,n5339 ,n5428);
    not g1515(n797 ,n1865);
    not g1516(n4853 ,n4852);
    nor g1517(n6921 ,n6835 ,n6893);
    or g1518(n1673 ,n1331 ,n1540);
    nor g1519(n6686 ,n6540 ,n6496);
    xnor g1520(n2724 ,n2511 ,n2640);
    not g1521(n508 ,n507);
    nor g1522(n4947 ,n4813 ,n4897);
    dff g1523(.RN(n1), .SN(1'b1), .CK(n0), .D(n1664), .Q(n35[4]));
    xnor g1524(n3075 ,n40[6] ,n7745);
    nor g1525(n5628 ,n5160 ,n5494);
    xnor g1526(n1048 ,n857 ,n818);
    xnor g1527(n4783 ,n4672 ,n4554);
    xnor g1528(n6977 ,n6858 ,n6829);
    nor g1529(n4836 ,n4750 ,n4775);
    nor g1530(n7458 ,n41[12] ,n7820);
    xnor g1531(n3960 ,n7787 ,n7772);
    not g1532(n4535 ,n4534);
    or g1533(n5335 ,n5092 ,n5100);
    not g1534(n5483 ,n5482);
    xnor g1535(n6259 ,n5790 ,n5286);
    not g1536(n5554 ,n5553);
    nor g1537(n7536 ,n7349 ,n7475);
    not g1538(n796 ,n1875);
    not g1539(n795 ,n1872);
    dff g1540(.RN(n1), .SN(1'b1), .CK(n0), .D(n1574), .Q(n25[0]));
    xnor g1541(n6130 ,n5817 ,n5330);
    not g1542(n719 ,n1832);
    xnor g1543(n3899 ,n41[6] ,n7807);
    nor g1544(n4812 ,n4704 ,n4764);
    nor g1545(n2894 ,n2865 ,n2841);
    nor g1546(n2125 ,n1968 ,n2083);
    nor g1547(n3193 ,n3013 ,n3072);
    xnor g1548(n6300 ,n5226 ,n6048);
    nor g1549(n2455 ,n21[2] ,n21[1]);
    or g1550(n1619 ,n1283 ,n1444);
    nor g1551(n3499 ,n3446 ,n3462);
    nor g1552(n3091 ,n3012 ,n3039);
    xor g1553(n2430 ,n2671 ,n2677);
    nor g1554(n7552 ,n7414 ,n7478);
    nor g1555(n3771 ,n3714 ,n3744);
    not g1556(n4248 ,n4247);
    not g1557(n2663 ,n2662);
    nor g1558(n3231 ,n3095 ,n3186);
    not g1559(n4107 ,n4106);
    xnor g1560(n4370 ,n4234 ,n4168);
    nor g1561(n1988 ,n1893 ,n1978);
    or g1562(n1621 ,n1285 ,n1490);
    nor g1563(n195 ,n156 ,n149);
    not g1564(n4687 ,n4686);
    nor g1565(n3924 ,n3894 ,n3923);
    not g1566(n5407 ,n5406);
    nor g1567(n1492 ,n798 ,n639);
    not g1568(n4122 ,n4121);
    not g1569(n1901 ,n37[1]);
    nor g1570(n4327 ,n4175 ,n4209);
    not g1571(n1902 ,n37[6]);
    nor g1572(n5978 ,n5722 ,n5865);
    not g1573(n4982 ,n4981);
    not g1574(n2165 ,n2164);
    nor g1575(n6895 ,n6632 ,n6795);
    nor g1576(n1454 ,n832 ,n634);
    nor g1577(n6308 ,n6265 ,n6253);
    nor g1578(n7528 ,n7714 ,n7475);
    not g1579(n3634 ,n7811);
    nor g1580(n3651 ,n3592 ,n3624);
    not g1581(n6162 ,n6161);
    not g1582(n900 ,n28[11]);
    nor g1583(n1272 ,n864 ,n640);
    nor g1584(n7266 ,n7243 ,n7174);
    or g1585(n5347 ,n5096 ,n5114);
    nor g1586(n619 ,n605 ,n612);
    not g1587(n6906 ,n6905);
    xnor g1588(n6640 ,n6403 ,n6274);
    not g1589(n826 ,n35[3]);
    nor g1590(n392 ,n318 ,n368);
    not g1591(n578 ,n577);
    not g1592(n348 ,n347);
    or g1593(n1699 ,n1348 ,n1462);
    or g1594(n1840 ,n33[6] ,n96);
    nor g1595(n1471 ,n763 ,n639);
    xnor g1596(n4550 ,n4364 ,n4361);
    not g1597(n740 ,n1878);
    xnor g1598(n3355 ,n3122 ,n3265);
    not g1599(n127 ,n33[2]);
    nor g1600(n7177 ,n7123 ,n7153);
    nor g1601(n6610 ,n6527 ,n6519);
    nor g1602(n7598 ,n7328 ,n7481);
    not g1603(n5108 ,n22[6]);
    not g1604(n844 ,n23[0]);
    xor g1605(n7789 ,n5072 ,n5079);
    nor g1606(n5892 ,n5556 ,n5592);
    nor g1607(n5905 ,n5582 ,n5656);
    nor g1608(n71 ,n66 ,n70);
    not g1609(n2432 ,n7765);
    not g1610(n2947 ,n2946);
    nor g1611(n7583 ,n7329 ,n7481);
    xnor g1612(n6618 ,n6395 ,n6183);
    nor g1613(n1187 ,n1005 ,n1104);
    or g1614(n1829 ,n1811 ,n1828);
    not g1615(n3246 ,n3245);
    or g1616(n1794 ,n1204 ,n1561);
    not g1617(n50 ,n19[3]);
    xnor g1618(n2482 ,n21[1] ,n22[1]);
    dff g1619(.RN(n1), .SN(1'b1), .CK(n0), .D(n1650), .Q(n35[13]));
    not g1620(n637 ,n634);
    nor g1621(n4491 ,n4217 ,n4402);
    xnor g1622(n2685 ,n2502 ,n2655);
    not g1623(n5157 ,n5156);
    nor g1624(n6561 ,n6270 ,n6432);
    not g1625(n5471 ,n5470);
    nor g1626(n315 ,n234 ,n172);
    not g1627(n7356 ,n38[2]);
    not g1628(n3240 ,n3239);
    nor g1629(n6269 ,n5708 ,n6009);
    not g1630(n2205 ,n2204);
    nor g1631(n4321 ,n4073 ,n4229);
    not g1632(n4531 ,n4530);
    nor g1633(n2914 ,n2877 ,n2891);
    nor g1634(n5882 ,n5340 ,n5604);
    nor g1635(n1198 ,n1012 ,n1104);
    not g1636(n2483 ,n2482);
    nor g1637(n4807 ,n4631 ,n4722);
    nor g1638(n7517 ,n7372 ,n7479);
    nor g1639(n1140 ,n641 ,n1045);
    nor g1640(n5543 ,n5118 ,n5107);
    nor g1641(n4665 ,n4490 ,n4574);
    nor g1642(n6660 ,n6484 ,n6563);
    nor g1643(n54 ,n37[6] ,n19[6]);
    nor g1644(n5222 ,n5112 ,n5104);
    dff g1645(.RN(n1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n29[2]));
    nor g1646(n6465 ,n6175 ,n6322);
    nor g1647(n7226 ,n7186 ,n7195);
    nor g1648(n143 ,n33[6] ,n141);
    nor g1649(n1260 ,n710 ,n636);
    nor g1650(n107 ,n25[2] ,n105);
    nor g1651(n2601 ,n2443 ,n2549);
    xor g1652(n1887 ,n2114 ,n2125);
    buf g1653(n13[13], n10[13]);
    nor g1654(n1194 ,n1007 ,n1104);
    nor g1655(n3404 ,n3310 ,n3366);
    or g1656(n1771 ,n1408 ,n1134);
    xnor g1657(n6255 ,n5795 ,n5130);
    xnor g1658(n6490 ,n6092 ,n6330);
    xnor g1659(n7728 ,n3553 ,n3548);
    xor g1660(n4368 ,n4140 ,n4224);
    not g1661(n430 ,n429);
    xnor g1662(n6792 ,n6596 ,n6426);
    nor g1663(n3354 ,n3235 ,n3273);
    nor g1664(n6609 ,n6334 ,n6555);
    nor g1665(n3988 ,n3943 ,n3987);
    nor g1666(n3048 ,n2994 ,n3041);
    xor g1667(n7792 ,n5018 ,n5085);
    xnor g1668(n4513 ,n4400 ,n4351);
    nor g1669(n3909 ,n3901 ,n3908);
    nor g1670(n2246 ,n2107 ,n2222);
    nor g1671(n5077 ,n5076 ,n5066);
    not g1672(n4551 ,n4550);
    xnor g1673(n6122 ,n5847 ,n5288);
    xnor g1674(n7805 ,n2317 ,n2302);
    nor g1675(n3755 ,n3696 ,n3733);
    nor g1676(n7197 ,n7104 ,n7184);
    xnor g1677(n6148 ,n5800 ,n5482);
    xnor g1678(n6253 ,n5785 ,n5358);
    not g1679(n5564 ,n5563);
    nor g1680(n6417 ,n6000 ,n6348);
    or g1681(n7610 ,n7607 ,n7606);
    nor g1682(n4837 ,n4712 ,n4811);
    nor g1683(n7564 ,n7399 ,n7475);
    not g1684(n6333 ,n6332);
    or g1685(n1803 ,n1439 ,n1514);
    or g1686(n1086 ,n23[1] ,n977);
    nor g1687(n5452 ,n5115 ,n5102);
    nor g1688(n6372 ,n6151 ,n6083);
    xnor g1689(n6708 ,n6541 ,n6586);
    or g1690(n7625 ,n7551 ,n7550);
    xnor g1691(n6521 ,n6283 ,n6148);
    nor g1692(n5934 ,n5625 ,n5846);
    not g1693(n4203 ,n4202);
    not g1694(n5445 ,n5444);
    nor g1695(n6050 ,n5717 ,n5866);
    nor g1696(n5738 ,n5413 ,n5155);
    nor g1697(n3636 ,n39[8] ,n7809);
    xnor g1698(n3454 ,n3393 ,n3416);
    or g1699(n1717 ,n1359 ,n1558);
    xnor g1700(n1044 ,n866 ,n646);
    dff g1701(.RN(n1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n20[6]));
    not g1702(n6853 ,n6852);
    nor g1703(n3224 ,n3085 ,n3191);
    xnor g1704(n6944 ,n6780 ,n6648);
    xnor g1705(n2515 ,n2492 ,n2480);
    not g1706(n7373 ,n7789);
    xnor g1707(n528 ,n480 ,n458);
    nor g1708(n5240 ,n5091 ,n5094);
    not g1709(n703 ,n19[7]);
    xor g1710(n7751 ,n7813 ,n7790);
    nor g1711(n235 ,n146 ,n148);
    nor g1712(n5593 ,n5132 ,n5482);
    dff g1713(.RN(n1), .SN(1'b1), .CK(n0), .D(n1710), .Q(n32[3]));
    xnor g1714(n6992 ,n6846 ,n6786);
    nor g1715(n471 ,n430 ,n414);
    nor g1716(n6663 ,n6471 ,n6579);
    not g1717(n4692 ,n4691);
    nor g1718(n7103 ,n7005 ,n7048);
    nor g1719(n6670 ,n6428 ,n6567);
    nor g1720(n3235 ,n3115 ,n3141);
    xor g1721(n40[11] ,n39[12] ,n7828);
    nor g1722(n3357 ,n3232 ,n3276);
    not g1723(n2899 ,n2898);
    nor g1724(n5692 ,n5173 ,n5357);
    xnor g1725(n4402 ,n4118 ,n4130);
    nor g1726(n3586 ,n3544 ,n3585);
    nor g1727(n7121 ,n7029 ,n7074);
    not g1728(n4243 ,n4242);
    not g1729(n4354 ,n4353);
    nor g1730(n7175 ,n7114 ,n7150);
    xnor g1731(n3787 ,n3749 ,n3720);
    xnor g1732(n6501 ,n6299 ,n5944);
    nor g1733(n2526 ,n2443 ,n2523);
    nor g1734(n6224 ,n5961 ,n6043);
    nor g1735(n445 ,n422 ,n439);
    nor g1736(n7314 ,n7313 ,n7306);
    not g1737(n937 ,n10[10]);
    nor g1738(n2304 ,n2260 ,n2280);
    not g1739(n6256 ,n6255);
    dff g1740(.RN(n1), .SN(1'b1), .CK(n0), .D(n1633), .Q(n11[2]));
    not g1741(n7442 ,n39[10]);
    nor g1742(n6969 ,n6766 ,n6886);
    nor g1743(n5911 ,n5570 ,n5661);
    not g1744(n5149 ,n5148);
    nor g1745(n1359 ,n890 ,n1107);
    xnor g1746(n2660 ,n2502 ,n2582);
    xnor g1747(n1930 ,n1906 ,n19[6]);
    xnor g1748(n1852 ,n566 ,n554);
    nor g1749(n5700 ,n5493 ,n5199);
    nor g1750(n6685 ,n6497 ,n6572);
    nor g1751(n311 ,n186 ,n182);
    nor g1752(n2358 ,n2311 ,n2328);
    nor g1753(n2618 ,n2441 ,n2547);
    xor g1754(n331 ,n272 ,n233);
    nor g1755(n2337 ,n2202 ,n2307);
    not g1756(n7327 ,n26[2]);
    xor g1757(n7749 ,n7811 ,n7788);
    buf g1758(n14[6], n10[6]);
    nor g1759(n2991 ,n2960 ,n2990);
    not g1760(n2909 ,n2908);
    nor g1761(n5182 ,n5096 ,n5092);
    nor g1762(n3195 ,n3097 ,n3127);
    nor g1763(n6347 ,n6054 ,n6224);
    xnor g1764(n4409 ,n4265 ,n4245);
    nor g1765(n3367 ,n3288 ,n3353);
    nor g1766(n2097 ,n2013 ,n2055);
    not g1767(n1890 ,n37[5]);
    xnor g1768(n7067 ,n6994 ,n6967);
    nor g1769(n3437 ,n3275 ,n3406);
    nor g1770(n2617 ,n2434 ,n2549);
    xor g1771(n7747 ,n7809 ,n7786);
    nor g1772(n2886 ,n2815 ,n2872);
    nor g1773(n1983 ,n1892 ,n1974);
    nor g1774(n6966 ,n6797 ,n6870);
    nor g1775(n3920 ,n3890 ,n3919);
    xnor g1776(n4717 ,n4603 ,n4528);
    xnor g1777(n6656 ,n6404 ,n6163);
    dff g1778(.RN(n1), .SN(1'b1), .CK(n0), .D(n1680), .Q(n34[6]));
    nor g1779(n144 ,n121 ,n142);
    nor g1780(n3290 ,n3157 ,n3216);
    nor g1781(n2055 ,n1893 ,n2003);
    dff g1782(.RN(n1), .SN(1'b1), .CK(n0), .D(n1601), .Q(n12[5]));
    dff g1783(.RN(n1), .SN(1'b1), .CK(n0), .D(n1606), .Q(n19[1]));
    nor g1784(n290 ,n247 ,n187);
    xnor g1785(n2209 ,n2106 ,n2164);
    nor g1786(n5586 ,n5246 ,n5268);
    nor g1787(n2417 ,n2416 ,n2400);
    nor g1788(n2968 ,n2921 ,n2948);
    nor g1789(n7185 ,n7098 ,n7146);
    not g1790(n6244 ,n6243);
    or g1791(n7695 ,n7644 ,n7643);
    xnor g1792(n7164 ,n7118 ,n7135);
    nor g1793(n6903 ,n6629 ,n6832);
    nor g1794(n5866 ,n5314 ,n5603);
    nor g1795(n6236 ,n5973 ,n5939);
    or g1796(n1577 ,n1240 ,n1340);
    nor g1797(n7064 ,n6957 ,n7003);
    nor g1798(n3280 ,n3147 ,n3247);
    xnor g1799(n2466 ,n2436 ,n22[1]);
    nor g1800(n4660 ,n4535 ,n4533);
    nor g1801(n3459 ,n3365 ,n3448);
    not g1802(n7376 ,n40[1]);
    nor g1803(n6443 ,n6274 ,n6323);
    xnor g1804(n2116 ,n1958 ,n2032);
    nor g1805(n7724 ,n3314 ,n3298);
    not g1806(n7421 ,n7759);
    not g1807(n4159 ,n4158);
    nor g1808(n1374 ,n962 ,n1105);
    nor g1809(n4338 ,n4037 ,n4157);
    dff g1810(.RN(n1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n20[3]));
    not g1811(n83 ,n25[4]);
    not g1812(n6651 ,n6650);
    nor g1813(n6759 ,n6641 ,n6638);
    dff g1814(.RN(n1), .SN(1'b1), .CK(n0), .D(n1637), .Q(n10[14]));
    xnor g1815(n4534 ,n4367 ,n4194);
    xnor g1816(n1061 ,n653 ,n861);
    xnor g1817(n6158 ,n5828 ,n5468);
    nor g1818(n1466 ,n803 ,n639);
    xnor g1819(n1847 ,n618 ,n624);
    nor g1820(n513 ,n463 ,n485);
    not g1821(n2719 ,n2718);
    or g1822(n985 ,n27[1] ,n27[2]);
    nor g1823(n5715 ,n5205 ,n5121);
    nor g1824(n3125 ,n3012 ,n3074);
    or g1825(n5339 ,n5108 ,n5109);
    nor g1826(n6363 ,n6011 ,n6186);
    not g1827(n4268 ,n4267);
    nor g1828(n4942 ,n4832 ,n4906);
    not g1829(n4496 ,n4495);
    dff g1830(.RN(n1), .SN(1'b1), .CK(n0), .D(n1724), .Q(n31[3]));
    nor g1831(n2048 ,n1903 ,n2003);
    xnor g1832(n3486 ,n3395 ,n3439);
    not g1833(n7424 ,n7797);
    nor g1834(n2799 ,n2732 ,n2742);
    or g1835(n1742 ,n1380 ,n1192);
    nor g1836(n5130 ,n5099 ,n5090);
    nor g1837(n5988 ,n5710 ,n5872);
    or g1838(n7710 ,n7617 ,n7689);
    nor g1839(n2258 ,n2108 ,n2223);
    not g1840(n7397 ,n7818);
    not g1841(n4128 ,n4127);
    nor g1842(n5724 ,n5191 ,n5355);
    nor g1843(n5727 ,n5189 ,n5147);
    xnor g1844(n7833 ,n3962 ,n3974);
    dff g1845(.RN(n1), .SN(1'b1), .CK(n0), .D(n1605), .Q(n12[3]));
    not g1846(n4710 ,n4709);
    not g1847(n7444 ,n7730);
    not g1848(n5269 ,n5268);
    nor g1849(n2178 ,n2154 ,n2139);
    xnor g1850(n5062 ,n5030 ,n5037);
    nor g1851(n5557 ,n5114 ,n5097);
    nor g1852(n6590 ,n6383 ,n6460);
    nor g1853(n3528 ,n3499 ,n3507);
    nor g1854(n6591 ,n6366 ,n6464);
    nor g1855(n5374 ,n5095 ,n5102);
    not g1856(n260 ,n259);
    nor g1857(n3416 ,n3296 ,n3369);
    nor g1858(n3769 ,n3712 ,n3740);
    nor g1859(n7117 ,n7032 ,n7081);
    nor g1860(n4299 ,n4164 ,n4064);
    not g1861(n5457 ,n5456);
    not g1862(n6019 ,n6018);
    xnor g1863(n2211 ,n2141 ,n2080);
    not g1864(n5125 ,n5124);
    xnor g1865(n2772 ,n2692 ,n2718);
    nor g1866(n1410 ,n663 ,n638);
    nor g1867(n5927 ,n5337 ,n5629);
    not g1868(n6435 ,n6434);
    nor g1869(n1564 ,n873 ,n1103);
    dff g1870(.RN(n1), .SN(1'b1), .CK(n0), .D(n1595), .Q(n12[7]));
    nor g1871(n6696 ,n6390 ,n6534);
    nor g1872(n3756 ,n3704 ,n3727);
    xnor g1873(n4820 ,n4735 ,n4762);
    not g1874(n4594 ,n4593);
    not g1875(n733 ,n1867);
    nor g1876(n2233 ,n2113 ,n2196);
    nor g1877(n5350 ,n5090 ,n5094);
    dff g1878(.RN(n1), .SN(1'b1), .CK(n0), .D(n1592), .Q(n12[9]));
    or g1879(n1774 ,n1413 ,n1501);
    or g1880(n7483 ,n7459 ,n7480);
    nor g1881(n1314 ,n919 ,n636);
    nor g1882(n1346 ,n699 ,n636);
    nor g1883(n4430 ,n4124 ,n4283);
    nor g1884(n4312 ,n4262 ,n4241);
    xnor g1885(n4366 ,n4082 ,n4040);
    nor g1886(n2498 ,n2432 ,n2477);
    not g1887(n4685 ,n4684);
    not g1888(n1903 ,n37[4]);
    nor g1889(n4760 ,n4660 ,n4679);
    nor g1890(n1214 ,n826 ,n1101);
    xnor g1891(n3844 ,n37[6] ,n19[6]);
    nor g1892(n3191 ,n3013 ,n3068);
    nor g1893(n4328 ,n4071 ,n4063);
    nor g1894(n3530 ,n3489 ,n3505);
    or g1895(n1006 ,n666 ,n657);
    or g1896(n1830 ,n1825 ,n1829);
    not g1897(n7172 ,n7171);
    not g1898(n5363 ,n5362);
    nor g1899(n2733 ,n2671 ,n2678);
    not g1900(n4126 ,n4125);
    nor g1901(n2335 ,n1888 ,n2296);
    xor g1902(n4396 ,n4253 ,n4174);
    nor g1903(n5341 ,n5112 ,n5094);
    nor g1904(n3180 ,n3013 ,n3063);
    not g1905(n2933 ,n2932);
    xnor g1906(n6120 ,n5766 ,n5350);
    xnor g1907(n2117 ,n1958 ,n2030);
    not g1908(n531 ,n530);
    dff g1909(.RN(n1), .SN(1'b1), .CK(n0), .D(n1619), .Q(n11[12]));
    not g1910(n5397 ,n5396);
    nor g1911(n2253 ,n2180 ,n2233);
    nor g1912(n3742 ,n39[1] ,n3716);
    nor g1913(n4753 ,n4709 ,n4626);
    not g1914(n6474 ,n6473);
    not g1915(n5475 ,n5474);
    nor g1916(n568 ,n551 ,n554);
    dff g1917(.RN(n1), .SN(1'b1), .CK(n0), .D(n1672), .Q(n34[14]));
    nor g1918(n7295 ,n7262 ,n7285);
    or g1919(n1625 ,n1291 ,n1492);
    nor g1920(n7188 ,n7062 ,n7142);
    or g1921(n7620 ,n7535 ,n7512);
    nor g1922(n4910 ,n4850 ,n4890);
    nor g1923(n2930 ,n2894 ,n2915);
    nor g1924(n6005 ,n5740 ,n5886);
    xnor g1925(n1865 ,n63 ,n57);
    not g1926(n4931 ,n4930);
    not g1927(n1898 ,n19[6]);
    xnor g1928(n2672 ,n2511 ,n2600);
    nor g1929(n4432 ,n4269 ,n4292);
    xor g1930(n5793 ,n5582 ,n5376);
    nor g1931(n3194 ,n2995 ,n3066);
    nor g1932(n3306 ,n3158 ,n3244);
    nor g1933(n5087 ,n4994 ,n5086);
    xnor g1934(n3379 ,n3327 ,n3354);
    nor g1935(n5524 ,n5118 ,n5089);
    not g1936(n3007 ,n7739);
    nor g1937(n2918 ,n2783 ,n2890);
    not g1938(n4980 ,n4979);
    not g1939(n7399 ,n38[3]);
    nor g1940(n3936 ,n7780 ,n38[3]);
    not g1941(n5249 ,n5248);
    xor g1942(n7750 ,n7812 ,n7789);
    nor g1943(n6360 ,n5948 ,n6125);
    not g1944(n2433 ,n7767);
    not g1945(n776 ,n1848);
    nor g1946(n7838 ,n3950 ,n3949);
    nor g1947(n3564 ,n3520 ,n3536);
    nor g1948(n3178 ,n2995 ,n3063);
    not g1949(n4209 ,n4208);
    nor g1950(n6193 ,n5852 ,n6066);
    nor g1951(n6740 ,n6556 ,n6609);
    nor g1952(n6493 ,n6373 ,n6449);
    not g1953(n4211 ,n4210);
    nor g1954(n3212 ,n3050 ,n3136);
    not g1955(n659 ,n36[6]);
    xnor g1956(n4688 ,n4515 ,n4472);
    xnor g1957(n584 ,n544 ,n528);
    nor g1958(n5066 ,n5035 ,n5051);
    not g1959(n2286 ,n2285);
    nor g1960(n5614 ,n5152 ,n5486);
    nor g1961(n3880 ,n7813 ,n41[12]);
    not g1962(n7343 ,n7803);
    nor g1963(n1316 ,n695 ,n637);
    not g1964(n5449 ,n5448);
    dff g1965(.RN(n1), .SN(1'b1), .CK(n0), .D(n1661), .Q(n35[5]));
    not g1966(n3426 ,n3425);
    xor g1967(n6182 ,n5775 ,n5571);
    not g1968(n902 ,n11[3]);
    not g1969(n2363 ,n2362);
    nor g1970(n4566 ,n4457 ,n4465);
    not g1971(n5271 ,n5270);
    nor g1972(n486 ,n458 ,n470);
    nor g1973(n4240 ,n4015 ,n4007);
    not g1974(n4018 ,n37[0]);
    nor g1975(n7723 ,n2994 ,n3074);
    nor g1976(n3295 ,n3105 ,n3241);
    not g1977(n5951 ,n5950);
    nor g1978(n4863 ,n4801 ,n4841);
    xnor g1979(n7290 ,n7254 ,n7227);
    nor g1980(n3649 ,n7802 ,n7779);
    xnor g1981(n7818 ,n3794 ,n3821);
    not g1982(n828 ,n34[9]);
    nor g1983(n3439 ,n3272 ,n3404);
    xnor g1984(n4855 ,n4777 ,n4731);
    xnor g1985(n501 ,n442 ,n433);
    not g1986(n154 ,n37[1]);
    xnor g1987(n1042 ,n36[14] ,n34[14]);
    nor g1988(n3173 ,n2995 ,n3074);
    not g1989(n4023 ,n19[3]);
    nor g1990(n4568 ,n4460 ,n4501);
    nor g1991(n5428 ,n5096 ,n5110);
    not g1992(n6157 ,n6156);
    not g1993(n959 ,n25[7]);
    xnor g1994(n6883 ,n6709 ,n6583);
    nor g1995(n2872 ,n2811 ,n2833);
    nor g1996(n6355 ,n6147 ,n6144);
    nor g1997(n3851 ,n3834 ,n3850);
    or g1998(n5517 ,n5101 ,n5107);
    nor g1999(n3948 ,n7783 ,n38[6]);
    nor g2000(n1818 ,n1102 ,n1813);
    or g2001(n5346 ,n5093 ,n5111);
    xor g2002(n4376 ,n4137 ,n4218);
    nor g2003(n1220 ,n649 ,n1101);
    not g2004(n665 ,n35[0]);
    or g2005(n1705 ,n1209 ,n1533);
    not g2006(n2931 ,n2930);
    nor g2007(n2294 ,n1887 ,n2275);
    nor g2008(n4300 ,n4072 ,n4228);
    not g2009(n5481 ,n5480);
    nor g2010(n199 ,n159 ,n153);
    xnor g2011(n409 ,n335 ,n329);
    nor g2012(n5956 ,n5729 ,n5901);
    nor g2013(n4442 ,n4305 ,n4362);
    nor g2014(n189 ,n156 ,n148);
    xnor g2015(n7771 ,n3890 ,n3919);
    nor g2016(n7154 ,n7042 ,n7130);
    not g2017(n4009 ,n20[4]);
    nor g2018(n2487 ,n2431 ,n2477);
    not g2019(n226 ,n225);
    nor g2020(n1917 ,n19[2] ,n19[1]);
    not g2021(n760 ,n6[3]);
    not g2022(n915 ,n11[4]);
    not g2023(n847 ,n34[3]);
    nor g2024(n5645 ,n5498 ,n5478);
    not g2025(n3614 ,n7808);
    or g2026(n1000 ,n652 ,n650);
    xnor g2027(n6286 ,n5970 ,n6020);
    nor g2028(n2001 ,n1891 ,n1976);
    xor g2029(n5822 ,n5542 ,n5168);
    dff g2030(.RN(n1), .SN(1'b1), .CK(n0), .D(n1693), .Q(n33[6]));
    not g2031(n4028 ,n20[3]);
    nor g2032(n5332 ,n5089 ,n5100);
    not g2033(n7349 ,n38[4]);
    or g2034(n7482 ,n7458 ,n7480);
    xnor g2035(n7782 ,n4958 ,n4917);
    xnor g2036(n4821 ,n4526 ,n4739);
    nor g2037(n1236 ,n660 ,n634);
    nor g2038(n6704 ,n6367 ,n6552);
    not g2039(n3157 ,n3156);
    nor g2040(n6962 ,n6791 ,n6861);
    nor g2041(n6313 ,n6003 ,n6228);
    nor g2042(n1421 ,n677 ,n642);
    nor g2043(n2040 ,n1901 ,n2004);
    not g2044(n576 ,n575);
    nor g2045(n6274 ,n5692 ,n5935);
    not g2046(n6021 ,n6020);
    or g2047(n1089 ,n17[1] ,n990);
    nor g2048(n7003 ,n6842 ,n6956);
    nor g2049(n5707 ,n5499 ,n5479);
    xnor g2050(n344 ,n257 ,n203);
    nor g2051(n7593 ,n7364 ,n7477);
    or g2052(n1591 ,n1254 ,n1475);
    not g2053(n5151 ,n5150);
    not g2054(n268 ,n267);
    or g2055(n1810 ,n1343 ,n1457);
    not g2056(n3026 ,n7747);
    nor g2057(n3208 ,n3098 ,n3134);
    xnor g2058(n6110 ,n5825 ,n5326);
    xor g2059(n2428 ,n2668 ,n2726);
    nor g2060(n3884 ,n3870 ,n3866);
    nor g2061(n4218 ,n4008 ,n4028);
    nor g2062(n1496 ,n753 ,n639);
    nor g2063(n7194 ,n7185 ,n7180);
    buf g2064(n13[7], n11[7]);
    not g2065(n850 ,n22[0]);
    nor g2066(n4484 ,n4351 ,n4401);
    xnor g2067(n2155 ,n1972 ,n2089);
    xnor g2068(n4919 ,n4891 ,n4852);
    not g2069(n729 ,n1861);
    nor g2070(n4112 ,n4021 ,n4016);
    xnor g2071(n3783 ,n3731 ,n3705);
    nor g2072(n4622 ,n4585 ,n4589);
    nor g2073(n6060 ,n5672 ,n5900);
    not g2074(n651 ,n17[1]);
    nor g2075(n6030 ,n5716 ,n5887);
    nor g2076(n6899 ,n6643 ,n6823);
    xnor g2077(n6932 ,n6785 ,n6585);
    xnor g2078(n2137 ,n1970 ,n2069);
    nor g2079(n6747 ,n6548 ,n6693);
    not g2080(n5183 ,n5182);
    not g2081(n4601 ,n4600);
    not g2082(n4755 ,n4754);
    not g2083(n6075 ,n6074);
    xnor g2084(n7827 ,n3952 ,n3986);
    nor g2085(n3150 ,n2994 ,n3077);
    nor g2086(n3472 ,n3436 ,n3442);
    xnor g2087(n7808 ,n2380 ,n2403);
    not g2088(n2723 ,n2722);
    nor g2089(n3641 ,n7808 ,n7785);
    xnor g2090(n3509 ,n3457 ,n3379);
    xnor g2091(n5847 ,n5464 ,n5444);
    or g2092(n7323 ,n7327 ,n7391);
    not g2093(n1928 ,n1927);
    xnor g2094(n2380 ,n2350 ,n2337);
    xnor g2095(n6978 ,n6796 ,n6911);
    nor g2096(n5749 ,n5523 ,n5514);
    nor g2097(n4743 ,n4659 ,n4699);
    nor g2098(n6349 ,n5950 ,n6119);
    nor g2099(n7554 ,n7407 ,n7476);
    nor g2100(n6585 ,n6355 ,n6444);
    not g2101(n711 ,n30[3]);
    not g2102(n7277 ,n7276);
    xnor g2103(n6134 ,n5778 ,n5394);
    xnor g2104(n441 ,n324 ,n381);
    not g2105(n961 ,n25[1]);
    nor g2106(n6817 ,n6582 ,n6757);
    xnor g2107(n3325 ,n3196 ,n3195);
    xnor g2108(n65 ,n37[5] ,n19[5]);
    nor g2109(n4412 ,n4096 ,n4357);
    nor g2110(n1546 ,n922 ,n641);
    xnor g2111(n2771 ,n2665 ,n2722);
    nor g2112(n5360 ,n5114 ,n5091);
    nor g2113(n4800 ,n4684 ,n4718);
    not g2114(n3254 ,n3253);
    nor g2115(n2079 ,n1993 ,n2061);
    not g2116(n3826 ,n37[5]);
    not g2117(n4142 ,n4141);
    or g2118(n1751 ,n1391 ,n1154);
    nor g2119(n3264 ,n3089 ,n3193);
    not g2120(n861 ,n32[3]);
    nor g2121(n7522 ,n7415 ,n7477);
    not g2122(n5298 ,n5297);
    nor g2123(n3837 ,n37[0] ,n19[0]);
    nor g2124(n4317 ,n4185 ,n4159);
    nor g2125(n5033 ,n5013 ,n5027);
    nor g2126(n6987 ,n6811 ,n6960);
    not g2127(n3536 ,n3535);
    nor g2128(n1366 ,n881 ,n1107);
    xnor g2129(n7238 ,n7202 ,n7157);
    nor g2130(n2196 ,n2081 ,n2142);
    nor g2131(n6562 ,n6269 ,n6433);
    nor g2132(n7542 ,n7368 ,n7474);
    xnor g2133(n7256 ,n7224 ,n7214);
    nor g2134(n1289 ,n974 ,n638);
    not g2135(n3631 ,n7778);
    nor g2136(n3148 ,n2994 ,n3067);
    nor g2137(n1503 ,n780 ,n639);
    xnor g2138(n7085 ,n6979 ,n6876);
    xor g2139(n5796 ,n5568 ,n5452);
    nor g2140(n5470 ,n5092 ,n5098);
    nor g2141(n4084 ,n4023 ,n4018);
    not g2142(n6851 ,n6850);
    not g2143(n7263 ,n7262);
    not g2144(n2945 ,n2944);
    nor g2145(n4737 ,n4642 ,n4677);
    nor g2146(n7502 ,n7444 ,n7476);
    not g2147(n5437 ,n5436);
    nor g2148(n5696 ,n5235 ,n5467);
    nor g2149(n2982 ,n2954 ,n2981);
    nor g2150(n7219 ,n7204 ,n7207);
    nor g2151(n3314 ,n3165 ,n3268);
    xnor g2152(n4938 ,n4858 ,n4836);
    nor g2153(n4186 ,n4008 ,n4026);
    nor g2154(n425 ,n190 ,n378);
    xor g2155(n40[7] ,n39[8] ,n7832);
    or g2156(n1588 ,n1252 ,n1474);
    not g2157(n2813 ,n2812);
    xnor g2158(n4516 ,n4410 ,n4080);
    not g2159(n7252 ,n7251);
    nor g2160(n447 ,n429 ,n413);
    xnor g2161(n3067 ,n40[9] ,n7748);
    not g2162(n7410 ,n38[6]);
    nor g2163(n3053 ,n2994 ,n3034);
    xor g2164(n40[0] ,n38[0] ,n39[1]);
    nor g2165(n3054 ,n2994 ,n3040);
    nor g2166(n3823 ,n3770 ,n3822);
    not g2167(n2171 ,n2170);
    not g2168(n3627 ,n7786);
    or g2169(n1630 ,n1294 ,n1231);
    nor g2170(n4892 ,n4808 ,n4839);
    not g2171(n6574 ,n6573);
    nor g2172(n6548 ,n6380 ,n6455);
    nor g2173(n5176 ,n5101 ,n5089);
    not g2174(n6970 ,n6969);
    nor g2175(n6315 ,n6136 ,n6122);
    nor g2176(n4909 ,n4791 ,n4875);
    not g2177(n7261 ,n7260);
    not g2178(n5544 ,n5543);
    nor g2179(n7305 ,n7298 ,n7291);
    nor g2180(n5074 ,n5059 ,n5073);
    nor g2181(n7495 ,n7408 ,n7474);
    nor g2182(n5693 ,n5201 ,n5389);
    not g2183(n379 ,n378);
    nor g2184(n7497 ,n7402 ,n7480);
    xor g2185(n38[4] ,n39[4] ,n7842);
    nor g2186(n4417 ,n4243 ,n4291);
    xnor g2187(n597 ,n532 ,n575);
    or g2188(n1666 ,n1214 ,n1155);
    xnor g2189(n5812 ,n5404 ,n5238);
    nor g2190(n5658 ,n5370 ,n5168);
    nor g2191(n5683 ,n5177 ,n5245);
    not g2192(n4788 ,n4787);
    nor g2193(n2978 ,n2934 ,n2975);
    not g2194(n5116 ,n21[6]);
    or g2195(n5567 ,n5108 ,n5104);
    nor g2196(n6391 ,n6012 ,n6196);
    not g2197(n654 ,n35[5]);
    xnor g2198(n2266 ,n2108 ,n2222);
    xnor g2199(n3848 ,n37[2] ,n19[2]);
    xnor g2200(n6654 ,n6405 ,n6140);
    nor g2201(n6322 ,n6096 ,n6074);
    not g2202(n3480 ,n3479);
    or g2203(n7635 ,n7538 ,n7537);
    nor g2204(n6608 ,n6420 ,n6501);
    not g2205(n6993 ,n6992);
    xor g2206(n7796 ,n7024 ,n7023);
    nor g2207(n4462 ,n4322 ,n4416);
    dff g2208(.RN(n1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n21[1]));
    nor g2209(n4915 ,n4846 ,n4876);
    nor g2210(n3986 ,n3942 ,n3985);
    xor g2211(n5826 ,n5338 ,n5200);
    or g2212(n7489 ,n7463 ,n7480);
    xnor g2213(n2835 ,n2773 ,n2805);
    not g2214(n5171 ,n5170);
    nor g2215(n6008 ,n5652 ,n5842);
    nor g2216(n3458 ,n3439 ,n3421);
    xnor g2217(n7200 ,n7137 ,n7161);
    not g2218(n5165 ,n5164);
    or g2219(n1692 ,n989 ,n1183);
    nor g2220(n3164 ,n2994 ,n3063);
    xnor g2221(n7075 ,n6980 ,n6944);
    nor g2222(n6046 ,n5673 ,n5868);
    xnor g2223(n5030 ,n4983 ,n4992);
    nor g2224(n3913 ,n3879 ,n3912);
    nor g2225(n7129 ,n7078 ,n7076);
    not g2226(n2144 ,n2143);
    xnor g2227(n6280 ,n5988 ,n5990);
    not g2228(n3601 ,n7809);
    nor g2229(n5506 ,n5108 ,n5117);
    xnor g2230(n1927 ,n1909 ,n19[7]);
    not g2231(n5092 ,n37[5]);
    nor g2232(n6015 ,n5748 ,n5835);
    nor g2233(n589 ,n532 ,n576);
    nor g2234(n7283 ,n7260 ,n7252);
    nor g2235(n2791 ,n2634 ,n2764);
    nor g2236(n4489 ,n4360 ,n4404);
    nor g2237(n6057 ,n5706 ,n5892);
    xor g2238(n7765 ,n3846 ,n3856);
    nor g2239(n2607 ,n2432 ,n2574);
    xnor g2240(n39[4] ,n2884 ,n2869);
    nor g2241(n5579 ,n5108 ,n5113);
    or g2242(n36[13] ,n7703 ,n7712);
    nor g2243(n424 ,n392 ,n389);
    not g2244(n1976 ,n1975);
    nor g2245(n7527 ,n7429 ,n7474);
    dff g2246(.RN(n1), .SN(1'b1), .CK(n0), .D(n1613), .Q(n1836));
    or g2247(n271 ,n146 ,n151);
    nor g2248(n5448 ,n5097 ,n5109);
    not g2249(n672 ,n20[7]);
    xnor g2250(n2884 ,n2843 ,n2765);
    not g2251(n5327 ,n5326);
    nor g2252(n6354 ,n6146 ,n6145);
    not g2253(n4814 ,n4813);
    not g2254(n3934 ,n38[1]);
    not g2255(n5439 ,n5438);
    nor g2256(n5571 ,n5112 ,n5119);
    xor g2257(n1884 ,n1972 ,n2082);
    xnor g2258(n7836 ,n3957 ,n3966);
    or g2259(n1614 ,n1277 ,n1441);
    nor g2260(n4954 ,n4879 ,n4909);
    dff g2261(.RN(n1), .SN(1'b1), .CK(n0), .D(n1632), .Q(n11[3]));
    nor g2262(n4286 ,n4088 ,n4196);
    not g2263(n266 ,n265);
    nor g2264(n1223 ,n820 ,n1105);
    xor g2265(n40[14] ,n39[15] ,n7825);
    xnor g2266(n5014 ,n4924 ,n4984);
    xnor g2267(n1970 ,n1947 ,n1925);
    nor g2268(n6837 ,n6670 ,n6730);
    or g2269(n5555 ,n5102 ,n5093);
    nor g2270(n6768 ,n6537 ,n6613);
    nor g2271(n4226 ,n4023 ,n4021);
    not g2272(n2687 ,n2686);
    nor g2273(n2758 ,n2706 ,n2701);
    nor g2274(n2537 ,n2442 ,n2523);
    nor g2275(n7095 ,n6970 ,n7065);
    nor g2276(n3758 ,n3706 ,n3731);
    or g2277(n1797 ,n1205 ,n1563);
    nor g2278(n4272 ,n4092 ,n4230);
    xnor g2279(n6396 ,n6128 ,n6126);
    nor g2280(n2415 ,n2414 ,n2405);
    xnor g2281(n4585 ,n4365 ,n4256);
    nor g2282(n1487 ,n765 ,n639);
    xnor g2283(n3427 ,n3334 ,n3366);
    not g2284(n4026 ,n20[2]);
    nor g2285(n7019 ,n6888 ,n6946);
    xnor g2286(n6112 ,n5770 ,n5543);
    xnor g2287(n6071 ,n5930 ,n5741);
    nor g2288(n4950 ,n4852 ,n4904);
    or g2289(n7709 ,n7631 ,n7678);
    nor g2290(n3996 ,n37[0] ,n20[0]);
    not g2291(n6736 ,n6735);
    not g2292(n4740 ,n4739);
    not g2293(n5459 ,n5458);
    nor g2294(n5326 ,n5117 ,n5103);
    nor g2295(n1411 ,n678 ,n642);
    nor g2296(n7161 ,n7092 ,n7116);
    dff g2297(.RN(n1), .SN(1'b1), .CK(n0), .D(n1702), .Q(n32[7]));
    not g2298(n6865 ,n6864);
    nor g2299(n423 ,n293 ,n383);
    not g2300(n7433 ,n7724);
    nor g2301(n3519 ,n3473 ,n3488);
    or g2302(n5510 ,n5096 ,n5099);
    or g2303(n1763 ,n1402 ,n1545);
    nor g2304(n5006 ,n4932 ,n4974);
    nor g2305(n2655 ,n2559 ,n2612);
    nor g2306(n6232 ,n6033 ,n5985);
    nor g2307(n367 ,n280 ,n286);
    xnor g2308(n6616 ,n6394 ,n6273);
    nor g2309(n1170 ,n1102 ,n1034);
    not g2310(n6113 ,n6112);
    not g2311(n669 ,n20[3]);
    xnor g2312(n4384 ,n4048 ,n4202);
    nor g2313(n5430 ,n5088 ,n5092);
    nor g2314(n4490 ,n4352 ,n4400);
    nor g2315(n6565 ,n6388 ,n6468);
    nor g2316(n7547 ,n7443 ,n7476);
    nor g2317(n6461 ,n6092 ,n6331);
    nor g2318(n1522 ,n748 ,n641);
    not g2319(n5261 ,n5260);
    nor g2320(n4423 ,n4257 ,n4277);
    nor g2321(n131 ,n33[2] ,n129);
    xnor g2322(n6082 ,n5762 ,n5260);
    nor g2323(n2022 ,n1894 ,n1980);
    nor g2324(n421 ,n289 ,n393);
    not g2325(n2651 ,n2652);
    nor g2326(n494 ,n382 ,n466);
    xnor g2327(n332 ,n239 ,n169);
    xnor g2328(n5845 ,n5295 ,n5575);
    nor g2329(n5964 ,n5684 ,n5912);
    xnor g2330(n7216 ,n7171 ,n7132);
    nor g2331(n111 ,n100 ,n109);
    nor g2332(n7186 ,n7040 ,n7144);
    nor g2333(n6687 ,n6431 ,n6510);
    nor g2334(n1148 ,n1100 ,n1071);
    not g2335(n5233 ,n5232);
    not g2336(n5113 ,n19[0]);
    nor g2337(n6668 ,n6475 ,n6513);
    nor g2338(n7550 ,n7341 ,n7474);
    nor g2339(n5400 ,n5115 ,n5092);
    nor g2340(n3049 ,n2994 ,n3033);
    not g2341(n835 ,n20[4]);
    nor g2342(n2854 ,n2740 ,n2808);
    not g2343(n4929 ,n4928);
    not g2344(n3715 ,n3714);
    nor g2345(n1169 ,n1102 ,n1036);
    or g2346(n5311 ,n5108 ,n5089);
    xor g2347(n6160 ,n5764 ,n5190);
    nor g2348(n2182 ,n2110 ,n1884);
    nor g2349(n6017 ,n5747 ,n5836);
    nor g2350(n7053 ,n6997 ,n6990);
    nor g2351(n4424 ,n4244 ,n4294);
    dff g2352(.RN(n1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n17[0]));
    dff g2353(.RN(n1), .SN(1'b1), .CK(n0), .D(n1670), .Q(n35[0]));
    nor g2354(n6452 ,n6179 ,n6317);
    not g2355(n3748 ,n3747);
    not g2356(n5441 ,n5440);
    xor g2357(n1860 ,n62 ,n78);
    xnor g2358(n5848 ,n5540 ,n5178);
    not g2359(n6137 ,n6136);
    nor g2360(n372 ,n288 ,n351);
    nor g2361(n1122 ,n635 ,n1019);
    xnor g2362(n2349 ,n2291 ,n2275);
    nor g2363(n3563 ,n3524 ,n3540);
    or g2364(n3028 ,n3019 ,n3027);
    or g2365(n5581 ,n5092 ,n5103);
    nor g2366(n1912 ,n19[1] ,n20[1]);
    nor g2367(n4678 ,n4509 ,n4641);
    or g2368(n1579 ,n1245 ,n1470);
    xnor g2369(n7826 ,n3956 ,n3988);
    or g2370(n96 ,n33[7] ,n95);
    xnor g2371(n403 ,n341 ,n351);
    xnor g2372(n2948 ,n2904 ,n2854);
    nor g2373(n3365 ,n3291 ,n3345);
    xnor g2374(n7193 ,n7141 ,n7062);
    nor g2375(n4801 ,n4737 ,n4726);
    not g2376(n6512 ,n6511);
    nor g2377(n5904 ,n5517 ,n5644);
    or g2378(n3039 ,n3017 ,n2997);
    nor g2379(n6209 ,n6040 ,n5942);
    not g2380(n7076 ,n7075);
    not g2381(n5239 ,n5238);
    nor g2382(n3288 ,n3111 ,n3210);
    nor g2383(n2575 ,n2443 ,n2517);
    nor g2384(n4825 ,n4743 ,n4807);
    not g2385(n4227 ,n4226);
    nor g2386(n6338 ,n6104 ,n6110);
    xnor g2387(n6632 ,n6397 ,n6100);
    nor g2388(n5045 ,n4987 ,n5021);
    not g2389(n3256 ,n3255);
    xnor g2390(n3679 ,n7801 ,n7778);
    or g2391(n1738 ,n1378 ,n1168);
    xnor g2392(n6850 ,n6717 ,n6612);
    not g2393(n436 ,n435);
    nor g2394(n3417 ,n3283 ,n3362);
    nor g2395(n6888 ,n6827 ,n6808);
    not g2396(n5091 ,n21[5]);
    dff g2397(.RN(n1), .SN(1'b1), .CK(n0), .D(n1644), .Q(n10[7]));
    xnor g2398(n2812 ,n2652 ,n2768);
    not g2399(n4350 ,n4349);
    nor g2400(n6028 ,n5704 ,n5895);
    nor g2401(n1552 ,n911 ,n1100);
    not g2402(n807 ,n1860);
    nor g2403(n3056 ,n3012 ,n3037);
    nor g2404(n296 ,n165 ,n249);
    nor g2405(n4877 ,n4793 ,n4847);
    nor g2406(n569 ,n510 ,n561);
    nor g2407(n2822 ,n2770 ,n2794);
    xor g2408(n1855 ,n396 ,n328);
    not g2409(n931 ,n29[2]);
    nor g2410(n3112 ,n3013 ,n3032);
    not g2411(n7435 ,n7795);
    xnor g2412(n7309 ,n7290 ,n7298);
    or g2413(n1805 ,n1440 ,n1516);
    not g2414(n5135 ,n5134);
    nor g2415(n5043 ,n4997 ,n5023);
    nor g2416(n5859 ,n5518 ,n5620);
    not g2417(n4183 ,n4182);
    nor g2418(n3078 ,n3013 ,n3031);
    not g2419(n7409 ,n7719);
    or g2420(n1608 ,n1269 ,n1118);
    nor g2421(n6234 ,n6029 ,n6027);
    nor g2422(n5146 ,n5088 ,n5106);
    not g2423(n2240 ,n2239);
    xnor g2424(n3678 ,n7806 ,n7783);
    nor g2425(n3573 ,n3541 ,n3572);
    xnor g2426(n2696 ,n2514 ,n2639);
    not g2427(n2834 ,n2833);
    xnor g2428(n610 ,n584 ,n591);
    nor g2429(n7276 ,n7257 ,n7245);
    xnor g2430(n3731 ,n39[3] ,n3666);
    xnor g2431(n1047 ,n655 ,n855);
    not g2432(n5281 ,n5280);
    not g2433(n4527 ,n4526);
    nor g2434(n5083 ,n5056 ,n5082);
    nor g2435(n2028 ,n1892 ,n1978);
    not g2436(n2136 ,n2135);
    not g2437(n6437 ,n6436);
    or g2438(n7702 ,n7658 ,n7656);
    not g2439(n6037 ,n6036);
    nor g2440(n5734 ,n5403 ,n5251);
    nor g2441(n6814 ,n6739 ,n6733);
    xor g2442(n5814 ,n5533 ,n5440);
    nor g2443(n4296 ,n4174 ,n4208);
    nor g2444(n4293 ,n4184 ,n4158);
    not g2445(n5523 ,n5522);
    not g2446(n1974 ,n1973);
    nor g2447(n6774 ,n6562 ,n6669);
    not g2448(n823 ,n24[2]);
    nor g2449(n2388 ,n2369 ,n2365);
    nor g2450(n1456 ,n662 ,n634);
    nor g2451(n1216 ,n822 ,n642);
    or g2452(n1597 ,n1259 ,n1478);
    not g2453(n5111 ,n19[2]);
    xnor g2454(n3745 ,n39[8] ,n3675);
    nor g2455(n5627 ,n5186 ,n5390);
    nor g2456(n2486 ,n2434 ,n2477);
    nor g2457(n3266 ,n3079 ,n3188);
    not g2458(n644 ,n18[1]);
    nor g2459(n518 ,n471 ,n489);
    xnor g2460(n6646 ,n6412 ,n6084);
    nor g2461(n5023 ,n5012 ,n5004);
    nor g2462(n4208 ,n4008 ,n4017);
    nor g2463(n5196 ,n5112 ,n5107);
    nor g2464(n5315 ,n5096 ,n5113);
    not g2465(n6250 ,n6249);
    not g2466(n2386 ,n2385);
    nor g2467(n5679 ,n5359 ,n5249);
    not g2468(n7352 ,n7776);
    nor g2469(n6378 ,n6262 ,n6133);
    xnor g2470(n3791 ,n3737 ,n3722);
    or g2471(n1672 ,n1361 ,n1572);
    nor g2472(n6223 ,n5959 ,n5963);
    nor g2473(n261 ,n147 ,n152);
    not g2474(n4061 ,n4060);
    not g2475(n2274 ,n1886);
    xor g2476(n4385 ,n4260 ,n4092);
    not g2477(n418 ,n417);
    or g2478(n7645 ,n7556 ,n7554);
    xnor g2479(n6285 ,n5966 ,n6022);
    not g2480(n7404 ,n39[0]);
    not g2481(n897 ,n29[4]);
    nor g2482(n4773 ,n4630 ,n4721);
    xnor g2483(n7719 ,n3784 ,n3809);
    nor g2484(n3741 ,n3599 ,n3717);
    nor g2485(n6352 ,n5975 ,n6148);
    not g2486(n1909 ,n20[7]);
    not g2487(n4020 ,n37[6]);
    xnor g2488(n499 ,n453 ,n191);
    nor g2489(n2190 ,n2102 ,n2167);
    or g2490(n1817 ,n1136 ,n1812);
    nor g2491(n462 ,n390 ,n416);
    nor g2492(n4696 ,n4473 ,n4655);
    nor g2493(n5714 ,n5247 ,n5269);
    not g2494(n7018 ,n7017);
    or g2495(n1804 ,n1432 ,n1512);
    nor g2496(n2397 ,n2351 ,n2391);
    not g2497(n4907 ,n4906);
    nor g2498(n1511 ,n773 ,n639);
    not g2499(n698 ,n10[7]);
    nor g2500(n5426 ,n5112 ,n5113);
    nor g2501(n6424 ,n6213 ,n6347);
    xnor g2502(n4680 ,n4514 ,n4479);
    xnor g2503(n3077 ,n7753 ,n40[14]);
    nor g2504(n4148 ,n4012 ,n4008);
    nor g2505(n4996 ,n4967 ,n4990);
    xnor g2506(n4000 ,n37[2] ,n20[2]);
    xnor g2507(n2780 ,n2688 ,n2705);
    not g2508(n2393 ,n2392);
    not g2509(n7144 ,n7143);
    dff g2510(.RN(n1), .SN(1'b1), .CK(n0), .D(n1667), .Q(n35[2]));
    nor g2511(n6664 ,n6525 ,n6523);
    nor g2512(n3907 ,n3900 ,n3906);
    nor g2513(n6821 ,n6684 ,n6751);
    not g2514(n6151 ,n6150);
    nor g2515(n1432 ,n686 ,n638);
    not g2516(n4041 ,n4040);
    not g2517(n7156 ,n7155);
    not g2518(n3315 ,n3314);
    nor g2519(n72 ,n59 ,n71);
    nor g2520(n1451 ,n701 ,n1106);
    xnor g2521(n1097 ,n656 ,n883);
    not g2522(n5551 ,n5550);
    xnor g2523(n2167 ,n1968 ,n2086);
    nor g2524(n1144 ,n1100 ,n1043);
    xnor g2525(n6399 ,n6261 ,n6132);
    nor g2526(n2628 ,n2540 ,n2593);
    or g2527(n7649 ,n7563 ,n7560);
    xnor g2528(n7302 ,n7262 ,n7285);
    not g2529(n222 ,n221);
    xor g2530(n1886 ,n2211 ,n2113);
    nor g2531(n3276 ,n3236 ,n3264);
    nor g2532(n2098 ,n1998 ,n2067);
    nor g2533(n5299 ,n5088 ,n5094);
    nor g2534(n6989 ,n6882 ,n6920);
    nor g2535(n1506 ,n802 ,n639);
    nor g2536(n3580 ,n3545 ,n3579);
    nor g2537(n1295 ,n717 ,n640);
    dff g2538(.RN(n1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n23[1]));
    or g2539(n1632 ,n1297 ,n1233);
    nor g2540(n7668 ,n7470 ,n7484);
    xnor g2541(n6294 ,n5958 ,n5998);
    xnor g2542(n6620 ,n6410 ,n6156);
    xnor g2543(n5048 ,n5001 ,n5028);
    or g2544(n1586 ,n1250 ,n1472);
    not g2545(n6526 ,n6525);
    not g2546(n244 ,n243);
    dff g2547(.RN(n1), .SN(1'b1), .CK(n0), .D(n1593), .Q(n12[8]));
    xnor g2548(n3671 ,n7805 ,n7782);
    not g2549(n4631 ,n4630);
    nor g2550(n6954 ,n6907 ,n6867);
    nor g2551(n4802 ,n4736 ,n4733);
    xnor g2552(n7716 ,n3796 ,n3716);
    nor g2553(n5666 ,n5434 ,n5504);
    not g2554(n901 ,n10[0]);
    not g2555(n4193 ,n4192);
    not g2556(n7168 ,n7167);
    dff g2557(.RN(n1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n28[12]));
    xnor g2558(n2942 ,n2908 ,n2898);
    not g2559(n7418 ,n40[8]);
    nor g2560(n3487 ,n3438 ,n3474);
    not g2561(n200 ,n199);
    nor g2562(n1353 ,n880 ,n1103);
    not g2563(n3466 ,n3465);
    dff g2564(.RN(n1), .SN(1'b1), .CK(n0), .D(n1725), .Q(n23[7]));
    not g2565(n6522 ,n6521);
    or g2566(n1617 ,n1282 ,n1443);
    or g2567(n1655 ,n1397 ,n1555);
    not g2568(n2838 ,n2837);
    nor g2569(n5584 ,n5452 ,n5206);
    not g2570(n2956 ,n2955);
    nor g2571(n3294 ,n3119 ,n3204);
    nor g2572(n5248 ,n5101 ,n5110);
    not g2573(n178 ,n177);
    xnor g2574(n7819 ,n3793 ,n3819);
    not g2575(n4161 ,n4160);
    not g2576(n3201 ,n3200);
    nor g2577(n286 ,n179 ,n241);
    xnor g2578(n5071 ,n5052 ,n5043);
    not g2579(n2481 ,n2480);
    nor g2580(n7004 ,n6911 ,n6966);
    nor g2581(n2562 ,n2445 ,n2519);
    not g2582(n941 ,n11[14]);
    nor g2583(n4829 ,n4762 ,n4802);
    nor g2584(n6196 ,n6059 ,n6010);
    buf g2585(n13[14], n10[14]);
    or g2586(n1687 ,n1339 ,n1527);
    dff g2587(.RN(n1), .SN(1'b1), .CK(n0), .D(n1717), .Q(n31[7]));
    or g2588(n1633 ,n1299 ,n1236);
    nor g2589(n2093 ,n2001 ,n2056);
    nor g2590(n3975 ,n3962 ,n3974);
    not g2591(n6242 ,n6241);
    nor g2592(n3346 ,n3225 ,n3299);
    nor g2593(n1571 ,n682 ,n634);
    not g2594(n3021 ,n40[8]);
    nor g2595(n1172 ,n1102 ,n1031);
    xnor g2596(n2130 ,n2084 ,n2028);
    or g2597(n1693 ,n1315 ,n1458);
    nor g2598(n3886 ,n3868 ,n3865);
    nor g2599(n6676 ,n6517 ,n6516);
    xnor g2600(n1963 ,n1952 ,n1938);
    nor g2601(n3541 ,n3501 ,n3509);
    nor g2602(n5484 ,n5101 ,n5099);
    nor g2603(n1254 ,n715 ,n638);
    nor g2604(n1460 ,n734 ,n634);
    or g2605(n1784 ,n1421 ,n1142);
    nor g2606(n4078 ,n4011 ,n4007);
    or g2607(n1674 ,n1357 ,n1566);
    nor g2608(n3223 ,n3086 ,n3182);
    not g2609(n810 ,n27[0]);
    nor g2610(n6901 ,n6624 ,n6822);
    xnor g2611(n6185 ,n5792 ,n5306);
    not g2612(n742 ,n4[0]);
    or g2613(n1646 ,n1342 ,n1549);
    nor g2614(n5597 ,n5256 ,n5432);
    nor g2615(n3283 ,n3139 ,n3214);
    nor g2616(n4791 ,n4701 ,n4748);
    nor g2617(n5272 ,n5115 ,n5107);
    not g2618(n4757 ,n4756);
    xor g2619(n1881 ,n1912 ,n1929);
    xnor g2620(n41[4] ,n7136 ,n7103);
    nor g2621(n114 ,n99 ,n112);
    nor g2622(n3712 ,n3650 ,n3685);
    not g2623(n4199 ,n4198);
    not g2624(n4266 ,n4265);
    nor g2625(n6840 ,n6665 ,n6746);
    or g2626(n7681 ,n7604 ,n7672);
    nor g2627(n1494 ,n770 ,n1099);
    nor g2628(n2407 ,n2371 ,n2403);
    xnor g2629(n6440 ,n6071 ,n6185);
    not g2630(n4085 ,n4084);
    nor g2631(n2282 ,n2119 ,n2252);
    nor g2632(n3470 ,n3414 ,n3433);
    nor g2633(n1914 ,n19[4] ,n19[3]);
    nor g2634(n6216 ,n5754 ,n6036);
    nor g2635(n4324 ,n4089 ,n4197);
    xor g2636(n38[2] ,n39[2] ,n7844);
    not g2637(n4177 ,n4176);
    or g2638(n1599 ,n1262 ,n1479);
    xnor g2639(n4727 ,n4607 ,n4544);
    nor g2640(n7020 ,n6896 ,n6921);
    dff g2641(.RN(n1), .SN(1'b1), .CK(n0), .D(n1739), .Q(n30[3]));
    xnor g2642(n5835 ,n5577 ,n5299);
    or g2643(n1759 ,n1398 ,n1543);
    nor g2644(n7205 ,n7113 ,n7182);
    nor g2645(n7124 ,n7058 ,n7086);
    nor g2646(n1213 ,n654 ,n1101);
    xnor g2647(n4975 ,n4923 ,n4906);
    dff g2648(.RN(n1), .SN(1'b1), .CK(n0), .D(n1700), .Q(n33[1]));
    not g2649(n7440 ,n38[1]);
    nor g2650(n2757 ,n2696 ,n2699);
    xnor g2651(n7173 ,n7109 ,n7083);
    nor g2652(n3473 ,n3388 ,n3430);
    nor g2653(n3902 ,n3886 ,n3893);
    nor g2654(n5667 ,n5157 ,n5185);
    not g2655(n7430 ,n7805);
    nor g2656(n76 ,n58 ,n75);
    nor g2657(n5575 ,n5095 ,n5094);
    or g2658(n7484 ,n7456 ,n7480);
    xnor g2659(n479 ,n415 ,n390);
    not g2660(n2436 ,n22[2]);
    xor g2661(n6284 ,n5759 ,n5982);
    nor g2662(n5924 ,n5545 ,n5595);
    xnor g2663(n2718 ,n2511 ,n2624);
    nor g2664(n3312 ,n3209 ,n3201);
    or g2665(n198 ,n159 ,n157);
    nor g2666(n2534 ,n2441 ,n2523);
    xnor g2667(n3063 ,n40[1] ,n7740);
    xnor g2668(n4819 ,n4725 ,n4737);
    or g2669(n7703 ,n7659 ,n7653);
    nor g2670(n7470 ,n7329 ,n7335);
    nor g2671(n6825 ,n6699 ,n6761);
    nor g2672(n3576 ,n3564 ,n3575);
    nor g2673(n313 ,n236 ,n176);
    not g2674(n3250 ,n3249);
    xor g2675(n4771 ,n4681 ,n4597);
    not g2676(n4075 ,n4074);
    nor g2677(n3812 ,n3756 ,n3811);
    not g2678(n926 ,n25[5]);
    nor g2679(n1992 ,n1902 ,n1980);
    nor g2680(n7519 ,n7421 ,n7478);
    not g2681(n893 ,n1836);
    nor g2682(n1369 ,n862 ,n1107);
    nor g2683(n6319 ,n6086 ,n6076);
    not g2684(n160 ,n37[2]);
    nor g2685(n1248 ,n866 ,n640);
    nor g2686(n1933 ,n1896 ,n1914);
    xnor g2687(n566 ,n524 ,n495);
    not g2688(n7355 ,n7760);
    nor g2689(n1372 ,n913 ,n1105);
    nor g2690(n2739 ,n2718 ,n2692);
    nor g2691(n6449 ,n6188 ,n6309);
    nor g2692(n7232 ,n7158 ,n7202);
    not g2693(n101 ,n25[1]);
    nor g2694(n7600 ,n7331 ,n7481);
    nor g2695(n5086 ,n5011 ,n5085);
    not g2696(n5754 ,n5753);
    xnor g2697(n1019 ,n647 ,n873);
    nor g2698(n5047 ,n5002 ,n5029);
    nor g2699(n6761 ,n6677 ,n6655);
    not g2700(n2901 ,n2900);
    not g2701(n202 ,n201);
    not g2702(n770 ,n6[7]);
    nor g2703(n7501 ,n7386 ,n7478);
    not g2704(n5291 ,n5290);
    xnor g2705(n4591 ,n4373 ,n4158);
    nor g2706(n3931 ,n3874 ,n3930);
    nor g2707(n2195 ,n2152 ,n2138);
    nor g2708(n2019 ,n1893 ,n1982);
    nor g2709(n2050 ,n1894 ,n2004);
    nor g2710(n5330 ,n5114 ,n5098);
    xor g2711(n7753 ,n7815 ,n7792);
    not g2712(n4502 ,n4501);
    nor g2713(n2199 ,n2163 ,n2144);
    nor g2714(n6467 ,n6167 ,n6345);
    xnor g2715(n3674 ,n7808 ,n7785);
    not g2716(n377 ,n376);
    xnor g2717(n7204 ,n7138 ,n7105);
    not g2718(n6580 ,n6579);
    not g2719(n6186 ,n6185);
    xor g2720(n6393 ,n6182 ,n6122);
    nor g2721(n3299 ,n3116 ,n3219);
    nor g2722(n356 ,n183 ,n326);
    nor g2723(n7592 ,n7455 ,n7474);
    or g2724(n7699 ,n7651 ,n7650);
    nor g2725(n4160 ,n4013 ,n4019);
    not g2726(n7039 ,n7038);
    nor g2727(n1499 ,n787 ,n639);
    nor g2728(n75 ,n64 ,n74);
    nor g2729(n3225 ,n3060 ,n3168);
    nor g2730(n4963 ,n4864 ,n4931);
    nor g2731(n7461 ,n41[5] ,n7823);
    not g2732(n849 ,n20[1]);
    nor g2733(n5370 ,n5119 ,n5097);
    nor g2734(n3863 ,n3836 ,n3862);
    nor g2735(n3268 ,n3054 ,n3125);
    not g2736(n7330 ,n41[12]);
    not g2737(n5213 ,n5212);
    nor g2738(n4344 ,n4043 ,n4045);
    not g2739(n2682 ,n2681);
    nor g2740(n2207 ,n2115 ,n2173);
    xnor g2741(n4532 ,n4388 ,n4127);
    nor g2742(n4314 ,n4193 ,n4219);
    nor g2743(n2070 ,n1989 ,n2038);
    nor g2744(n1558 ,n666 ,n1106);
    xor g2745(n1844 ,n564 ,n630);
    nor g2746(n5680 ,n5431 ,n5373);
    not g2747(n122 ,n33[0]);
    nor g2748(n5535 ,n5096 ,n5106);
    nor g2749(n5232 ,n5115 ,n5119);
    nor g2750(n7584 ,n7446 ,n7474);
    nor g2751(n6213 ,n5960 ,n6042);
    xnor g2752(n6495 ,n6298 ,n6003);
    nor g2753(n1228 ,n825 ,n642);
    xnor g2754(n7718 ,n3783 ,n3799);
    nor g2755(n4146 ,n4015 ,n4008);
    xnor g2756(n4682 ,n4565 ,n4507);
    nor g2757(n4940 ,n4753 ,n4895);
    xnor g2758(n2245 ,n2079 ,n2206);
    nor g2759(n3232 ,n3113 ,n3143);
    nor g2760(n53 ,n37[7] ,n19[7]);
    not g2761(n4734 ,n4733);
    not g2762(n3708 ,n3707);
    nor g2763(n6690 ,n6429 ,n6568);
    not g2764(n3356 ,n3355);
    nor g2765(n3947 ,n7790 ,n7775);
    not g2766(n6031 ,n6030);
    nor g2767(n3451 ,n3373 ,n3409);
    nor g2768(n6764 ,n6702 ,n6621);
    xor g2769(n7767 ,n3844 ,n3860);
    nor g2770(n6731 ,n6486 ,n6691);
    nor g2771(n2816 ,n2744 ,n2791);
    dff g2772(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[1]), .Q(n15[5]));
    nor g2773(n1480 ,n788 ,n639);
    or g2774(n993 ,n17[4] ,n17[5]);
    xnor g2775(n2219 ,n2168 ,n2134);
    not g2776(n4165 ,n4164);
    xor g2777(n2427 ,n2515 ,n2636);
    nor g2778(n1179 ,n1106 ,n1079);
    nor g2779(n7122 ,n7030 ,n7084);
    not g2780(n7420 ,n7813);
    not g2781(n932 ,n10[3]);
    not g2782(n3211 ,n3210);
    nor g2783(n2603 ,n2431 ,n2548);
    nor g2784(n1416 ,n870 ,n642);
    or g2785(n994 ,n9[1] ,n9[0]);
    nor g2786(n2538 ,n2441 ,n2521);
    not g2787(n3518 ,n3517);
    nor g2788(n4123 ,n4007 ,n4010);
    nor g2789(n5328 ,n5112 ,n5117);
    not g2790(n7382 ,n40[14]);
    nor g2791(n6453 ,n6176 ,n6318);
    nor g2792(n3092 ,n3012 ,n3033);
    nor g2793(n2032 ,n1943 ,n2020);
    xnor g2794(n7163 ,n7120 ,n7040);
    xnor g2795(n2173 ,n1968 ,n2077);
    nor g2796(n7578 ,n7427 ,n7478);
    or g2797(n1740 ,n1379 ,n1191);
    nor g2798(n277 ,n147 ,n151);
    xnor g2799(n4600 ,n4366 ,n4125);
    xnor g2800(n4898 ,n4821 ,n4765);
    or g2801(n5345 ,n5088 ,n5099);
    or g2802(n1091 ,n996 ,n995);
    nor g2803(n2096 ,n2025 ,n2058);
    xnor g2804(n6720 ,n6523 ,n6525);
    not g2805(n7367 ,n38[7]);
    not g2806(n2442 ,n7766);
    not g2807(n7029 ,n7028);
    nor g2808(n4839 ,n4765 ,n4774);
    nor g2809(n1541 ,n740 ,n641);
    nor g2810(n1954 ,n1931 ,n1932);
    or g2811(n1716 ,n1434 ,n1165);
    nor g2812(n1349 ,n924 ,n636);
    xnor g2813(n4520 ,n4384 ,n4106);
    nor g2814(n4485 ,n4216 ,n4403);
    nor g2815(n1415 ,n882 ,n642);
    not g2816(n121 ,n33[6]);
    nor g2817(n3561 ,n3522 ,n3534);
    or g2818(n1727 ,n1364 ,n1185);
    nor g2819(n3642 ,n3613 ,n3622);
    nor g2820(n6882 ,n6770 ,n6818);
    not g2821(n4726 ,n4725);
    nor g2822(n2553 ,n2432 ,n2517);
    not g2823(n882 ,n28[5]);
    xnor g2824(n7254 ,n7220 ,n7177);
    nor g2825(n4597 ,n4431 ,n4454);
    nor g2826(n4135 ,n4015 ,n4020);
    nor g2827(n2581 ,n2486 ,n2573);
    nor g2828(n7123 ,n7031 ,n7083);
    or g2829(n7659 ,n7583 ,n7573);
    xnor g2830(n6519 ,n6278 ,n5964);
    xor g2831(n7764 ,n3849 ,n3854);
    nor g2832(n6575 ,n6385 ,n6465);
    not g2833(n4831 ,n4830);
    nor g2834(n3467 ,n3385 ,n3423);
    not g2835(n164 ,n163);
    nor g2836(n3966 ,n3939 ,n3965);
    or g2837(n988 ,n27[5] ,n27[6]);
    nor g2838(n2295 ,n2257 ,n2281);
    xnor g2839(n7292 ,n7255 ,n7243);
    not g2840(n867 ,n31[6]);
    not g2841(n256 ,n255);
    not g2842(n818 ,n24[6]);
    nor g2843(n2499 ,n2445 ,n2477);
    not g2844(n707 ,n11[0]);
    nor g2845(n6900 ,n6736 ,n6800);
    nor g2846(n4614 ,n4321 ,n4570);
    nor g2847(n6446 ,n6053 ,n6368);
    buf g2848(n14[2], n11[2]);
    xnor g2849(n3887 ,n7816 ,n41[15]);
    nor g2850(n7469 ,n7392 ,n7336);
    not g2851(n5429 ,n5428);
    nor g2852(n469 ,n431 ,n418);
    nor g2853(n2458 ,n21[1] ,n22[1]);
    not g2854(n159 ,n37[3]);
    not g2855(n3608 ,n7801);
    nor g2856(n1990 ,n1903 ,n1980);
    nor g2857(n5907 ,n5533 ,n5607);
    xnor g2858(n2287 ,n2213 ,n2137);
    nor g2859(n4090 ,n4029 ,n4020);
    nor g2860(n3447 ,n3317 ,n3392);
    xnor g2861(n7069 ,n7022 ,n7015);
    nor g2862(n4961 ,n4918 ,n4944);
    nor g2863(n2740 ,n2720 ,n2694);
    not g2864(n2350 ,n2349);
    xnor g2865(n3735 ,n39[4] ,n3671);
    not g2866(n1895 ,n19[5]);
    not g2867(n2448 ,n22[6]);
    nor g2868(n5454 ,n5098 ,n5106);
    nor g2869(n7320 ,n7295 ,n7319);
    xor g2870(n38[0] ,n39[0] ,n7846);
    nor g2871(n4655 ,n4494 ,n4593);
    not g2872(n6855 ,n6854);
    nor g2873(n7500 ,n7345 ,n7475);
    dff g2874(.RN(n1), .SN(1'b1), .CK(n0), .D(n1643), .Q(n10[8]));
    nor g2875(n2462 ,n2450 ,n2449);
    nor g2876(n2418 ,n2398 ,n2417);
    nor g2877(n5406 ,n5100 ,n5111);
    nor g2878(n2614 ,n2444 ,n2547);
    dff g2879(.RN(n1), .SN(1'b1), .CK(n0), .D(n1697), .Q(n33[3]));
    not g2880(n761 ,n1846);
    not g2881(n594 ,n593);
    nor g2882(n1315 ,n963 ,n637);
    not g2883(n6504 ,n6503);
    not g2884(n450 ,n449);
    not g2885(n819 ,n17[6]);
    nor g2886(n3688 ,n3630 ,n3637);
    not g2887(n4555 ,n4554);
    nor g2888(n468 ,n347 ,n402);
    or g2889(n4255 ,n4021 ,n4024);
    nor g2890(n6918 ,n6740 ,n6891);
    nor g2891(n7155 ,n7089 ,n7112);
    not g2892(n5967 ,n5966);
    xnor g2893(n3895 ,n7795 ,n7803);
    not g2894(n5987 ,n5986);
    nor g2895(n3442 ,n3411 ,n3413);
    not g2896(n4013 ,n19[2]);
    not g2897(n785 ,n1852);
    not g2898(n151 ,n19[7]);
    xnor g2899(n3781 ,n3724 ,n3709);
    nor g2900(n7058 ,n6968 ,n6995);
    xnor g2901(n6712 ,n6501 ,n6420);
    nor g2902(n2570 ,n2444 ,n2525);
    nor g2903(n2024 ,n1894 ,n1974);
    not g2904(n640 ,n639);
    nor g2905(n577 ,n537 ,n549);
    nor g2906(n376 ,n308 ,n369);
    not g2907(n5296 ,n5295);
    nor g2908(n5306 ,n5115 ,n5117);
    xnor g2909(n3330 ,n3104 ,n3241);
    nor g2910(n1115 ,n635 ,n1049);
    nor g2911(n4878 ,n4788 ,n4835);
    nor g2912(n1985 ,n1893 ,n1974);
    xor g2913(n338 ,n197 ,n251);
    nor g2914(n4811 ,n4633 ,n4759);
    xnor g2915(n6780 ,n6650 ,n6592);
    nor g2916(n1300 ,n688 ,n1103);
    or g2917(n7474 ,n26[0] ,n7325);
    not g2918(n4500 ,n4499);
    not g2919(n3591 ,n39[13]);
    not g2920(n4133 ,n4132);
    or g2921(n84 ,n25[1] ,n25[0]);
    nor g2922(n4245 ,n4013 ,n4022);
    nor g2923(n6763 ,n6703 ,n6620);
    nor g2924(n1438 ,n836 ,n638);
    not g2925(n7386 ,n40[2]);
    xnor g2926(n7289 ,n7258 ,n7241);
    xnor g2927(n3796 ,n39[1] ,n3766);
    nor g2928(n2021 ,n1894 ,n1978);
    not g2929(n7119 ,n7118);
    not g2930(n4012 ,n19[0]);
    not g2931(n156 ,n37[5]);
    xnor g2932(n339 ,n229 ,n221);
    nor g2933(n5438 ,n5097 ,n5094);
    not g2934(n506 ,n505);
    not g2935(n4197 ,n4196);
    xnor g2936(n7101 ,n6982 ,n6802);
    xnor g2937(n4934 ,n4769 ,n4892);
    not g2938(n5038 ,n5037);
    not g2939(n133 ,n132);
    not g2940(n738 ,n1851);
    nor g2941(n1962 ,n1926 ,n1947);
    nor g2942(n4427 ,n4122 ,n4276);
    not g2943(n744 ,n1857);
    nor g2944(n4285 ,n4070 ,n4062);
    not g2945(n5305 ,n5304);
    xnor g2946(n3953 ,n38[7] ,n7784);
    nor g2947(n7179 ,n7129 ,n7152);
    dff g2948(.RN(n1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n22[4]));
    nor g2949(n6450 ,n6184 ,n6312);
    nor g2950(n6813 ,n6585 ,n6759);
    nor g2951(n4651 ,n4498 ,n4556);
    xnor g2952(n6915 ,n6800 ,n6838);
    nor g2953(n5723 ,n5481 ,n5151);
    nor g2954(n1381 ,n839 ,n637);
    xnor g2955(n4858 ,n4727 ,n4789);
    nor g2956(n6361 ,n6240 ,n6120);
    nor g2957(n1409 ,n845 ,n640);
    not g2958(n6502 ,n6501);
    not g2959(n7449 ,n7731);
    or g2960(n5569 ,n5091 ,n5104);
    not g2961(n3217 ,n3216);
    nor g2962(n3450 ,n3301 ,n3408);
    nor g2963(n605 ,n578 ,n582);
    not g2964(n7443 ,n7736);
    not g2965(n6159 ,n6158);
    not g2966(n4553 ,n4552);
    nor g2967(n4576 ,n4288 ,n4512);
    not g2968(n1936 ,n1937);
    not g2969(n1971 ,n1972);
    nor g2970(n1210 ,n824 ,n1101);
    nor g2971(n6584 ,n6387 ,n6467);
    xnor g2972(n1068 ,n810 ,n842);
    nor g2973(n627 ,n607 ,n626);
    not g2974(n6145 ,n6144);
    not g2975(n4014 ,n19[5]);
    nor g2976(n4319 ,n4201 ,n4091);
    not g2977(n5237 ,n5236);
    xor g2978(n4389 ,n4120 ,n4088);
    not g2979(n7041 ,n7040);
    nor g2980(n2873 ,n2765 ,n2844);
    or g2981(n980 ,n35[8] ,n35[15]);
    not g2982(n5175 ,n5174);
    nor g2983(n4810 ,n4681 ,n4724);
    nor g2984(n5035 ,n5007 ,n5024);
    nor g2985(n2966 ,n2956 ,n2945);
    nor g2986(n292 ,n251 ,n177);
    not g2987(n6972 ,n6971);
    xnor g2988(n6785 ,n6640 ,n6638);
    not g2989(n5127 ,n5126);
    xnor g2990(n6126 ,n5849 ,n5146);
    nor g2991(n2089 ,n1986 ,n2065);
    nor g2992(n3236 ,n3112 ,n3142);
    not g2993(n4119 ,n4118);
    nor g2994(n4703 ,n4562 ,n4646);
    buf g2995(n13[2], n10[2]);
    nor g2996(n3202 ,n3048 ,n3133);
    nor g2997(n257 ,n145 ,n152);
    nor g2998(n4570 ,n4300 ,n4480);
    not g2999(n345 ,n344);
    nor g3000(n1920 ,n1898 ,n1895);
    nor g3001(n5456 ,n5118 ,n5119);
    nor g3002(n5174 ,n5118 ,n5114);
    nor g3003(n7052 ,n6967 ,n6994);
    nor g3004(n6955 ,n6796 ,n6871);
    nor g3005(n1394 ,n709 ,n1101);
    xnor g3006(n2858 ,n2502 ,n2829);
    nor g3007(n6727 ,n6505 ,n6622);
    nor g3008(n573 ,n518 ,n550);
    nor g3009(n5960 ,n5723 ,n5854);
    or g3010(n7646 ,n7557 ,n7500);
    or g3011(n1575 ,n1238 ,n1466);
    xnor g3012(n39[11] ,n2972 ,n2985);
    nor g3013(n3639 ,n39[10] ,n7788);
    or g3014(n1798 ,n1435 ,n1511);
    not g3015(n180 ,n179);
    nor g3016(n4458 ,n4329 ,n4419);
    nor g3017(n5515 ,n5096 ,n5111);
    not g3018(n4191 ,n4190);
    nor g3019(n3273 ,n3197 ,n3224);
    not g3020(n4469 ,n4468);
    nor g3021(n1163 ,n1102 ,n1066);
    nor g3022(n5220 ,n5103 ,n5106);
    xor g3023(n41[13] ,n7302 ,n7318);
    nor g3024(n2319 ,n2251 ,n2308);
    or g3025(n7705 ,n7635 ,n7634);
    nor g3026(n7579 ,n7432 ,n7476);
    nor g3027(n5745 ,n5300 ,n5578);
    nor g3028(n6557 ,n6242 ,n6426);
    not g3029(n5750 ,n5749);
    not g3030(n1906 ,n20[6]);
    xnor g3031(n6599 ,n6442 ,n6006);
    not g3032(n4407 ,n4406);
    nor g3033(n3883 ,n7807 ,n41[6]);
    not g3034(n439 ,n438);
    nor g3035(n4421 ,n4144 ,n4301);
    or g3036(n1779 ,n1416 ,n1139);
    nor g3037(n4943 ,n4885 ,n4899);
    nor g3038(n4416 ,n4263 ,n4302);
    nor g3039(n6680 ,n6177 ,n6564);
    not g3040(n6272 ,n6271);
    xnor g3041(n3901 ,n41[4] ,n7805);
    nor g3042(n1486 ,n759 ,n639);
    nor g3043(n1527 ,n736 ,n641);
    xnor g3044(n6934 ,n6784 ,n6836);
    nor g3045(n3444 ,n3382 ,n3380);
    buf g3046(n15[3], 1'b0);
    not g3047(n6135 ,n6134);
    nor g3048(n4764 ,n4649 ,n4694);
    nor g3049(n2594 ,n2433 ,n2549);
    nor g3050(n6885 ,n6672 ,n6819);
    not g3051(n862 ,n31[1]);
    not g3052(n853 ,n34[10]);
    nor g3053(n2546 ,n2433 ,n2523);
    not g3054(n7403 ,n7722);
    or g3055(n999 ,n808 ,n644);
    not g3056(n3599 ,n39[1]);
    not g3057(n806 ,n1869);
    xnor g3058(n4777 ,n4676 ,n4602);
    not g3059(n635 ,n636);
    nor g3060(n5496 ,n5112 ,n5110);
    nor g3061(n3928 ,n3896 ,n3927);
    or g3062(n1704 ,n1351 ,n1159);
    nor g3063(n7596 ,n7355 ,n7479);
    nor g3064(n4488 ,n4359 ,n4405);
    nor g3065(n7313 ,n7312 ,n7307);
    or g3066(n1703 ,n1215 ,n1532);
    or g3067(n7689 ,n7502 ,n7666);
    nor g3068(n5902 ,n5561 ,n5645);
    not g3069(n174 ,n173);
    nor g3070(n4642 ,n4468 ,n4545);
    or g3071(n1610 ,n1274 ,n1485);
    nor g3072(n2333 ,n2226 ,n2295);
    nor g3073(n3970 ,n3964 ,n3969);
    dff g3074(.RN(n1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n28[5]));
    xnor g3075(n2725 ,n2511 ,n2629);
    nor g3076(n3476 ,n3394 ,n3426);
    nor g3077(n6667 ,n6389 ,n6533);
    nor g3078(n3493 ,n3464 ,n3465);
    xnor g3079(n6291 ,n5995 ,n6032);
    nor g3080(n3249 ,n3087 ,n3183);
    xor g3081(n5763 ,n5347 ,n5396);
    nor g3082(n6756 ,n6577 ,n6627);
    xor g3083(n5799 ,n5555 ,n5390);
    or g3084(n7692 ,n7639 ,n7636);
    nor g3085(n132 ,n127 ,n130);
    nor g3086(n4879 ,n4756 ,n4830);
    not g3087(n4899 ,n4898);
    nor g3088(n6920 ,n6790 ,n6860);
    or g3089(n1780 ,n1226 ,n1197);
    nor g3090(n3973 ,n3961 ,n3972);
    xnor g3091(n3324 ,n3118 ,n3204);
    nor g3092(n3255 ,n3052 ,n3135);
    nor g3093(n4475 ,n4314 ,n4422);
    nor g3094(n2056 ,n1893 ,n2004);
    not g3095(n6127 ,n6126);
    not g3096(n7441 ,n7718);
    not g3097(n6131 ,n6130);
    xnor g3098(n1025 ,n870 ,n835);
    nor g3099(n448 ,n381 ,n427);
    not g3100(n4006 ,n37[3]);
    nor g3101(n6444 ,n6273 ,n6354);
    nor g3102(n173 ,n156 ,n158);
    nor g3103(n3047 ,n2994 ,n3030);
    not g3104(n4022 ,n37[7]);
    nor g3105(n591 ,n559 ,n570);
    or g3106(n1982 ,n1936 ,n1964);
    not g3107(n6939 ,n6938);
    nor g3108(n3286 ,n3110 ,n3211);
    or g3109(n7674 ,n7641 ,n7623);
    xor g3110(n5769 ,n5562 ,n5430);
    xnor g3111(n4902 ,n4817 ,n4721);
    xnor g3112(n2833 ,n2772 ,n2733);
    nor g3113(n6555 ,n6098 ,n6419);
    not g3114(n5263 ,n5262);
    not g3115(n147 ,n37[4]);
    not g3116(n7332 ,n41[14]);
    nor g3117(n4707 ,n4575 ,n4638);
    xnor g3118(n2837 ,n2777 ,n2653);
    dff g3119(.RN(n1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n27[5]));
    nor g3120(n5152 ,n5112 ,n5099);
    not g3121(n4115 ,n4114);
    not g3122(n2208 ,n2207);
    xnor g3123(n2779 ,n2667 ,n2427);
    or g3124(n1686 ,n1338 ,n1525);
    xnor g3125(n6717 ,n6537 ,n6591);
    xnor g3126(n6299 ,n5997 ,n5940);
    not g3127(n668 ,n22[4]);
    not g3128(n2997 ,n7744);
    nor g3129(n3940 ,n7786 ,n7771);
    xnor g3130(n4860 ,n4791 ,n4756);
    nor g3131(n298 ,n168 ,n164);
    nor g3132(n3543 ,n3490 ,n3506);
    nor g3133(n3817 ,n3777 ,n3816);
    not g3134(n99 ,n25[4]);
    xnor g3135(n2339 ,n2215 ,n2304);
    nor g3136(n3044 ,n2994 ,n3031);
    nor g3137(n4497 ,n4323 ,n4442);
    nor g3138(n1553 ,n900 ,n1100);
    not g3139(n2659 ,n2658);
    xnor g3140(n4542 ,n4370 ,n4121);
    nor g3141(n4096 ,n4006 ,n4016);
    or g3142(n3032 ,n3010 ,n3006);
    not g3143(n5941 ,n5940);
    nor g3144(n5172 ,n5114 ,n5116);
    nor g3145(n4036 ,n4027 ,n4008);
    nor g3146(n1989 ,n1903 ,n1976);
    xor g3147(n5779 ,n5548 ,n5138);
    nor g3148(n1961 ,n1927 ,n1949);
    xnor g3149(n3344 ,n3114 ,n3224);
    xnor g3150(n2149 ,n2092 ,n1970);
    nor g3151(n5950 ,n5676 ,n5861);
    not g3152(n581 ,n580);
    nor g3153(n2598 ,n2445 ,n2548);
    xnor g3154(n4408 ,n4249 ,n4148);
    dff g3155(.RN(n1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n34[15]));
    nor g3156(n4806 ,n4665 ,n4742);
    not g3157(n90 ,n33[5]);
    not g3158(n5742 ,n5741);
    xnor g3159(n7149 ,n7066 ,n6973);
    nor g3160(n2328 ,n2306 ,n2302);
    xnor g3161(n1938 ,n20[3] ,n19[3]);
    not g3162(n3933 ,n7778);
    nor g3163(n3187 ,n3013 ,n3075);
    nor g3164(n1302 ,n692 ,n1101);
    nor g3165(n2265 ,n2184 ,n2230);
    nor g3166(n3108 ,n3013 ,n3041);
    not g3167(n7225 ,n7224);
    nor g3168(n7273 ,n7246 ,n7270);
    nor g3169(n3658 ,n3600 ,n3625);
    nor g3170(n2232 ,n2172 ,n2193);
    not g3171(n7340 ,n7780);
    xnor g3172(n2727 ,n2511 ,n2642);
    xnor g3173(n440 ,n347 ,n382);
    xnor g3174(n3894 ,n7800 ,n7812);
    nor g3175(n3122 ,n3013 ,n3040);
    nor g3176(n1186 ,n1006 ,n1104);
    nor g3177(n3562 ,n3518 ,n3538);
    not g3178(n5401 ,n5400);
    nor g3179(n6579 ,n6356 ,n6445);
    not g3180(n155 ,n19[4]);
    not g3181(n5981 ,n5980);
    not g3182(n2148 ,n2147);
    xnor g3183(n1966 ,n1953 ,n1928);
    nor g3184(n5356 ,n5116 ,n5113);
    nor g3185(n632 ,n548 ,n631);
    nor g3186(n4847 ,n4730 ,n4781);
    not g3187(n4883 ,n4882);
    or g3188(n1736 ,n1220 ,n1151);
    nor g3189(n4747 ,n4710 ,n4627);
    not g3190(n7158 ,n7157);
    not g3191(n756 ,n3[1]);
    not g3192(n3380 ,n3379);
    nor g3193(n285 ,n219 ,n281);
    nor g3194(n4945 ,n4872 ,n4902);
    dff g3195(.RN(n1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n18[1]));
    nor g3196(n7047 ,n6917 ,n7001);
    xnor g3197(n2516 ,n2454 ,n2504);
    xnor g3198(n7799 ,n7308 ,n7312);
    nor g3199(n3697 ,n3659 ,n3692);
    nor g3200(n6823 ,n6664 ,n6747);
    nor g3201(n7265 ,n7253 ,n7228);
    nor g3202(n2351 ,n2262 ,n2324);
    nor g3203(n631 ,n562 ,n630);
    or g3204(n7628 ,n7558 ,n7508);
    nor g3205(n2307 ,n2185 ,n2288);
    not g3206(n3161 ,n3160);
    or g3207(n7691 ,n7638 ,n7637);
    dff g3208(.RN(n1), .SN(1'b1), .CK(n0), .D(n1585), .Q(n12[12]));
    or g3209(n1095 ,n978 ,n988);
    nor g3210(n2646 ,n2530 ,n2585);
    nor g3211(n4242 ,n4022 ,n4026);
    not g3212(n2632 ,n2631);
    nor g3213(n1329 ,n832 ,n637);
    not g3214(n5109 ,n19[5]);
    nor g3215(n1880 ,n105 ,n104);
    xnor g3216(n6845 ,n6642 ,n6776);
    nor g3217(n2391 ,n2305 ,n2370);
    not g3218(n2695 ,n2694);
    or g3219(n4269 ,n4021 ,n4026);
    nor g3220(n6056 ,n5732 ,n5911);
    xnor g3221(n5050 ,n5014 ,n5003);
    nor g3222(n5494 ,n5096 ,n5105);
    not g3223(n5507 ,n5506);
    nor g3224(n2005 ,n1958 ,n1981);
    nor g3225(n5270 ,n5090 ,n5113);
    nor g3226(n1910 ,n19[3] ,n20[3]);
    nor g3227(n5124 ,n5119 ,n5098);
    not g3228(n6701 ,n6700);
    xnor g3229(n6525 ,n6282 ,n6063);
    nor g3230(n1948 ,n1919 ,n1935);
    not g3231(n889 ,n24[8]);
    nor g3232(n3663 ,n3608 ,n3631);
    nor g3233(n4294 ,n4042 ,n4044);
    or g3234(n992 ,n23[4] ,n23[5]);
    xnor g3235(n1924 ,n1906 ,n20[5]);
    nor g3236(n3835 ,n37[7] ,n19[7]);
    xor g3237(n7734 ,n3568 ,n3581);
    nor g3238(n1309 ,n697 ,n642);
    xnor g3239(n2923 ,n2889 ,n2782);
    nor g3240(n1133 ,n641 ,n1057);
    dff g3241(.RN(n1), .SN(1'b1), .CK(n0), .D(n1618), .Q(n1835));
    nor g3242(n2025 ,n1890 ,n1980);
    xnor g3243(n7136 ,n7079 ,n6971);
    nor g3244(n3799 ,n3757 ,n3798);
    nor g3245(n5589 ,n5238 ,n5404);
    nor g3246(n3838 ,n3831 ,n3832);
    nor g3247(n7511 ,n7389 ,n7479);
    nor g3248(n3177 ,n2995 ,n3073);
    nor g3249(n6456 ,n6162 ,n6341);
    nor g3250(n4251 ,n4015 ,n4019);
    nor g3251(n7096 ,n6998 ,n7034);
    nor g3252(n4645 ,n4504 ,n4536);
    not g3253(n3002 ,n7743);
    xnor g3254(n2903 ,n2870 ,n2788);
    nor g3255(n2042 ,n1893 ,n2002);
    nor g3256(n4150 ,n4012 ,n4018);
    nor g3257(n2624 ,n2536 ,n2590);
    nor g3258(n5210 ,n5118 ,n5102);
    nor g3259(n5691 ,n5223 ,n5275);
    not g3260(n5961 ,n5960);
    nor g3261(n7590 ,n7448 ,n7475);
    nor g3262(n457 ,n387 ,n428);
    nor g3263(n6064 ,n5701 ,n5891);
    not g3264(n228 ,n227);
    xnor g3265(n4772 ,n4632 ,n4712);
    not g3266(n4045 ,n4044);
    or g3267(n7708 ,n7619 ,n7675);
    nor g3268(n7669 ,n7469 ,n7486);
    nor g3269(n1297 ,n902 ,n637);
    nor g3270(n7011 ,n6879 ,n6928);
    nor g3271(n6769 ,n6576 ,n6615);
    nor g3272(n5060 ,n4999 ,n5042);
    not g3273(n4155 ,n4154);
    not g3274(n2439 ,n22[0]);
    nor g3275(n2378 ,n2334 ,n2355);
    nor g3276(n3716 ,n3610 ,n3679);
    dff g3277(.RN(n1), .SN(1'b1), .CK(n0), .D(n1642), .Q(n10[9]));
    xnor g3278(n507 ,n441 ,n376);
    not g3279(n5351 ,n5350);
    nor g3280(n2312 ,n2264 ,n2286);
    nor g3281(n6971 ,n6750 ,n6887);
    not g3282(n643 ,n18[2]);
    nor g3283(n5420 ,n5093 ,n5110);
    nor g3284(n4060 ,n4023 ,n4019);
    nor g3285(n5010 ,n4927 ,n4979);
    or g3286(n7465 ,n26[2] ,n26[1]);
    nor g3287(n5995 ,n5733 ,n5884);
    xnor g3288(n41[6] ,n7238 ,n7234);
    not g3289(n3605 ,n39[2]);
    xnor g3290(n1037 ,n888 ,n852);
    nor g3291(n6776 ,n6559 ,n6662);
    xnor g3292(n4956 ,n4898 ,n4884);
    or g3293(n1786 ,n1424 ,n1133);
    nor g3294(n7491 ,n7366 ,n7477);
    nor g3295(n6336 ,n6090 ,n6259);
    nor g3296(n55 ,n37[0] ,n19[0]);
    nor g3297(n2092 ,n2012 ,n2054);
    not g3298(n7170 ,n7169);
    nor g3299(n2035 ,n1956 ,n2019);
    xnor g3300(n4871 ,n4768 ,n4713);
    xnor g3301(n1859 ,n61 ,n81);
    xnor g3302(n3328 ,n3237 ,n3253);
    nor g3303(n4479 ,n4345 ,n4439);
    nor g3304(n4865 ,n4800 ,n4824);
    nor g3305(n2764 ,n2654 ,n2686);
    not g3306(n836 ,n20[5]);
    not g3307(n5105 ,n19[7]);
    xnor g3308(n3327 ,n3138 ,n3214);
    xor g3309(n5767 ,n5534 ,n5128);
    not g3310(n4053 ,n4052);
    nor g3311(n3127 ,n3012 ,n3077);
    nor g3312(n2259 ,n2206 ,n2229);
    not g3313(n6155 ,n6154);
    xnor g3314(n7071 ,n6983 ,n6943);
    not g3315(n7379 ,n7772);
    xnor g3316(n7087 ,n6977 ,n6942);
    nor g3317(n5224 ,n5090 ,n5110);
    xnor g3318(n1088 ,n24[0] ,n35[0]);
    nor g3319(n5663 ,n5253 ,n5393);
    not g3320(n2667 ,n2666);
    not g3321(n5169 ,n5168);
    or g3322(n1783 ,n1422 ,n1505);
    xnor g3323(n1070 ,n24[6] ,n35[6]);
    or g3324(n1753 ,n1224 ,n1195);
    or g3325(n7673 ,n7582 ,n7579);
    xnor g3326(n3377 ,n3337 ,n3239);
    not g3327(n3603 ,n7804);
    nor g3328(n1235 ,n656 ,n634);
    nor g3329(n1237 ,n693 ,n638);
    nor g3330(n4448 ,n4129 ,n4293);
    nor g3331(n6309 ,n6108 ,n6106);
    nor g3332(n287 ,n253 ,n227);
    or g3333(n2477 ,n2463 ,n2457);
    or g3334(n1702 ,n1300 ,n1557);
    not g3335(n718 ,n24[14]);
    or g3336(n1661 ,n1213 ,n1158);
    nor g3337(n1273 ,n896 ,n636);
    not g3338(n920 ,n10[12]);
    nor g3339(n3925 ,n3877 ,n3924);
    xor g3340(n5816 ,n5312 ,n5484);
    not g3341(n4151 ,n4150);
    not g3342(n5385 ,n5384);
    or g3343(n1715 ,n1219 ,n1537);
    nor g3344(n7249 ,n7222 ,n7168);
    nor g3345(n7560 ,n7451 ,n7477);
    nor g3346(n318 ,n252 ,n178);
    dff g3347(.RN(n1), .SN(1'b1), .CK(n0), .D(n1615), .Q(n16[0]));
    nor g3348(n2496 ,n2470 ,n2466);
    nor g3349(n2895 ,n2864 ,n2842);
    not g3350(n4778 ,n4777);
    nor g3351(n5664 ,n5451 ,n5271);
    not g3352(n2128 ,n2127);
    xnor g3353(n5792 ,n5500 ,n5442);
    nor g3354(n5042 ,n5010 ,n5032);
    not g3355(n4101 ,n4100);
    not g3356(n2138 ,n2137);
    nor g3357(n5713 ,n5209 ,n5427);
    nor g3358(n7282 ,n7258 ,n7242);
    not g3359(n2811 ,n2810);
    nor g3360(n6842 ,n6681 ,n6744);
    nor g3361(n6014 ,n5758 ,n5837);
    or g3362(n1573 ,n1319 ,n1128);
    not g3363(n1106 ,n1107);
    nor g3364(n1993 ,n1903 ,n1978);
    nor g3365(n7151 ,n7103 ,n7125);
    nor g3366(n5040 ,n5009 ,n5025);
    not g3367(n6568 ,n6567);
    xnor g3368(n39[12] ,n2977 ,n2987);
    nor g3369(n1157 ,n1100 ,n1088);
    nor g3370(n5563 ,n5118 ,n5106);
    nor g3371(n2052 ,n1902 ,n2004);
    nor g3372(n6220 ,n5941 ,n5945);
    nor g3373(n5887 ,n5568 ,n5584);
    xnor g3374(n6529 ,n6296 ,n6116);
    not g3375(n7098 ,n7097);
    or g3376(n1012 ,n681 ,n709);
    xnor g3377(n2340 ,n2303 ,n2226);
    xnor g3378(n1052 ,n660 ,n851);
    xnor g3379(n6092 ,n5797 ,n5490);
    not g3380(n6797 ,n6796);
    dff g3381(.RN(n1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n29[0]));
    not g3382(n6649 ,n6648);
    not g3383(n139 ,n138);
    xnor g3384(n3425 ,n3322 ,n3374);
    nor g3385(n3409 ,n3315 ,n3372);
    nor g3386(n1111 ,n635 ,n1021);
    nor g3387(n5278 ,n5088 ,n5117);
    xnor g3388(n1057 ,n868 ,n825);
    not g3389(n109 ,n108);
    xnor g3390(n4981 ,n4920 ,n4938);
    nor g3391(n6894 ,n6735 ,n6801);
    not g3392(n3832 ,n19[3]);
    not g3393(n274 ,n273);
    or g3394(n1745 ,n1384 ,n1150);
    nor g3395(n613 ,n586 ,n601);
    not g3396(n2445 ,n7769);
    nor g3397(n5148 ,n5103 ,n5104);
    nor g3398(n2808 ,n2805 ,n2761);
    or g3399(n1004 ,n820 ,n824);
    xnor g3400(n6136 ,n5788 ,n5292);
    not g3401(n5307 ,n5306);
    not g3402(n6033 ,n6032);
    not g3403(n7338 ,n40[6]);
    nor g3404(n7529 ,n7390 ,n7476);
    not g3405(n7436 ,n7770);
    dff g3406(.RN(n1), .SN(1'b1), .CK(n0), .D(n1685), .Q(n34[3]));
    not g3407(n4241 ,n4240);
    not g3408(n3392 ,n3391);
    nor g3409(n1270 ,n720 ,n638);
    nor g3410(n4420 ,n4253 ,n4296);
    nor g3411(n1167 ,n1102 ,n1041);
    not g3412(n7452 ,n7812);
    dff g3413(.RN(n1), .SN(1'b1), .CK(n0), .D(n1631), .Q(n11[4]));
    nor g3414(n1448 ,n854 ,n634);
    or g3415(n991 ,n17[6] ,n17[7]);
    xnor g3416(n6975 ,n6872 ,n6825);
    xnor g3417(n1845 ,n597 ,n628);
    xnor g3418(n39[5] ,n2882 ,n2922);
    xnor g3419(n6985 ,n6790 ,n6882);
    nor g3420(n5725 ,n5507 ,n5139);
    nor g3421(n4464 ,n4335 ,n4434);
    not g3422(n7275 ,n7274);
    not g3423(n3149 ,n3148);
    xnor g3424(n5054 ,n5015 ,n4991);
    xor g3425(n7754 ,n7816 ,n7760);
    nor g3426(n7017 ,n6902 ,n6947);
    not g3427(n4081 ,n4080);
    xnor g3428(n6297 ,n6062 ,n5954);
    not g3429(n7329 ,n41[13]);
    not g3430(n5836 ,n5835);
    nor g3431(n3146 ,n2994 ,n3070);
    nor g3432(n1401 ,n834 ,n638);
    nor g3433(n6241 ,n5928 ,n6007);
    nor g3434(n203 ,n150 ,n153);
    nor g3435(n3298 ,n3164 ,n3269);
    nor g3436(n3950 ,n3933 ,n3934);
    or g3437(n1776 ,n1415 ,n1138);
    nor g3438(n6018 ,n5734 ,n5910);
    xnor g3439(n3786 ,n3747 ,n3718);
    xnor g3440(n6710 ,n6521 ,n6473);
    nor g3441(n3259 ,n3096 ,n3131);
    nor g3442(n2582 ,n2489 ,n2560);
    nor g3443(n5236 ,n5118 ,n5092);
    xnor g3444(n2303 ,n2245 ,n2190);
    nor g3445(n2237 ,n2171 ,n2182);
    not g3446(n484 ,n483);
    not g3447(n3244 ,n3243);
    not g3448(n6995 ,n6994);
    nor g3449(n1387 ,n829 ,n1103);
    xor g3450(n5808 ,n5294 ,n5282);
    not g3451(n3510 ,n3509);
    nor g3452(n1124 ,n635 ,n1055);
    nor g3453(n4656 ,n4493 ,n4594);
    not g3454(n184 ,n183);
    xnor g3455(n407 ,n336 ,n205);
    nor g3456(n5863 ,n5327 ,n5622);
    not g3457(n6863 ,n6862);
    not g3458(n4225 ,n4224);
    not g3459(n6147 ,n6146);
    not g3460(n695 ,n10[5]);
    xnor g3461(n1077 ,n645 ,n671);
    xnor g3462(n7145 ,n7068 ,n7017);
    not g3463(n4229 ,n4228);
    nor g3464(n3081 ,n2995 ,n3040);
    or g3465(n91 ,n33[4] ,n33[3]);
    nor g3466(n3872 ,n7808 ,n41[7]);
    dff g3467(.RN(n1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n28[2]));
    xnor g3468(n6644 ,n6411 ,n6096);
    or g3469(n3030 ,n3021 ,n3026);
    nor g3470(n1202 ,n645 ,n1107);
    not g3471(n2325 ,n2324);
    nor g3472(n7135 ,n7049 ,n7094);
    nor g3473(n4840 ,n4804 ,n4792);
    xnor g3474(n7829 ,n3960 ,n3982);
    not g3475(n2126 ,n2125);
    nor g3476(n1951 ,n1892 ,n1937);
    nor g3477(n614 ,n594 ,n602);
    nor g3478(n2284 ,n2176 ,n2265);
    nor g3479(n95 ,n90 ,n94);
    or g3480(n7627 ,n7570 ,n7526);
    nor g3481(n3128 ,n3012 ,n3075);
    nor g3482(n4578 ,n4312 ,n4467);
    not g3483(n6999 ,n6998);
    not g3484(n966 ,n30[5]);
    nor g3485(n2595 ,n2432 ,n2548);
    not g3486(n4533 ,n4532);
    dff g3487(.RN(n1), .SN(1'b1), .CK(n0), .D(n1727), .Q(n17[7]));
    nor g3488(n1279 ,n893 ,n638);
    or g3489(n1724 ,n1366 ,n1175);
    nor g3490(n1393 ,n844 ,n1103);
    nor g3491(n5056 ,n5037 ,n5030);
    not g3492(n4887 ,n4886);
    nor g3493(n1143 ,n1100 ,n1028);
    not g3494(n204 ,n203);
    not g3495(n3262 ,n3261);
    nor g3496(n2308 ,n2187 ,n2276);
    not g3497(n4903 ,n4902);
    not g3498(n3606 ,n7791);
    buf g3499(n37[5] ,n1836);
    xnor g3500(n3389 ,n3336 ,n3357);
    xnor g3501(n4404 ,n4251 ,n4247);
    nor g3502(n1269 ,n898 ,n636);
    nor g3503(n314 ,n246 ,n174);
    nor g3504(n1396 ,n724 ,n642);
    nor g3505(n2950 ,n2912 ,n2928);
    not g3506(n4117 ,n4116);
    nor g3507(n509 ,n461 ,n487);
    xnor g3508(n5817 ,n5266 ,n5162);
    dff g3509(.RN(n1), .SN(1'b1), .CK(n0), .D(n1743), .Q(n23[3]));
    nor g3510(n2677 ,n2511 ,n2635);
    nor g3511(n6682 ,n6504 ,n6573);
    not g3512(n6476 ,n6475);
    not g3513(n2431 ,n7762);
    nor g3514(n6758 ,n6477 ,n6631);
    nor g3515(n7183 ,n7127 ,n7149);
    not g3516(n5245 ,n5244);
    not g3517(n726 ,n5[0]);
    nor g3518(n3802 ,n3765 ,n3801);
    nor g3519(n2989 ,n2988 ,n2974);
    nor g3520(n2550 ,n2501 ,n2524);
    or g3521(n1596 ,n1258 ,n1477);
    nor g3522(n6000 ,n5711 ,n5908);
    nor g3523(n1367 ,n871 ,n1107);
    not g3524(n5969 ,n5968);
    nor g3525(n2204 ,n2124 ,n2155);
    not g3526(n968 ,n11[9]);
    nor g3527(n3237 ,n3056 ,n3169);
    xnor g3528(n5825 ,n5426 ,n5208);
    xnor g3529(n5815 ,n5436 ,n5446);
    nor g3530(n1809 ,n985 ,n1181);
    nor g3531(n6350 ,n5759 ,n6229);
    nor g3532(n4851 ,n4732 ,n4778);
    not g3533(n5251 ,n5250);
    or g3534(n5552 ,n5093 ,n5106);
    not g3535(n913 ,n30[7]);
    nor g3536(n2767 ,n2683 ,n2714);
    nor g3537(n3691 ,n3609 ,n3648);
    not g3538(n130 ,n129);
    nor g3539(n2063 ,n1890 ,n2027);
    xnor g3540(n4932 ,n4856 ,n4793);
    nor g3541(n3243 ,n3101 ,n3179);
    nor g3542(n1436 ,n945 ,n1101);
    or g3543(n1601 ,n1263 ,n1116);
    nor g3544(n5057 ,n5038 ,n5031);
    nor g3545(n1226 ,n651 ,n1105);
    or g3546(n1677 ,n1352 ,n1569);
    dff g3547(.RN(n1), .SN(1'b1), .CK(n0), .D(n1760), .Q(n22[6]));
    xnor g3548(n2910 ,n2858 ,n2801);
    not g3549(n6252 ,n6251);
    xnor g3550(n349 ,n261 ,n199);
    nor g3551(n6897 ,n6633 ,n6794);
    nor g3552(n2067 ,n1903 ,n2027);
    xnor g3553(n6790 ,n6595 ,n6469);
    nor g3554(n2600 ,n2445 ,n2547);
    not g3555(n6510 ,n6509);
    xnor g3556(n5819 ,n5416 ,n5456);
    nor g3557(n1282 ,n958 ,n637);
    not g3558(n5137 ,n5136);
    nor g3559(n5228 ,n5097 ,n5111);
    not g3560(n5163 ,n5162);
    dff g3561(.RN(n1), .SN(1'b1), .CK(n0), .D(n1735), .Q(n30[5]));
    dff g3562(.RN(n1), .SN(1'b1), .CK(n0), .D(n1658), .Q(n35[7]));
    not g3563(n2443 ,n7761);
    nor g3564(n6673 ,n6329 ,n6511);
    not g3565(n5423 ,n5422);
    nor g3566(n6909 ,n6772 ,n6812);
    nor g3567(n288 ,n243 ,n237);
    nor g3568(n6838 ,n6663 ,n6728);
    xnor g3569(n3359 ,n3270 ,n3231);
    not g3570(n3500 ,n3499);
    or g3571(n1009 ,n863 ,n948);
    nor g3572(n5875 ,n5542 ,n5658);
    not g3573(n6742 ,n6741);
    nor g3574(n2241 ,n2121 ,n2183);
    not g3575(n504 ,n503);
    or g3576(n1648 ,n1302 ,n1550);
    nor g3577(n4744 ,n4643 ,n4678);
    nor g3578(n6369 ,n6018 ,n6117);
    nor g3579(n81 ,n54 ,n80);
    nor g3580(n1164 ,n1102 ,n1067);
    not g3581(n6109 ,n6108);
    nor g3582(n7562 ,n7416 ,n7481);
    nor g3583(n7591 ,n7344 ,n7478);
    not g3584(n655 ,n36[7]);
    xnor g3585(n401 ,n338 ,n177);
    nor g3586(n3443 ,n3351 ,n3418);
    xor g3587(n5800 ,n5547 ,n5132);
    nor g3588(n3855 ,n3849 ,n3854);
    xnor g3589(n2188 ,n2122 ,n2103);
    or g3590(n1697 ,n1347 ,n1461);
    not g3591(n6828 ,n6827);
    or g3592(n7611 ,n7490 ,n7608);
    xnor g3593(n4388 ,n4068 ,n4166);
    not g3594(n6655 ,n6654);
    nor g3595(n308 ,n162 ,n196);
    nor g3596(n1192 ,n1001 ,n1104);
    not g3597(n6174 ,n6173);
    xnor g3598(n411 ,n354 ,n249);
    nor g3599(n3405 ,n3289 ,n3367);
    nor g3600(n3090 ,n2995 ,n3036);
    dff g3601(.RN(n1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n28[0]));
    not g3602(n2949 ,n2948);
    xnor g3603(n342 ,n195 ,n161);
    not g3604(n2551 ,n2550);
    nor g3605(n4444 ,n4126 ,n4281);
    not g3606(n4870 ,n4869);
    nor g3607(n2675 ,n2502 ,n2656);
    nor g3608(n3850 ,n3839 ,n3845);
    not g3609(n404 ,n403);
    xnor g3610(n2859 ,n2810 ,n2815);
    nor g3611(n4158 ,n4007 ,n4017);
    not g3612(n4401 ,n4400);
    xnor g3613(n2662 ,n2501 ,n2577);
    xor g3614(n40[4] ,n39[5] ,n7835);
    nor g3615(n5709 ,n5133 ,n5483);
    not g3616(n827 ,n24[0]);
    xnor g3617(n4383 ,n4100 ,n4078);
    nor g3618(n6353 ,n6039 ,n6243);
    nor g3619(n5731 ,n5443 ,n5501);
    not g3620(n6141 ,n6140);
    nor g3621(n6339 ,n6052 ,n6219);
    xnor g3622(n6102 ,n5791 ,n5240);
    buf g3623(n13[15], n10[15]);
    nor g3624(n5862 ,n5527 ,n5589);
    not g3625(n6085 ,n6084);
    nor g3626(n1399 ,n843 ,n638);
    xnor g3627(n5775 ,n5360 ,n5400);
    xnor g3628(n3423 ,n3326 ,n3375);
    nor g3629(n5565 ,n5100 ,n5106);
    not g3630(n5259 ,n5258);
    xnor g3631(n2946 ,n2902 ,n2910);
    nor g3632(n3449 ,n3308 ,n3407);
    nor g3633(n165 ,n160 ,n158);
    nor g3634(n2588 ,n2433 ,n2548);
    nor g3635(n4693 ,n4483 ,n4645);
    not g3636(n1892 ,n37[0]);
    nor g3637(n604 ,n595 ,n580);
    not g3638(n2828 ,n2827);
    nor g3639(n6744 ,n6587 ,n6679);
    dff g3640(.RN(n1), .SN(1'b1), .CK(n0), .D(n1654), .Q(n35[10]));
    nor g3641(n1497 ,n741 ,n639);
    not g3642(n5197 ,n5196);
    nor g3643(n5990 ,n5677 ,n5874);
    xor g3644(n1862 ,n64 ,n74);
    not g3645(n4557 ,n4556);
    nor g3646(n2937 ,n2898 ,n2909);
    nor g3647(n3998 ,n3994 ,n3993);
    nor g3648(n2590 ,n2431 ,n2547);
    nor g3649(n3556 ,n3519 ,n3535);
    nor g3650(n7553 ,n7356 ,n7475);
    xnor g3651(n4589 ,n4389 ,n4196);
    xnor g3652(n39[6] ,n2924 ,n2957);
    not g3653(n7358 ,n39[15]);
    not g3654(n746 ,n3[7]);
    not g3655(n5221 ,n5220);
    xor g3656(n7741 ,n7803 ,n7780);
    not g3657(n152 ,n19[0]);
    or g3658(n1664 ,n1210 ,n1145);
    nor g3659(n3882 ,n7809 ,n7797);
    or g3660(n1706 ,n1261 ,n1160);
    xnor g3661(n2217 ,n2149 ,n2146);
    xnor g3662(n1090 ,n656 ,n837);
    not g3663(n5357 ,n5356);
    nor g3664(n3311 ,n3254 ,n3238);
    nor g3665(n2737 ,n2674 ,n2728);
    nor g3666(n5687 ,n5261 ,n5411);
    nor g3667(n1428 ,n874 ,n638);
    not g3668(n6248 ,n6247);
    xnor g3669(n6408 ,n6094 ,n6245);
    not g3670(n196 ,n195);
    nor g3671(n2862 ,n2823 ,n2852);
    xnor g3672(n4725 ,n4606 ,n4520);
    xnor g3673(n6593 ,n6249 ,n6484);
    nor g3674(n6428 ,n6191 ,n6313);
    nor g3675(n6767 ,n6538 ,n6612);
    not g3676(n6123 ,n6122);
    not g3677(n4732 ,n4731);
    nor g3678(n1350 ,n889 ,n642);
    nor g3679(n1147 ,n1100 ,n1074);
    xnor g3680(n6622 ,n6396 ,n6178);
    xnor g3681(n6716 ,n6590 ,n6479);
    nor g3682(n3438 ,n3290 ,n3405);
    not g3683(n741 ,n6[4]);
    not g3684(n3613 ,n39[12]);
    nor g3685(n3692 ,n3629 ,n3641);
    not g3686(n6045 ,n6044);
    nor g3687(n5678 ,n5371 ,n5169);
    xnor g3688(n4556 ,n4375 ,n4112);
    xnor g3689(n6267 ,n5819 ,n5313);
    or g3690(n989 ,n23[6] ,n23[7]);
    not g3691(n7401 ,n7734);
    nor g3692(n2331 ,n2300 ,n2277);
    nor g3693(n7007 ,n6910 ,n6958);
    nor g3694(n7021 ,n6899 ,n6926);
    nor g3695(n2898 ,n2850 ,n2871);
    not g3696(n6049 ,n6048);
    nor g3697(n2352 ,n2336 ,n2327);
    not g3698(n757 ,n8[2]);
    not g3699(n5469 ,n5468);
    nor g3700(n3134 ,n3012 ,n3076);
    nor g3701(n2566 ,n2444 ,n2523);
    or g3702(n7655 ,n7609 ,n7575);
    not g3703(n5403 ,n5402);
    xor g3704(n7842 ,n3901 ,n3908);
    or g3705(n1730 ,n1370 ,n1177);
    nor g3706(n616 ,n587 ,n600);
    not g3707(n6524 ,n6523);
    nor g3708(n1204 ,n809 ,n1107);
    not g3709(n2824 ,n2823);
    nor g3710(n2640 ,n2546 ,n2596);
    not g3711(n706 ,n29[1]);
    xnor g3712(n4406 ,n4110 ,n4138);
    not g3713(n7074 ,n7073);
    nor g3714(n5198 ,n5088 ,n5105);
    nor g3715(n4210 ,n4027 ,n4018);
    nor g3716(n4070 ,n4014 ,n4019);
    not g3717(n4588 ,n4587);
    not g3718(n839 ,n34[15]);
    not g3719(n964 ,n30[2]);
    xnor g3720(n5820 ,n5134 ,n5362);
    buf g3721(n14[1], n11[1]);
    nor g3722(n2649 ,n2535 ,n2604);
    not g3723(n168 ,n167);
    nor g3724(n2584 ,n2500 ,n2556);
    not g3725(n5746 ,n5745);
    dff g3726(.RN(n1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n29[4]));
    nor g3727(n4287 ,n4078 ,n4100);
    nor g3728(n5500 ,n5117 ,n5090);
    not g3729(n2732 ,n2731);
    nor g3730(n2674 ,n2513 ,n2632);
    xnor g3731(n1029 ,n882 ,n836);
    nor g3732(n2976 ,n2970 ,n2964);
    nor g3733(n4290 ,n4094 ,n4098);
    nor g3734(n6726 ,n6575 ,n6614);
    nor g3735(n4206 ,n4029 ,n4019);
    dff g3736(.RN(n1), .SN(1'b1), .CK(n0), .D(n1629), .Q(n11[6]));
    nor g3737(n5974 ,n5691 ,n5881);
    not g3738(n3726 ,n3725);
    nor g3739(n74 ,n56 ,n73);
    xnor g3740(n6511 ,n6277 ,n6118);
    nor g3741(n1446 ,n853 ,n634);
    nor g3742(n2065 ,n1892 ,n2004);
    or g3743(n7656 ,n7581 ,n7580);
    nor g3744(n4046 ,n4013 ,n4006);
    nor g3745(n2235 ,n2175 ,n2199);
    nor g3746(n1243 ,n833 ,n640);
    or g3747(n3041 ,n3023 ,n3025);
    or g3748(n1764 ,n1403 ,n1546);
    not g3749(n6528 ,n6527);
    or g3750(n1685 ,n1337 ,n1123);
    nor g3751(n3816 ,n3772 ,n3815);
    not g3752(n2327 ,n2326);
    nor g3753(n4809 ,n4531 ,n4720);
    nor g3754(n1490 ,n782 ,n639);
    nor g3755(n6368 ,n6019 ,n6116);
    nor g3756(n6820 ,n6619 ,n6738);
    not g3757(n814 ,n27[2]);
    nor g3758(n3104 ,n3013 ,n3030);
    xnor g3759(n39[3] ,n2831 ,n2814);
    not g3760(n963 ,n33[6]);
    not g3761(n3413 ,n3412);
    nor g3762(n1987 ,n1901 ,n1974);
    xnor g3763(n1054 ,n686 ,n815);
    not g3764(n3865 ,n7793);
    nor g3765(n7062 ,n6963 ,n7013);
    nor g3766(n161 ,n160 ,n157);
    xnor g3767(n1035 ,n36[11] ,n34[11]);
    not g3768(n929 ,n11[7]);
    xor g3769(n5764 ,n5517 ,n5354);
    xnor g3770(n6187 ,n5767 ,n5276);
    nor g3771(n6328 ,n5850 ,n6193);
    nor g3772(n5719 ,n5159 ,n5243);
    not g3773(n5265 ,n5264);
    nor g3774(n1015 ,n643 ,n18[1]);
    or g3775(n1701 ,n1350 ,n1531);
    nor g3776(n5434 ,n5119 ,n5091);
    xor g3777(n7733 ,n3550 ,n3579);
    nor g3778(n2554 ,n2442 ,n2525);
    nor g3779(n5653 ,n5210 ,n5462);
    nor g3780(n7153 ,n7044 ,n7122);
    nor g3781(n4999 ,n4926 ,n4980);
    xnor g3782(n6597 ,n6389 ,n6481);
    not g3783(n970 ,n35[9]);
    nor g3784(n5388 ,n5118 ,n5104);
    not g3785(n939 ,n11[1]);
    nor g3786(n5757 ,n5560 ,n5580);
    not g3787(n5367 ,n5366);
    nor g3788(n7575 ,n7379 ,n7475);
    xnor g3789(n6784 ,n6644 ,n6700);
    not g3790(n7381 ,n40[7]);
    xnor g3791(n341 ,n237 ,n243);
    nor g3792(n2988 ,n2976 ,n2987);
    not g3793(n2913 ,n2912);
    nor g3794(n5986 ,n5688 ,n5885);
    nor g3795(n1389 ,n917 ,n1101);
    nor g3796(n5655 ,n5402 ,n5250);
    xnor g3797(n2135 ,n1971 ,n2087);
    not g3798(n4039 ,n4038);
    not g3799(n2994 ,n7755);
    xnor g3800(n2518 ,n2425 ,n2503);
    nor g3801(n4305 ,n4066 ,n4076);
    xnor g3802(n5839 ,n5535 ,n5553);
    not g3803(n5117 ,n37[1]);
    nor g3804(n1812 ,n1100 ,n1807);
    or g3805(n1770 ,n1409 ,n1499);
    not g3806(n527 ,n526);
    nor g3807(n1422 ,n860 ,n640);
    xnor g3808(n1848 ,n617 ,n622);
    or g3809(n1606 ,n1268 ,n1482);
    nor g3810(n5208 ,n5118 ,n5094);
    nor g3811(n1570 ,n679 ,n634);
    xnor g3812(n1940 ,n20[1] ,n19[1]);
    dff g3813(.RN(n1), .SN(1'b1), .CK(n0), .D(n1651), .Q(n35[12]));
    not g3814(n4761 ,n4760);
    nor g3815(n6010 ,n5755 ,n5840);
    nor g3816(n366 ,n198 ,n295);
    nor g3817(n1203 ,n813 ,n1107);
    not g3818(n3293 ,n3292);
    xor g3819(n40[13] ,n39[14] ,n7826);
    not g3820(n686 ,n16[7]);
    not g3821(n3502 ,n3501);
    nor g3822(n2250 ,n2178 ,n2236);
    nor g3823(n7212 ,n7100 ,n7165);
    not g3824(n4008 ,n37[4]);
    nor g3825(n1286 ,n921 ,n637);
    not g3826(n895 ,n24[15]);
    nor g3827(n5641 ,n5442 ,n5500);
    nor g3828(n5860 ,n5564 ,n5626);
    not g3829(n7438 ,n7815);
    nor g3830(n3313 ,n3148 ,n3207);
    nor g3831(n7285 ,n7265 ,n7229);
    dff g3832(.RN(n1), .SN(1'b1), .CK(n0), .D(n1584), .Q(n20[1]));
    not g3833(n6478 ,n6477);
    nor g3834(n3491 ,n3445 ,n3458);
    nor g3835(n3220 ,n3057 ,n3174);
    not g3836(n3384 ,n3383);
    not g3837(n3628 ,n39[4]);
    nor g3838(n497 ,n426 ,n448);
    nor g3839(n7268 ,n7240 ,n7196);
    xnor g3840(n2113 ,n1971 ,n2050);
    not g3841(n765 ,n2[5]);
    xnor g3842(n6505 ,n6287 ,n6061);
    not g3843(n7377 ,n7781);
    dff g3844(.RN(n1), .SN(1'b1), .CK(n0), .D(n1636), .Q(n10[15]));
    nor g3845(n2807 ,n2660 ,n2784);
    nor g3846(n1953 ,n1930 ,n1924);
    nor g3847(n3174 ,n2995 ,n3067);
    xnor g3848(n6535 ,n6289 ,n6052);
    not g3849(n6789 ,n6788);
    xnor g3850(n2471 ,n2448 ,n21[6]);
    or g3851(n1756 ,n1394 ,n1157);
    nor g3852(n4698 ,n4598 ,n4640);
    xnor g3853(n7024 ,n6868 ,n6938);
    nor g3854(n4156 ,n4014 ,n4006);
    nor g3855(n7585 ,n7392 ,n7481);
    nor g3856(n5876 ,n5539 ,n5609);
    xnor g3857(n3952 ,n7789 ,n7774);
    nor g3858(n7229 ,n7199 ,n7148);
    nor g3859(n3918 ,n3888 ,n3917);
    not g3860(n3001 ,n7748);
    nor g3861(n3086 ,n2995 ,n3031);
    not g3862(n6427 ,n6426);
    nor g3863(n3529 ,n3491 ,n3511);
    nor g3864(n2061 ,n1891 ,n2027);
    nor g3865(n6811 ,n6606 ,n6754);
    not g3866(n5560 ,n5559);
    nor g3867(n3303 ,n3103 ,n3249);
    nor g3868(n2047 ,n1901 ,n2003);
    nor g3869(n5410 ,n5118 ,n5105);
    nor g3870(n4455 ,n4303 ,n4408);
    nor g3871(n3152 ,n2994 ,n3072);
    nor g3872(n5631 ,n5444 ,n5464);
    xnor g3873(n2882 ,n2853 ,n2823);
    nor g3874(n3546 ,n3502 ,n3510);
    nor g3875(n2545 ,n2441 ,n2519);
    nor g3876(n7506 ,n7380 ,n7475);
    xnor g3877(n4386 ,n4090 ,n4200);
    nor g3878(n7056 ,n7015 ,n6935);
    nor g3879(n5027 ,n4908 ,n5000);
    nor g3880(n1385 ,n700 ,n642);
    or g3881(n1726 ,n1367 ,n1176);
    xnor g3882(n7825 ,n3959 ,n3990);
    nor g3883(n1521 ,n781 ,n641);
    not g3884(n2853 ,n2852);
    or g3885(n1092 ,n981 ,n980);
    dff g3886(.RN(n1), .SN(1'b1), .CK(n0), .D(n1744), .Q(n29[7]));
    xnor g3887(n481 ,n395 ,n419);
    nor g3888(n1127 ,n635 ,n1058);
    nor g3889(n5620 ,n5202 ,n5468);
    nor g3890(n3300 ,n3146 ,n3248);
    nor g3891(n3182 ,n3013 ,n3071);
    nor g3892(n2074 ,n2022 ,n2053);
    not g3893(n801 ,n1873);
    xnor g3894(n354 ,n165 ,n201);
    nor g3895(n2069 ,n2011 ,n2037);
    or g3896(n1590 ,n1248 ,n1473);
    nor g3897(n5942 ,n5712 ,n5924);
    nor g3898(n5522 ,n5108 ,n5111);
    xnor g3899(n7301 ,n7278 ,n7276);
    nor g3900(n2500 ,n2444 ,n2477);
    not g3901(n2766 ,n2765);
    xor g3902(n5805 ,n5345 ,n5234);
    not g3903(n4093 ,n4092);
    buf g3904(n15[7], 1'b0);
    nor g3905(n6356 ,n5974 ,n6149);
    not g3906(n2161 ,n1884);
    or g3907(n1826 ,n1083 ,n1819);
    nor g3908(n3124 ,n2994 ,n3062);
    xnor g3909(n2729 ,n2513 ,n2637);
    not g3910(n4181 ,n4180);
    nor g3911(n3650 ,n3590 ,n3602);
    dff g3912(.RN(n1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n16[7]));
    not g3913(n2278 ,n2277);
    nor g3914(n6034 ,n5727 ,n5914);
    not g3915(n3018 ,n40[11]);
    nor g3916(n2060 ,n1901 ,n2027);
    not g3917(n7350 ,n40[13]);
    not g3918(n731 ,n1880);
    not g3919(n5034 ,n5033);
    nor g3920(n3912 ,n3898 ,n3911);
    not g3921(n5353 ,n5352);
    xnor g3922(n3378 ,n3355 ,n3243);
    not g3923(n661 ,n17[3]);
    nor g3924(n1425 ,n842 ,n1105);
    not g3925(n5161 ,n5160);
    nor g3926(n3410 ,n3285 ,n3371);
    not g3927(n3604 ,n7802);
    nor g3928(n2054 ,n1892 ,n2002);
    not g3929(n3269 ,n3268);
    not g3930(n3242 ,n3241);
    nor g3931(n7038 ,n6919 ,n6988);
    xnor g3932(n3551 ,n3505 ,n3489);
    xnor g3933(n4856 ,n4729 ,n4781);
    dff g3934(.RN(n1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n21[2]));
    nor g3935(n6849 ,n6769 ,n6810);
    nor g3936(n7504 ,n7367 ,n7475);
    nor g3937(n2493 ,n2464 ,n2483);
    xnor g3938(n6709 ,n6579 ,n6471);
    not g3939(n282 ,n281);
    not g3940(n7102 ,n7101);
    xor g3941(n6392 ,n6160 ,n6265);
    nor g3942(n1414 ,n887 ,n638);
    xnor g3943(n3270 ,n3124 ,n3078);
    nor g3944(n6911 ,n6760 ,n6813);
    nor g3945(n5490 ,n5101 ,n5102);
    not g3946(n4029 ,n19[7]);
    or g3947(n36[3] ,n7699 ,n7698);
    xor g3948(n1888 ,n2115 ,n2173);
    xnor g3949(n1864 ,n66 ,n69);
    nor g3950(n5650 ,n5156 ,n5184);
    not g3951(n232 ,n231);
    nor g3952(n556 ,n501 ,n523);
    xor g3953(n40[3] ,n39[4] ,n7836);
    nor g3954(n2100 ,n1994 ,n2062);
    nor g3955(n7518 ,n7423 ,n7479);
    nor g3956(n2657 ,n2553 ,n2610);
    or g3957(n36[9] ,n7696 ,n7692);
    xnor g3958(n1045 ,n877 ,n817);
    xor g3959(n1853 ,n520 ,n509);
    nor g3960(n5909 ,n5581 ,n5616);
    nor g3961(n1508 ,n758 ,n639);
    not g3962(n666 ,n17[7]);
    nor g3963(n5751 ,n5554 ,n5536);
    nor g3964(n5908 ,n5339 ,n5633);
    xnor g3965(n6864 ,n6706 ,n6573);
    nor g3966(n3662 ,n3620 ,n3601);
    nor g3967(n5065 ,n5036 ,n5050);
    nor g3968(n3978 ,n3938 ,n3977);
    not g3969(n955 ,n11[15]);
    xnor g3970(n7288 ,n7200 ,n7268);
    nor g3971(n2387 ,n2368 ,n2364);
    nor g3972(n4278 ,n4232 ,n4032);
    nor g3973(n5007 ,n4933 ,n4973);
    not g3974(n400 ,n399);
    xnor g3975(n4563 ,n4376 ,n4192);
    nor g3976(n1193 ,n1009 ,n1104);
    not g3977(n752 ,n1844);
    not g3978(n327 ,n326);
    not g3979(n4187 ,n4186);
    nor g3980(n606 ,n592 ,n585);
    not g3981(n854 ,n34[8]);
    not g3982(n7391 ,n26[1]);
    xnor g3983(n4603 ,n4509 ,n4462);
    nor g3984(n1162 ,n1102 ,n1065);
    xnor g3985(n6509 ,n6294 ,n5962);
    xnor g3986(n4832 ,n4716 ,n4637);
    xnor g3987(n4904 ,n4818 ,n4763);
    not g3988(n5520 ,n5519);
    dff g3989(.RN(n1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n16[5]));
    nor g3990(n7316 ,n7305 ,n7315);
    nor g3991(n488 ,n407 ,n456);
    not g3992(n3145 ,n3144);
    not g3993(n1942 ,n20[0]);
    nor g3994(n5852 ,n5382 ,n5751);
    not g3995(n6169 ,n6168);
    not g3996(n5179 ,n5178);
    not g3997(n4459 ,n4458);
    nor g3998(n6605 ,n6565 ,n6545);
    nor g3999(n5697 ,n5259 ,n5419);
    or g4000(n1605 ,n1267 ,n1117);
    xnor g4001(n6152 ,n5822 ,n5370);
    xor g4002(n6165 ,n5801 ,n5222);
    xnor g4003(n6976 ,n6874 ,n6798);
    nor g4004(n3815 ,n3769 ,n3814);
    nor g4005(n1290 ,n930 ,n636);
    nor g4006(n1263 ,n722 ,n636);
    xnor g4007(n2210 ,n2143 ,n2162);
    nor g4008(n1141 ,n641 ,n1087);
    dff g4009(.RN(n1), .SN(1'b1), .CK(n0), .D(n1690), .Q(n24[11]));
    not g4010(n7370 ,n39[3]);
    nor g4011(n4572 ,n4479 ,n4488);
    nor g4012(n4507 ,n4331 ,n4444);
    not g4013(n859 ,n28[1]);
    xnor g4014(n7787 ,n5070 ,n5075);
    nor g4015(n3275 ,n3253 ,n3237);
    or g4016(n1700 ,n1349 ,n1449);
    nor g4017(n362 ,n268 ,n299);
    not g4018(n7385 ,n7726);
    or g4019(n4253 ,n4007 ,n4026);
    xnor g4020(n7788 ,n5071 ,n5077);
    nor g4021(n7609 ,n7375 ,n7478);
    nor g4022(n4062 ,n4022 ,n4028);
    nor g4023(n7240 ,n7213 ,n7235);
    not g4024(n7259 ,n7258);
    not g4025(n3027 ,n7753);
    dff g4026(.RN(n1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n29[3]));
    or g4027(n36[10] ,n7701 ,n7700);
    not g4028(n2684 ,n2683);
    not g4029(n788 ,n1864);
    or g4030(n1096 ,n998 ,n984);
    nor g4031(n2823 ,n2752 ,n2795);
    xnor g4032(n438 ,n332 ,n277);
    nor g4033(n4121 ,n4007 ,n4016);
    xnor g4034(n1069 ,n810 ,n844);
    not g4035(n957 ,n12[7]);
    not g4036(n3664 ,n3663);
    xnor g4037(n3062 ,n7754 ,n7759);
    nor g4038(n1224 ,n661 ,n1105);
    nor g4039(n2563 ,n2443 ,n2525);
    xnor g4040(n1931 ,n1896 ,n19[4]);
    nor g4041(n3834 ,n37[1] ,n19[1]);
    nor g4042(n4492 ,n4414 ,n4409);
    nor g4043(n5202 ,n5096 ,n5117);
    nor g4044(n629 ,n589 ,n628);
    not g4045(n879 ,n32[2]);
    nor g4046(n6818 ,n6657 ,n6727);
    nor g4047(n1440 ,n933 ,n638);
    or g4048(n7479 ,n7326 ,n7465);
    nor g4049(n6698 ,n6566 ,n6546);
    nor g4050(n1371 ,n665 ,n1101);
    not g4051(n952 ,n35[13]);
    not g4052(n2911 ,n2910);
    nor g4053(n1384 ,n948 ,n1101);
    not g4054(n2078 ,n2079);
    nor g4055(n5997 ,n5739 ,n5905);
    xnor g4056(n2111 ,n1959 ,n2033);
    not g4057(n1893 ,n37[2]);
    not g4058(n4207 ,n4206);
    nor g4059(n6607 ,n6539 ,n6495);
    not g4060(n6871 ,n6870);
    not g4061(n767 ,n3[6]);
    nor g4062(n110 ,n25[3] ,n108);
    dff g4063(.RN(n1), .SN(1'b1), .CK(n0), .D(n1707), .Q(n24[5]));
    nor g4064(n4888 ,n4794 ,n4837);
    not g4065(n4627 ,n4626);
    not g4066(n876 ,n32[5]);
    not g4067(n6246 ,n6245);
    nor g4068(n1123 ,n634 ,n1061);
    or g4069(n1749 ,n1389 ,n1147);
    not g4070(n2464 ,n2463);
    nor g4071(n6214 ,n5744 ,n5956);
    nor g4072(n2118 ,n1958 ,n2100);
    not g4073(n3534 ,n3533);
    nor g4074(n3265 ,n3083 ,n3180);
    xnor g4075(n2315 ,n2277 ,n2254);
    not g4076(n856 ,n23[4]);
    nor g4077(n4579 ,n4177 ,n4470);
    xnor g4078(n2341 ,n1886 ,n2297);
    not g4079(n7160 ,n7159);
    nor g4080(n563 ,n495 ,n525);
    nor g4081(n3186 ,n3013 ,n3070);
    xnor g4082(n3896 ,n41[13] ,n7814);
    nor g4083(n3795 ,n3742 ,n3767);
    not g4084(n3717 ,n3716);
    not g4085(n3155 ,n3154);
    xnor g4086(n5788 ,n5124 ,n5474);
    nor g4087(n6486 ,n6192 ,n6327);
    xnor g4088(n6650 ,n6407 ,n6187);
    not g4089(n2734 ,n2733);
    nor g4090(n7499 ,n7438 ,n7477);
    xnor g4091(n7844 ,n3895 ,n3903);
    not g4092(n3464 ,n3463);
    nor g4093(n77 ,n65 ,n76);
    not g4094(n863 ,n21[6]);
    nor g4095(n2620 ,n2567 ,n2594);
    nor g4096(n6228 ,n6051 ,n5977);
    xnor g4097(n582 ,n545 ,n526);
    nor g4098(n5482 ,n5100 ,n5104);
    nor g4099(n3364 ,n3295 ,n3349);
    not g4100(n7405 ,n7784);
    nor g4101(n3495 ,n3419 ,n3470);
    not g4102(n2510 ,n2511);
    nor g4103(n5685 ,n5477 ,n5143);
    not g4104(n4205 ,n4204);
    not g4105(n5939 ,n5938);
    not g4106(n690 ,n16[5]);
    not g4107(n6635 ,n6634);
    nor g4108(n6919 ,n6829 ,n6858);
    nor g4109(n7463 ,n41[6] ,n7822);
    not g4110(n4901 ,n4900);
    not g4111(n787 ,n6[2]);
    nor g4112(n2533 ,n2434 ,n2521);
    xnor g4113(n7840 ,n3899 ,n3913);
    nor g4114(n3814 ,n3762 ,n3813);
    xnor g4115(n6636 ,n6401 ,n6259);
    nor g4116(n3350 ,n3230 ,n3287);
    xnor g4117(n3788 ,n3735 ,n3701);
    not g4118(n6805 ,n6804);
    xnor g4119(n1027 ,n889 ,n891);
    not g4120(n4833 ,n4832);
    or g4121(n7475 ,n26[0] ,n7324);
    nor g4122(n2000 ,n1890 ,n1976);
    nor g4123(n7544 ,n7437 ,n7481);
    not g4124(n3432 ,n3431);
    nor g4125(n4190 ,n4014 ,n4008);
    nor g4126(n7318 ,n7294 ,n7317);
    nor g4127(n3271 ,n3104 ,n3242);
    nor g4128(n3584 ,n3560 ,n3583);
    nor g4129(n7105 ,n7010 ,n7027);
    nor g4130(n6924 ,n6806 ,n6850);
    nor g4131(n265 ,n147 ,n157);
    xnor g4132(n1031 ,n869 ,n850);
    nor g4133(n1530 ,n776 ,n641);
    not g4134(n935 ,n12[13]);
    nor g4135(n138 ,n123 ,n136);
    nor g4136(n2170 ,n2006 ,n2117);
    nor g4137(n5865 ,n5347 ,n5621);
    xnor g4138(n6108 ,n5769 ,n5372);
    nor g4139(n105 ,n101 ,n98);
    not g4140(n5529 ,n5528);
    not g4141(n3109 ,n3108);
    nor g4142(n6323 ,n6154 ,n6152);
    nor g4143(n6730 ,n6441 ,n6690);
    or g4144(n85 ,n25[3] ,n25[2]);
    nor g4145(n2376 ,n2329 ,n2352);
    nor g4146(n3878 ,n7814 ,n41[13]);
    not g4147(n4131 ,n4130);
    nor g4148(n241 ,n145 ,n157);
    xnor g4149(n39[15] ,n2943 ,n2993);
    or g4150(n7485 ,n7460 ,n7480);
    nor g4151(n6061 ,n5695 ,n5897);
    nor g4152(n1173 ,n1102 ,n1030);
    nor g4153(n5643 ,n5252 ,n5392);
    not g4154(n7344 ,n40[5]);
    xnor g4155(n405 ,n340 ,n173);
    or g4156(n1618 ,n1284 ,n1489);
    nor g4157(n6202 ,n6022 ,n5966);
    not g4158(n768 ,n1879);
    nor g4159(n7090 ,n7022 ,n7054);
    xnor g4160(n4530 ,n4387 ,n4108);
    nor g4161(n2039 ,n1890 ,n2002);
    nor g4162(n3707 ,n3661 ,n3682);
    nor g4163(n4813 ,n4663 ,n4752);
    xnor g4164(n7794 ,n6602 ,n6239);
    nor g4165(n2491 ,n2462 ,n2474);
    not g4166(n3623 ,n39[11]);
    dff g4167(.RN(n1), .SN(1'b1), .CK(n0), .D(n1625), .Q(n1832));
    not g4168(n7412 ,n7787);
    xnor g4169(n2666 ,n2501 ,n2581);
    not g4170(n1899 ,n20[0]);
    dff g4171(.RN(n1), .SN(1'b1), .CK(n0), .D(n1639), .Q(n10[12]));
    nor g4172(n1276 ,n879 ,n1103);
    not g4173(n2927 ,n2926);
    xnor g4174(n4859 ,n4785 ,n4634);
    nor g4175(n4351 ,n4131 ,n4119);
    nor g4176(n5284 ,n5119 ,n5090);
    nor g4177(n3819 ,n3759 ,n3818);
    nor g4178(n5348 ,n5103 ,n5111);
    xnor g4179(n6844 ,n6599 ,n6743);
    or g4180(n7688 ,n7632 ,n7628);
    not g4181(n6542 ,n6541);
    dff g4182(.RN(n1), .SN(1'b1), .CK(n0), .D(n1609), .Q(n12[1]));
    not g4183(n5119 ,n37[3]);
    dff g4184(.RN(n1), .SN(1'b1), .CK(n0), .D(n1745), .Q(n29[6]));
    nor g4185(n2625 ,n2569 ,n2611);
    or g4186(n1721 ,n1227 ,n1539);
    nor g4187(n6381 ,n6143 ,n6139);
    or g4188(n1652 ,n1433 ,n1553);
    not g4189(n715 ,n19[6]);
    nor g4190(n361 ,n206 ,n287);
    not g4191(n4067 ,n4066);
    or g4192(n1181 ,n27[0] ,n1095);
    nor g4193(n1449 ,n801 ,n634);
    xnor g4194(n1049 ,n659 ,n670);
    not g4195(n673 ,n34[14]);
    not g4196(n3829 ,n19[0]);
    not g4197(n5101 ,n22[5]);
    not g4198(n4073 ,n4072);
    or g4199(n1734 ,n1374 ,n1187);
    nor g4200(n3118 ,n3013 ,n3036);
    or g4201(n7637 ,n7541 ,n7540);
    nor g4202(n2715 ,n2575 ,n2663);
    nor g4203(n6902 ,n6625 ,n6821);
    or g4204(n5338 ,n5100 ,n5110);
    not g4205(n923 ,n11[5]);
    xnor g4206(n3954 ,n7785 ,n7770);
    not g4207(n5293 ,n5292);
    not g4208(n240 ,n239);
    xnor g4209(n2147 ,n1970 ,n2096);
    nor g4210(n7272 ,n7268 ,n7200);
    nor g4211(n4194 ,n4014 ,n4018);
    xnor g4212(n4528 ,n4374 ,n4258);
    nor g4213(n4349 ,n4237 ,n4136);
    nor g4214(n4265 ,n4023 ,n4020);
    nor g4215(n6386 ,n6256 ,n6252);
    nor g4216(n1261 ,n876 ,n1103);
    nor g4217(n3701 ,n3653 ,n3686);
    nor g4218(n3342 ,n3233 ,n3274);
    nor g4219(n3768 ,n3715 ,n3743);
    not g4220(n4403 ,n4402);
    nor g4221(n1250 ,n852 ,n640);
    nor g4222(n3478 ,n3384 ,n3428);
    nor g4223(n7567 ,n7442 ,n7474);
    xor g4224(n5777 ,n5340 ,n5136);
    xnor g4225(n6422 ,n6073 ,n6058);
    xnor g4226(n6491 ,n6098 ,n6334);
    nor g4227(n6662 ,n6485 ,n6558);
    nor g4228(n633 ,n492 ,n632);
    nor g4229(n3097 ,n2994 ,n3028);
    nor g4230(n2849 ,n2820 ,n2829);
    nor g4231(n5204 ,n5092 ,n5116);
    nor g4232(n5352 ,n5108 ,n5094);
    xnor g4233(n2082 ,n1971 ,n2008);
    nor g4234(n1153 ,n1100 ,n1073);
    dff g4235(.RN(n1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n21[4]));
    xnor g4236(n2502 ,n2482 ,n2463);
    not g4237(n6647 ,n6646);
    xnor g4238(n2943 ,n2883 ,n2914);
    nor g4239(n3762 ,n3713 ,n3739);
    nor g4240(n459 ,n321 ,n434);
    not g4241(n100 ,n25[3]);
    not g4242(n596 ,n595);
    xnor g4243(n5774 ,n5384 ,n5272);
    nor g4244(n2330 ,n2289 ,n2292);
    nor g4245(n1549 ,n724 ,n1100);
    nor g4246(n5424 ,n5089 ,n5097);
    dff g4247(.RN(n1), .SN(1'b1), .CK(n0), .D(n1590), .Q(n16[4]));
    nor g4248(n193 ,n159 ,n148);
    nor g4249(n4341 ,n4051 ,n4189);
    xnor g4250(n4598 ,n4363 ,n4408);
    nor g4251(n2354 ,n2303 ,n2335);
    xnor g4252(n1072 ,n24[5] ,n35[5]);
    nor g4253(n2293 ,n2220 ,n2270);
    not g4254(n4541 ,n4540);
    nor g4255(n6589 ,n6369 ,n6446);
    not g4256(n4523 ,n4522);
    not g4257(n4136 ,n4135);
    not g4258(n2159 ,n2160);
    nor g4259(n7012 ,n6878 ,n6929);
    not g4260(n3508 ,n3507);
    not g4261(n4362 ,n4361);
    nor g4262(n4256 ,n4019 ,n4024);
    not g4263(n6791 ,n6790);
    nor g4264(n1452 ,n855 ,n634);
    nor g4265(n5402 ,n5119 ,n5093);
    xnor g4266(n5766 ,n5458 ,n5174);
    nor g4267(n3358 ,n3234 ,n3277);
    xnor g4268(n7077 ,n6978 ,n6870);
    not g4269(n7293 ,n7292);
    or g4270(n995 ,n35[1] ,n35[7]);
    dff g4271(.RN(n1), .SN(1'b1), .CK(n0), .D(n1741), .Q(n17[5]));
    or g4272(n36[1] ,n7691 ,n7705);
    not g4273(n4564 ,n4563);
    or g4274(n1791 ,n1202 ,n1559);
    nor g4275(n59 ,n45 ,n42);
    not g4276(n6822 ,n6821);
    not g4277(n2225 ,n2224);
    nor g4278(n3304 ,n3106 ,n3258);
    not g4279(n6637 ,n6636);
    not g4280(n3540 ,n3539);
    xnor g4281(n4526 ,n4386 ,n4238);
    nor g4282(n7565 ,n7351 ,n7478);
    xnor g4283(n6132 ,n5779 ,n5506);
    nor g4284(n2320 ,n1886 ,n2297);
    xnor g4285(n5837 ,n5315 ,n5352);
    nor g4286(n7210 ,n7118 ,n7170);
    not g4287(n638 ,n639);
    nor g4288(n4434 ,n4140 ,n4295);
    xnor g4289(n5021 ,n4955 ,n4977);
    nor g4290(n1947 ,n1918 ,n1933);
    xnor g4291(n3892 ,n41[14] ,n7815);
    xor g4292(n5768 ,n5308 ,n5476);
    xnor g4293(n333 ,n225 ,n223);
    xor g4294(n38[1] ,n7845 ,n39[1]);
    xnor g4295(n2509 ,n2495 ,n2478);
    not g4296(n2750 ,n2749);
    nor g4297(n6430 ,n6190 ,n6311);
    nor g4298(n2046 ,n1891 ,n2002);
    xnor g4299(n2157 ,n1968 ,n2076);
    nor g4300(n4890 ,n4798 ,n4838);
    nor g4301(n2461 ,n2451 ,n2435);
    xnor g4302(n6090 ,n5765 ,n5126);
    nor g4303(n5881 ,n5335 ,n5594);
    nor g4304(n2072 ,n2000 ,n2043);
    not g4305(n3390 ,n3389);
    dff g4306(.RN(n1), .SN(1'b1), .CK(n0), .D(n1653), .Q(n10[1]));
    nor g4307(n1485 ,n747 ,n639);
    not g4308(n3625 ,n7783);
    or g4309(n7480 ,n7326 ,n7323);
    not g4310(n1939 ,n1938);
    nor g4311(n3285 ,n3159 ,n3243);
    nor g4312(n1815 ,n993 ,n1808);
    nor g4313(n470 ,n405 ,n404);
    dff g4314(.RN(n1), .SN(1'b1), .CK(n0), .D(n1624), .Q(n11[9]));
    xnor g4315(n2704 ,n2514 ,n2628);
    xor g4316(n6177 ,n5832 ,n5160);
    not g4317(n123 ,n33[4]);
    nor g4318(n7505 ,n7381 ,n7478);
    or g4319(n36[2] ,n7695 ,n7693);
    or g4320(n7641 ,n7525 ,n7524);
    nor g4321(n4637 ,n4451 ,n4569);
    nor g4322(n2073 ,n1990 ,n2046);
    xnor g4323(n3361 ,n3292 ,n3212);
    xor g4324(n7732 ,n3567 ,n3577);
    or g4325(n1793 ,n1430 ,n1508);
    nor g4326(n78 ,n60 ,n77);
    not g4327(n2857 ,n2856);
    buf g4328(n14[11], n11[11]);
    nor g4329(n6311 ,n6055 ,n6226);
    or g4330(n639 ,n18[2] ,n979);
    nor g4331(n5737 ,n5161 ,n5495);
    xnor g4332(n7198 ,n7139 ,n7155);
    xnor g4333(n3737 ,n39[11] ,n3667);
    xnor g4334(n5016 ,n4981 ,n4951);
    not g4335(n4905 ,n4904);
    not g4336(n3492 ,n3491);
    xnor g4337(n7762 ,n3845 ,n3839);
    nor g4338(n3822 ,n3775 ,n3821);
    xnor g4339(n5841 ,n5290 ,n5341);
    not g4340(n705 ,n10[2]);
    dff g4341(.RN(n1), .SN(1'b1), .CK(n0), .D(n1688), .Q(n34[2]));
    xnor g4342(n3846 ,n37[4] ,n19[4]);
    nor g4343(n4198 ,n4008 ,n4024);
    dff g4344(.RN(n1), .SN(1'b1), .CK(n0), .D(n1747), .Q(n23[2]));
    xnor g4345(n398 ,n370 ,n183);
    or g4346(n1782 ,n1419 ,n1504);
    not g4347(n2191 ,n2190);
    or g4348(n36[14] ,n7694 ,n7707);
    xnor g4349(n3341 ,n3102 ,n3249);
    nor g4350(n7555 ,n7371 ,n7476);
    nor g4351(n120 ,n97 ,n118);
    nor g4352(n5889 ,n5312 ,n5602);
    not g4353(n679 ,n36[8]);
    not g4354(n3103 ,n3102);
    nor g4355(n5268 ,n5099 ,n5116);
    not g4356(n414 ,n413);
    nor g4357(n5464 ,n5091 ,n5113);
    nor g4358(n4850 ,n4816 ,n4780);
    not g4359(n3400 ,n3399);
    nor g4360(n1121 ,n634 ,n1047);
    or g4361(n1694 ,n1317 ,n1529);
    xnor g4362(n7308 ,n7292 ,n7274);
    nor g4363(n3839 ,n3828 ,n3829);
    nor g4364(n5069 ,n5041 ,n5055);
    nor g4365(n2986 ,n2985 ,n2967);
    xor g4366(n5832 ,n5510 ,n5494);
    xnor g4367(n2870 ,n2806 ,n2747);
    not g4368(n5993 ,n5992);
    nor g4369(n590 ,n533 ,n575);
    not g4370(n4087 ,n4086);
    not g4371(n6419 ,n6418);
    xnor g4372(n4830 ,n4715 ,n4719);
    nor g4373(n1377 ,n711 ,n1105);
    nor g4374(n6036 ,n5689 ,n5899);
    not g4375(n3317 ,n3316);
    not g4376(n871 ,n31[2]);
    dff g4377(.RN(n1), .SN(1'b1), .CK(n0), .D(n1738), .Q(n23[4]));
    nor g4378(n7667 ,n7466 ,n7482);
    nor g4379(n3309 ,n3252 ,n3262);
    xor g4380(n4562 ,n4381 ,n4242);
    nor g4381(n2644 ,n2543 ,n2603);
    nor g4382(n5362 ,n5088 ,n5114);
    nor g4383(n6058 ,n5728 ,n5877);
    nor g4384(n4238 ,n4022 ,n4010);
    nor g4385(n5673 ,n5263 ,n5365);
    nor g4386(n3373 ,n3239 ,n3338);
    not g4387(n734 ,n1870);
    nor g4388(n3289 ,n3156 ,n3217);
    xnor g4389(n3072 ,n40[8] ,n7747);
    nor g4390(n3637 ,n39[12] ,n7813);
    not g4391(n3428 ,n3427);
    nor g4392(n1208 ,n817 ,n642);
    nor g4393(n5869 ,n5538 ,n5666);
    nor g4394(n7042 ,n6955 ,n7004);
    xnor g4395(n2141 ,n2088 ,n1970);
    not g4396(n212 ,n211);
    xnor g4397(n6541 ,n6285 ,n6158);
    xnor g4398(n7099 ,n6984 ,n7020);
    nor g4399(n1321 ,n943 ,n637);
    or g4400(n1676 ,n1322 ,n1523);
    nor g4401(n6553 ,n6361 ,n6440);
    not g4402(n4059 ,n4058);
    nor g4403(n1333 ,n670 ,n637);
    xnor g4404(n6400 ,n6142 ,n6138);
    xor g4405(n7735 ,n3569 ,n3583);
    nor g4406(n1379 ,n964 ,n1105);
    nor g4407(n5711 ,n5181 ,n5429);
    xnor g4408(n7784 ,n5017 ,n5032);
    nor g4409(n2194 ,n2109 ,n2161);
    nor g4410(n3797 ,n3741 ,n3795);
    nor g4411(n6746 ,n6590 ,n6694);
    not g4412(n7166 ,n7165);
    xnor g4413(n2383 ,n2341 ,n2301);
    nor g4414(n6606 ,n6424 ,n6499);
    nor g4415(n2420 ,n2387 ,n2419);
    nor g4416(n7580 ,n7430 ,n7477);
    not g4417(n6023 ,n6022);
    nor g4418(n435 ,n319 ,n373);
    not g4419(n208 ,n207);
    not g4420(n7337 ,n7823);
    nor g4421(n2238 ,n1889 ,n2198);
    xor g4422(n4372 ,n4264 ,n4170);
    xnor g4423(n4921 ,n4867 ,n4865);
    or g4424(n1725 ,n1365 ,n1166);
    nor g4425(n5480 ,n5089 ,n5103);
    nor g4426(n2616 ,n2431 ,n2549);
    not g4427(n3719 ,n3718);
    xnor g4428(n2843 ,n2776 ,n2691);
    not g4429(n3017 ,n40[5]);
    nor g4430(n4679 ,n4602 ,n4616);
    nor g4431(n6042 ,n5690 ,n5926);
    xnor g4432(n7717 ,n3782 ,n3797);
    nor g4433(n4092 ,n4013 ,n4021);
    not g4434(n7065 ,n7064);
    nor g4435(n2012 ,n1901 ,n1980);
    not g4436(n1926 ,n1925);
    xnor g4437(n7772 ,n3897 ,n3921);
    nor g4438(n1537 ,n777 ,n641);
    xnor g4439(n1066 ,n814 ,n829);
    nor g4440(n6961 ,n6830 ,n6859);
    not g4441(n5302 ,n5301);
    xnor g4442(n2889 ,n2830 ,n2767);
    not g4443(n5491 ,n5490);
    or g4444(n7488 ,n7462 ,n7480);
    not g4445(n5744 ,n5743);
    not g4446(n662 ,n34[4]);
    xor g4447(n7745 ,n7807 ,n7784);
    or g4448(n1594 ,n1256 ,n1476);
    or g4449(n7676 ,n7547 ,n7668);
    nor g4450(n6001 ,n5694 ,n5860);
    xnor g4451(n3484 ,n3423 ,n3385);
    xnor g4452(n6602 ,n6120 ,n6440);
    not g4453(n6625 ,n6624);
    xor g4454(n5797 ,n5334 ,n5420);
    nor g4455(n6794 ,n6610 ,n6723);
    buf g4456(n14[10], n11[10]);
    nor g4457(n1136 ,n1841 ,n641);
    nor g4458(n463 ,n375 ,n411);
    nor g4459(n3903 ,n3873 ,n3902);
    not g4460(n6540 ,n6539);
    xnor g4461(n3747 ,n39[6] ,n3677);
    not g4462(n7082 ,n7081);
    xnor g4463(n2973 ,n2945 ,n2955);
    xnor g4464(n2480 ,n21[3] ,n22[3]);
    nor g4465(n2102 ,n1996 ,n2059);
    nor g4466(n1479 ,n779 ,n1099);
    nor g4467(n2257 ,n2160 ,n2240);
    xnor g4468(n4540 ,n4385 ,n4230);
    nor g4469(n5530 ,n5112 ,n5106);
    xor g4470(n1867 ,n33[7] ,n144);
    or g4471(n1593 ,n1255 ,n1114);
    nor g4472(n6766 ,n6700 ,n6645);
    nor g4473(n1435 ,n672 ,n640);
    nor g4474(n1271 ,n868 ,n640);
    nor g4475(n3094 ,n3012 ,n3036);
    not g4476(n6039 ,n6038);
    xnor g4477(n6847 ,n6632 ,n6775);
    nor g4478(n4288 ,n4034 ,n4162);
    not g4479(n763 ,n4[1]);
    xnor g4480(n3739 ,n39[10] ,n3668);
    nor g4481(n3100 ,n3012 ,n3035);
    nor g4482(n6819 ,n6685 ,n6742);
    xnor g4483(n4957 ,n4871 ,n4902);
    nor g4484(n5474 ,n5115 ,n5109);
    nor g4485(n5076 ,n5065 ,n5075);
    nor g4486(n4415 ,n4180 ,n4348);
    nor g4487(n388 ,n322 ,n350);
    or g4488(n1639 ,n1307 ,n1566);
    dff g4489(.RN(n1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n28[8]));
    or g4490(n1679 ,n1332 ,n1129);
    xor g4491(n5780 ,n5532 ,n5472);
    not g4492(n4939 ,n4938);
    xnor g4493(n3393 ,n3340 ,n3225);
    not g4494(n6935 ,n6934);
    xnor g4495(n41[5] ,n7193 ,n7191);
    dff g4496(.RN(n1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n17[2]));
    nor g4497(n5596 ,n5422 ,n5488);
    nor g4498(n4944 ,n4871 ,n4903);
    nor g4499(n3938 ,n7784 ,n38[7]);
    nor g4500(n7233 ,n7135 ,n7210);
    nor g4501(n1378 ,n856 ,n1103);
    nor g4502(n4699 ,n4561 ,n4623);
    not g4503(n689 ,n23[7]);
    or g4504(n7713 ,n7654 ,n7677);
    nor g4505(n2919 ,n2825 ,n2888);
    xnor g4506(n7804 ,n2266 ,n2249);
    not g4507(n3012 ,n7756);
    nor g4508(n6926 ,n6776 ,n6898);
    nor g4509(n7057 ,n7018 ,n6931);
    not g4510(n2691 ,n2690);
    nor g4511(n1126 ,n634 ,n1060);
    nor g4512(n4828 ,n4731 ,n4777);
    nor g4513(n3680 ,n3633 ,n3635);
    xnor g4514(n5015 ,n4975 ,n4915);
    nor g4515(n4765 ,n4654 ,n4693);
    or g4516(n1789 ,n1427 ,n1141);
    xnor g4517(n2115 ,n1969 ,n2049);
    not g4518(n6795 ,n6794);
    or g4519(n1592 ,n1253 ,n1113);
    nor g4520(n5432 ,n5103 ,n5105);
    nor g4521(n4435 ,n4105 ,n4285);
    nor g4522(n2850 ,n2430 ,n2827);
    dff g4523(.RN(n1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n18[0]));
    nor g4524(n1507 ,n774 ,n639);
    nor g4525(n4316 ,n4223 ,n4059);
    not g4526(n4506 ,n4505);
    nor g4527(n5703 ,n5445 ,n5465);
    nor g4528(n2878 ,n2766 ,n2843);
    xor g4529(n40[6] ,n39[7] ,n7833);
    not g4530(n5427 ,n5426);
    nor g4531(n7498 ,n7382 ,n7478);
    nor g4532(n284 ,n223 ,n225);
    not g4533(n2867 ,n2866);
    nor g4534(n3874 ,n7815 ,n41[14]);
    nor g4535(n3403 ,n3312 ,n3375);
    not g4536(n6997 ,n6996);
    xnor g4537(n2212 ,n1970 ,n2166);
    buf g4538(n13[11], n10[11]);
    xnor g4539(n4928 ,n4855 ,n4873);
    or g4540(n36[12] ,n7674 ,n7708);
    nor g4541(n263 ,n160 ,n153);
    nor g4542(n6552 ,n6482 ,n6365);
    nor g4543(n3517 ,n3477 ,n3495);
    nor g4544(n4495 ,n4325 ,n4438);
    xnor g4545(n6705 ,n6582 ,n6477);
    xnor g4546(n6628 ,n6398 ,n6173);
    nor g4547(n4477 ,n4341 ,n4433);
    nor g4548(n1361 ,n673 ,n637);
    dff g4549(.RN(n1), .SN(1'b1), .CK(n0), .D(n1701), .Q(n24[8]));
    not g4550(n106 ,n105);
    not g4551(n7427 ,n40[4]);
    not g4552(n6470 ,n6469);
    not g4553(n4985 ,n4984);
    nor g4554(n7601 ,n7354 ,n7478);
    not g4555(n3619 ,n39[10]);
    not g4556(n4043 ,n4042);
    nor g4557(n4234 ,n4019 ,n4009);
    not g4558(n325 ,n324);
    nor g4559(n4493 ,n4343 ,n4446);
    not g4560(n802 ,n5[3]);
    xnor g4561(n1030 ,n867 ,n843);
    xnor g4562(n520 ,n481 ,n435);
    xnor g4563(n6634 ,n6400 ,n6161);
    xnor g4564(n6603 ,n6328 ,n6438);
    not g4565(n2514 ,n2515);
    not g4566(n2787 ,n2786);
    nor g4567(n3140 ,n2994 ,n3064);
    xnor g4568(n483 ,n397 ,n392);
    nor g4569(n6325 ,n6064 ,n6234);
    not g4570(n7439 ,n7808);
    not g4571(n2338 ,n2337);
    nor g4572(n7245 ,n7221 ,n7177);
    or g4573(n4129 ,n4021 ,n4025);
    not g4574(n4784 ,n4783);
    nor g4575(n2556 ,n2433 ,n2525);
    nor g4576(n4967 ,n4883 ,n4928);
    nor g4577(n4436 ,n4145 ,n4284);
    nor g4578(n3981 ,n3958 ,n3980);
    xnor g4579(n417 ,n337 ,n265);
    nor g4580(n3871 ,n7811 ,n7799);
    nor g4581(n3854 ,n3841 ,n3853);
    nor g4582(n3821 ,n3774 ,n3820);
    not g4583(n146 ,n37[0]);
    xnor g4584(n1033 ,n862 ,n663);
    or g4585(n5340 ,n5116 ,n5106);
    xnor g4586(n3326 ,n3200 ,n3208);
    not g4587(n4173 ,n4172);
    not g4588(n1967 ,n1968);
    xor g4589(n1882 ,n1911 ,n1930);
    xor g4590(n5778 ,n5556 ,n5230);
    nor g4591(n6604 ,n6493 ,n6507);
    nor g4592(n2965 ,n2920 ,n2949);
    not g4593(n102 ,n25[5]);
    nor g4594(n2408 ,n2375 ,n2407);
    xor g4595(n5783 ,n5546 ,n5262);
    nor g4596(n3558 ,n3523 ,n3539);
    not g4597(n206 ,n205);
    nor g4598(n1400 ,n938 ,n642);
    nor g4599(n7534 ,n7426 ,n7480);
    nor g4600(n2821 ,n2661 ,n2785);
    nor g4601(n6771 ,n6637 ,n6635);
    xor g4602(n6176 ,n5783 ,n5364);
    not g4603(n5241 ,n5240);
    xnor g4604(n6180 ,n5808 ,n5408);
    xnor g4605(n3339 ,n3226 ,n3267);
    not g4606(n3526 ,n3525);
    not g4607(n2701 ,n2700);
    or g4608(n1616 ,n1280 ,n1442);
    dff g4609(.RN(n1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n28[9]));
    nor g4610(n5178 ,n5095 ,n5105);
    dff g4611(.RN(n1), .SN(1'b1), .CK(n0), .D(n1719), .Q(n34[13]));
    not g4612(n5514 ,n5513);
    not g4613(n4927 ,n4926);
    nor g4614(n5082 ,n5081 ,n5057);
    nor g4615(n6700 ,n6454 ,n6551);
    nor g4616(n4076 ,n4021 ,n4010);
    or g4617(n7697 ,n7633 ,n7615);
    not g4618(n927 ,n12[0]);
    not g4619(n800 ,n1871);
    dff g4620(.RN(n1), .SN(1'b1), .CK(n0), .D(n1684), .Q(n24[14]));
    xnor g4621(n6983 ,n6854 ,n6804);
    nor g4622(n4984 ,n4950 ,n4960);
    nor g4623(n7540 ,n7440 ,n7475);
    not g4624(n4933 ,n4932);
    not g4625(n7033 ,n7032);
    not g4626(n6431 ,n6430);
    xnor g4627(n1021 ,n36[13] ,n34[13]);
    nor g4628(n247 ,n159 ,n155);
    nor g4629(n6053 ,n5696 ,n5920);
    not g4630(n6081 ,n6080);
    xnor g4631(n7107 ,n6986 ,n7047);
    not g4632(n3004 ,n7750);
    nor g4633(n6945 ,n6775 ,n6895);
    nor g4634(n6011 ,n5741 ,n5931);
    nor g4635(n2345 ,n2294 ,n2319);
    nor g4636(n5037 ,n4995 ,n5026);
    xnor g4637(n3724 ,n3665 ,n39[15]);
    not g4638(n2517 ,n2516);
    nor g4639(n5921 ,n5562 ,n5647);
    not g4640(n7100 ,n7099);
    nor g4641(n52 ,n37[1] ,n19[1]);
    xor g4642(n5831 ,n5322 ,n5176);
    not g4643(n2998 ,n40[3]);
    nor g4644(n1557 ,n689 ,n1102);
    nor g4645(n6923 ,n6798 ,n6874);
    not g4646(n1018 ,n1017);
    not g4647(n6423 ,n6422);
    nor g4648(n5324 ,n5115 ,n5094);
    not g4649(n4596 ,n4595);
    dff g4650(.RN(n1), .SN(1'b1), .CK(n0), .D(n1733), .Q(n23[5]));
    nor g4651(n1354 ,n861 ,n1103);
    nor g4652(n464 ,n374 ,n412);
    not g4653(n5379 ,n5378);
    nor g4654(n1151 ,n1100 ,n1032);
    nor g4655(n4325 ,n4213 ,n4087);
    not g4656(n748 ,n1877);
    nor g4657(n3199 ,n3108 ,n3150);
    nor g4658(n1563 ,n711 ,n1106);
    nor g4659(n7576 ,n7343 ,n7477);
    nor g4660(n3043 ,n3012 ,n3041);
    nor g4661(n6754 ,n6584 ,n6678);
    xor g4662(n7726 ,n3453 ,n3451);
    nor g4663(n4658 ,n4539 ,n4596);
    nor g4664(n2080 ,n1988 ,n2060);
    or g4665(n5537 ,n5101 ,n5104);
    xnor g4666(n567 ,n530 ,n516);
    not g4667(n3615 ,n7812);
    not g4668(n4708 ,n4707);
    nor g4669(n386 ,n323 ,n349);
    nor g4670(n3241 ,n3084 ,n3190);
    not g4671(n2996 ,n40[12]);
    xnor g4672(n6414 ,n6086 ,n6076);
    not g4673(n2661 ,n2660);
    xnor g4674(n4538 ,n4396 ,n4208);
    dff g4675(.RN(n1), .SN(1'b1), .CK(n0), .D(n1662), .Q(n10[0]));
    nor g4676(n4130 ,n4012 ,n4007);
    not g4677(n754 ,n1863);
    nor g4678(n5264 ,n5115 ,n5104);
    nor g4679(n4854 ,n4745 ,n4795);
    not g4680(n46 ,n37[0]);
    xnor g4681(n3570 ,n3537 ,n3517);
    nor g4682(n7125 ,n6972 ,n7079);
    nor g4683(n6963 ,n6807 ,n6851);
    nor g4684(n104 ,n25[1] ,n25[0]);
    nor g4685(n5156 ,n5088 ,n5107);
    dff g4686(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[2]), .Q(n15[6]));
    nor g4687(n6249 ,n5738 ,n5934);
    xnor g4688(n5802 ,n5172 ,n5356);
    nor g4689(n5150 ,n5090 ,n5106);
    nor g4690(n2974 ,n2969 ,n2963);
    nor g4691(n6674 ,n6518 ,n6515);
    not g4692(n3630 ,n7790);
    nor g4693(n2192 ,n2028 ,n2131);
    nor g4694(n2261 ,n2179 ,n2238);
    nor g4695(n2869 ,n2821 ,n2846);
    nor g4696(n1307 ,n920 ,n636);
    xnor g4697(n1067 ,n812 ,n674);
    nor g4698(n3110 ,n3013 ,n3029);
    nor g4699(n2846 ,n2814 ,n2807);
    or g4700(n1808 ,n991 ,n1182);
    not g4701(n851 ,n34[2]);
    nor g4702(n1423 ,n946 ,n1101);
    or g4703(n1711 ,n1356 ,n1567);
    not g4704(n3010 ,n40[7]);
    xnor g4705(n4970 ,n4932 ,n4953);
    xnor g4706(n7224 ,n7164 ,n7169);
    nor g4707(n2815 ,n2741 ,n2797);
    xnor g4708(n4857 ,n4783 ,n4744);
    nor g4709(n1529 ,n749 ,n641);
    or g4710(n4260 ,n4018 ,n4028);
    not g4711(n7437 ,n7798);
    nor g4712(n4066 ,n4011 ,n4021);
    nor g4713(n1155 ,n1100 ,n1040);
    nor g4714(n4630 ,n4487 ,n4567);
    xnor g4715(n1060 ,n648 ,n876);
    dff g4716(.RN(n1), .SN(1'b1), .CK(n0), .D(n1699), .Q(n33[2]));
    not g4717(n6703 ,n6702);
    nor g4718(n1175 ,n1106 ,n1080);
    or g4719(n2548 ,n2509 ,n2518);
    nor g4720(n3079 ,n2995 ,n3039);
    nor g4721(n1310 ,n937 ,n636);
    nor g4722(n2647 ,n2533 ,n2616);
    xnor g4723(n7822 ,n3786 ,n3805);
    not g4724(n5285 ,n5284);
    nor g4725(n4505 ,n4344 ,n4424);
    nor g4726(n1308 ,n965 ,n636);
    dff g4727(.RN(n1), .SN(1'b1), .CK(n0), .D(n1687), .Q(n24[12]));
    nor g4728(n179 ,n150 ,n148);
    not g4729(n98 ,n25[0]);
    nor g4730(n3572 ,n3546 ,n3571);
    nor g4731(n7180 ,n7117 ,n7154);
    nor g4732(n2200 ,n2029 ,n2132);
    dff g4733(.RN(n1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n18[2]));
    nor g4734(n1482 ,n756 ,n1099);
    xor g4735(n5762 ,n5320 ,n5410);
    nor g4736(n2920 ,n2863 ,n2897);
    nor g4737(n140 ,n33[5] ,n138);
    nor g4738(n5011 ,n4935 ,n4989);
    nor g4739(n5376 ,n5116 ,n5104);
    not g4740(n4111 ,n4110);
    nor g4741(n4116 ,n4019 ,n4016);
    nor g4742(n4438 ,n4113 ,n4274);
    nor g4743(n5140 ,n5117 ,n5097);
    nor g4744(n6358 ,n6089 ,n6084);
    nor g4745(n2121 ,n1969 ,n2098);
    or g4746(n7654 ,n7578 ,n7536);
    or g4747(n1788 ,n1428 ,n1507);
    nor g4748(n273 ,n159 ,n152);
    nor g4749(n2456 ,n21[4] ,n21[3]);
    not g4750(n3115 ,n3114);
    not g4751(n118 ,n117);
    not g4752(n2836 ,n2835);
    nor g4753(n309 ,n254 ,n228);
    nor g4754(n5080 ,n5079 ,n5069);
    nor g4755(n328 ,n220 ,n282);
    nor g4756(n5595 ,n5216 ,n5192);
    or g4757(n1642 ,n1311 ,n1569);
    nor g4758(n3445 ,n3396 ,n3390);
    nor g4759(n6384 ,n6087 ,n6077);
    nor g4760(n2789 ,n2652 ,n2769);
    xnor g4761(n1959 ,n1940 ,n1921);
    not g4762(n7346 ,n7804);
    nor g4763(n1180 ,n1106 ,n1098);
    xnor g4764(n2786 ,n2725 ,n2633);
    nor g4765(n1285 ,n905 ,n638);
    xnor g4766(n473 ,n409 ,n437);
    xor g4767(n6409 ,n6167 ,n6267);
    xnor g4768(n1038 ,n884 ,n668);
    not g4769(n7411 ,n7783);
    nor g4770(n4478 ,n4320 ,n4432);
    nor g4771(n5446 ,n5115 ,n5106);
    nor g4772(n5067 ,n5044 ,n5052);
    xnor g4773(n5001 ,n4956 ,n4954);
    not g4774(n714 ,n28[10]);
    nor g4775(n7187 ,n7037 ,n7155);
    nor g4776(n2321 ,n2250 ,n2293);
    or g4777(n978 ,n27[3] ,n27[4]);
    nor g4778(n2399 ,n2363 ,n2384);
    not g4779(n4083 ,n4082);
    nor g4780(n4647 ,n4459 ,n4558);
    not g4781(n891 ,n16[8]);
    not g4782(n832 ,n34[1]);
    or g4783(n7632 ,n7530 ,n7545);
    nor g4784(n211 ,n154 ,n148);
    nor g4785(n5854 ,n5349 ,n5623);
    nor g4786(n4152 ,n4020 ,n4025);
    nor g4787(n5486 ,n5088 ,n5104);
    nor g4788(n6836 ,n6611 ,n6724);
    not g4789(n7341 ,n39[2]);
    not g4790(n3121 ,n3120);
    or g4791(n1765 ,n1405 ,n1497);
    nor g4792(n5450 ,n5114 ,n5090);
    not g4793(n4730 ,n4729);
    xor g4794(n7731 ,n3566 ,n3575);
    nor g4795(n307 ,n244 ,n238);
    not g4796(n7269 ,n7268);
    dff g4797(.RN(n1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n27[6]));
    nor g4798(n3648 ,n39[14] ,n7815);
    not g4799(n6181 ,n6180);
    xnor g4800(n6507 ,n6291 ,n5984);
    nor g4801(n2494 ,n2471 ,n2467);
    nor g4802(n3188 ,n3013 ,n3064);
    xnor g4803(n7781 ,n4859 ,n4854);
    nor g4804(n4946 ,n4814 ,n4896);
    xnor g4805(n7243 ,n7192 ,n7180);
    xnor g4806(n6265 ,n5777 ,n5214);
    nor g4807(n1542 ,n895 ,n641);
    nor g4808(n2489 ,n2441 ,n2477);
    nor g4809(n4483 ,n4337 ,n4428);
    not g4810(n833 ,n20[2]);
    nor g4811(n5252 ,n5108 ,n5102);
    xnor g4812(n7802 ,n2117 ,n2005);
    xor g4813(n4669 ,n4561 ,n4522);
    xnor g4814(n6543 ,n6295 ,n5986);
    not g4815(n7431 ,n39[13]);
    xnor g4816(n478 ,n407 ,n394);
    nor g4817(n7239 ,n7234 ,n7232);
    not g4818(n671 ,n23[6]);
    not g4819(n432 ,n431);
    nor g4820(n1358 ,n841 ,n637);
    or g4821(n1580 ,n1241 ,n1468);
    nor g4822(n3555 ,n3525 ,n3531);
    not g4823(n4233 ,n4232);
    xor g4824(n7111 ,n7033 ,n7042);
    not g4825(n7380 ,n7774);
    nor g4826(n465 ,n391 ,n415);
    nor g4827(n3183 ,n3013 ,n3069);
    nor g4828(n3703 ,n3662 ,n3683);
    xnor g4829(n7768 ,n3843 ,n3863);
    nor g4830(n1392 ,n706 ,n1101);
    or g4831(n5542 ,n5091 ,n5111);
    nor g4832(n3770 ,n3707 ,n3730);
    nor g4833(n4763 ,n4662 ,n4697);
    or g4834(n5545 ,n5107 ,n5098);
    not g4835(n6908 ,n6907);
    nor g4836(n2336 ,n2225 ,n2314);
    or g4837(n2004 ,n1963 ,n1975);
    not g4838(n2907 ,n2906);
    nor g4839(n6217 ,n5226 ,n6049);
    or g4840(n1688 ,n1326 ,n1127);
    nor g4841(n1911 ,n19[5] ,n20[5]);
    nor g4842(n1913 ,n19[0] ,n20[0]);
    not g4843(n4179 ,n4178);
    nor g4844(n217 ,n156 ,n152);
    xnor g4845(n7779 ,n4348 ,n4670);
    nor g4846(n1131 ,n634 ,n1085);
    xnor g4847(n7260 ,n7218 ,n7204);
    nor g4848(n2302 ,n2258 ,n2283);
    nor g4849(n2412 ,n2390 ,n2411);
    xnor g4850(n2122 ,n1968 ,n2051);
    nor g4851(n3571 ,n3547 ,n3557);
    xnor g4852(n4381 ,n4220 ,n4190);
    nor g4853(n4815 ,n4644 ,n4751);
    xor g4854(n5829 ,n5567 ,n5502);
    xnor g4855(n6078 ,n5806 ,n5180);
    nor g4856(n5466 ,n5095 ,n5104);
    nor g4857(n6893 ,n6834 ,n6792);
    xnor g4858(n6398 ,n6124 ,n5948);
    nor g4859(n4032 ,n4022 ,n4009);
    nor g4860(n4104 ,n4008 ,n4010);
    not g4861(n7347 ,n7794);
    not g4862(n1099 ,n638);
    nor g4863(n324 ,n204 ,n258);
    xnor g4864(n6279 ,n5938 ,n6004);
    nor g4865(n3245 ,n3051 ,n3137);
    nor g4866(n5605 ,n5476 ,n5142);
    nor g4867(n2900 ,n2763 ,n2875);
    nor g4868(n2009 ,n1902 ,n1978);
    xnor g4869(n6171 ,n5814 ,n5264);
    not g4870(n3622 ,n7813);
    dff g4871(.RN(n1), .SN(1'b1), .CK(n0), .D(n1669), .Q(n25[4]));
    not g4872(n6103 ,n6102);
    dff g4873(.RN(n1), .SN(1'b1), .CK(n0), .D(n1646), .Q(n35[15]));
    not g4874(n682 ,n36[15]);
    buf g4875(n14[15], n11[15]);
    not g4876(n650 ,n35[2]);
    nor g4877(n5871 ,n5525 ,n5598);
    or g4878(n7663 ,n7595 ,n7592);
    not g4879(n4019 ,n37[5]);
    not g4880(n162 ,n161);
    not g4881(n7453 ,n7779);
    not g4882(n6117 ,n6116);
    not g4883(n678 ,n28[7]);
    not g4884(n783 ,n1866);
    nor g4885(n359 ,n271 ,n290);
    not g4886(n3598 ,n7782);
    not g4887(n6518 ,n6517);
    nor g4888(n2398 ,n2376 ,n2385);
    xor g4889(n5794 ,n5537 ,n5218);
    not g4890(n5118 ,n22[1]);
    nor g4891(n4776 ,n4680 ,n4723);
    nor g4892(n2007 ,n1894 ,n1982);
    nor g4893(n4310 ,n4161 ,n4171);
    xnor g4894(n1051 ,n653 ,n847);
    nor g4895(n2018 ,n1890 ,n1982);
    nor g4896(n1265 ,n721 ,n636);
    nor g4897(n1995 ,n1902 ,n1974);
    xnor g4898(n1058 ,n660 ,n879);
    nor g4899(n1509 ,n786 ,n639);
    nor g4900(n2754 ,n2684 ,n2713);
    xnor g4901(n2131 ,n1971 ,n2090);
    nor g4902(n5916 ,n5322 ,n5608);
    nor g4903(n7014 ,n6951 ,n6944);
    xnor g4904(n1080 ,n811 ,n661);
    nor g4905(n4339 ,n4057 ,n4153);
    not g4906(n4109 ,n4108);
    nor g4907(n3082 ,n2995 ,n3037);
    xnor g4908(n6118 ,n5793 ,n5366);
    not g4909(n7408 ,n39[6]);
    nor g4910(n4422 ,n4137 ,n4298);
    nor g4911(n1572 ,n687 ,n634);
    not g4912(n5361 ,n5360);
    xnor g4913(n5833 ,n5378 ,n5232);
    nor g4914(n453 ,n317 ,n421);
    nor g4915(n1956 ,n1891 ,n1937);
    not g4916(n3868 ,n7801);
    nor g4917(n3945 ,n7782 ,n38[5]);
    nor g4918(n6385 ,n6097 ,n6075);
    nor g4919(n4508 ,n4336 ,n4447);
    not g4920(n7402 ,n7715);
    nor g4921(n1247 ,n849 ,n640);
    not g4922(n5273 ,n5272);
    nor g4923(n7130 ,n7033 ,n7082);
    xnor g4924(n2317 ,n2268 ,n2204);
    nor g4925(n1256 ,n918 ,n640);
    or g4926(n1800 ,n1437 ,n1513);
    xnor g4927(n1075 ,n24[2] ,n35[2]);
    nor g4928(n4501 ,n4310 ,n4425);
    nor g4929(n6459 ,n6181 ,n6307);
    nor g4930(n5502 ,n5096 ,n5109);
    xor g4931(n6412 ,n6189 ,n6088);
    nor g4932(n1502 ,n764 ,n639);
    not g4933(n877 ,n16[3]);
    or g4934(n7324 ,n7327 ,n26[1]);
    not g4935(n5389 ,n5388);
    dff g4936(.RN(n1), .SN(1'b1), .CK(n0), .D(n1679), .Q(n34[7]));
    nor g4937(n2362 ,n2331 ,n2342);
    nor g4938(n5468 ,n5116 ,n5111);
    nor g4939(n2075 ,n1985 ,n2047);
    dff g4940(.RN(n1), .SN(1'b1), .CK(n0), .D(n1587), .Q(n12[11]));
    nor g4941(n2765 ,n2680 ,n2712);
    xnor g4942(n2507 ,n2485 ,n2482);
    not g4943(n743 ,n1854);
    or g4944(n7644 ,n7577 ,n7555);
    xnor g4945(n1024 ,n36[8] ,n34[8]);
    dff g4946(.RN(n1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n21[3]));
    xor g4947(n2429 ,n2681 ,n2669);
    not g4948(n1894 ,n37[7]);
    not g4949(n3732 ,n3731);
    nor g4950(n3813 ,n3761 ,n3812);
    nor g4951(n5526 ,n5117 ,n5100);
    xnor g4952(n3849 ,n37[3] ,n19[3]);
    nor g4953(n7089 ,n6999 ,n7035);
    nor g4954(n2539 ,n2432 ,n2521);
    not g4955(n3013 ,n7758);
    or g4956(n1802 ,n1207 ,n1451);
    nor g4957(n7051 ,n7017 ,n6930);
    nor g4958(n2179 ,n2146 ,n2149);
    nor g4959(n6026 ,n5703 ,n5893);
    xnor g4960(n4517 ,n4409 ,n4198);
    not g4961(n5965 ,n5964);
    dff g4962(.RN(n1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n27[3]));
    not g4963(n7279 ,n7278);
    not g4964(n2134 ,n2133);
    not g4965(n3165 ,n3164);
    nor g4966(n326 ,n200 ,n262);
    xnor g4967(n2401 ,n2384 ,n2362);
    nor g4968(n3559 ,n3517 ,n3537);
    xor g4969(n4561 ,n4395 ,n4123);
    nor g4970(n4643 ,n4462 ,n4529);
    nor g4971(n1478 ,n732 ,n639);
    nor g4972(n312 ,n194 ,n256);
    nor g4973(n5897 ,n5544 ,n5590);
    nor g4974(n380 ,n314 ,n366);
    nor g4975(n3877 ,n7812 ,n7800);
    not g4976(n692 ,n35[14]);
    nor g4977(n2505 ,n2479 ,n2491);
    nor g4978(n3284 ,n3117 ,n3218);
    nor g4979(n5903 ,n5510 ,n5628);
    xnor g4980(n3429 ,n3323 ,n3367);
    not g4981(n1905 ,n19[1]);
    nor g4982(n5085 ,n5084 ,n5039);
    nor g4983(n4711 ,n4449 ,n4653);
    xnor g4984(n2928 ,n2881 ,n2835);
    nor g4985(n2568 ,n2444 ,n2519);
    not g4986(n3000 ,n40[9]);
    nor g4987(n431 ,n307 ,n372);
    xnor g4988(n2692 ,n2643 ,n2513);
    nor g4989(n1915 ,n19[6] ,n19[5]);
    xor g4990(n6401 ,n6170 ,n6090);
    nor g4991(n446 ,n320 ,n433);
    xor g4992(n5810 ,n5570 ,n5228);
    nor g4993(n5609 ,n5280 ,n5148);
    nor g4994(n2026 ,n1892 ,n1982);
    xnor g4995(n2839 ,n2775 ,n2631);
    xnor g4996(n7721 ,n3790 ,n3813);
    nor g4997(n4623 ,n4524 ,n4522);
    xnor g4998(n618 ,n600 ,n586);
    not g4999(n5337 ,n5336);
    xnor g5000(n4398 ,n4135 ,n4236);
    nor g5001(n3638 ,n7803 ,n7780);
    not g5002(n3711 ,n3710);
    not g5003(n5455 ,n5454);
    nor g5004(n3206 ,n3061 ,n3177);
    not g5005(n936 ,n1837);
    nor g5006(n3310 ,n3203 ,n3221);
    not g5007(n647 ,n36[1]);
    not g5008(n5756 ,n5755);
    not g5009(n2348 ,n2347);
    or g5010(n1735 ,n1375 ,n1188);
    dff g5011(.RN(n1), .SN(1'b1), .CK(n0), .D(n1588), .Q(n19[7]));
    not g5012(n6115 ,n6114);
    nor g5013(n4270 ,n4018 ,n4017);
    nor g5014(n6927 ,n6838 ,n6894);
    nor g5015(n7043 ,n6962 ,n6989);
    xnor g5016(n3387 ,n3324 ,n3227);
    nor g5017(n2452 ,n21[3] ,n22[3]);
    dff g5018(.RN(n1), .SN(1'b1), .CK(n0), .D(n1602), .Q(n19[2]));
    nor g5019(n7672 ,n7467 ,n7489);
    xor g5020(n4394 ,n4263 ,n4054);
    nor g5021(n2411 ,n2389 ,n2410);
    nor g5022(n7531 ,n7332 ,n7481);
    nor g5023(n6040 ,n5583 ,n5898);
    nor g5024(n1481 ,n778 ,n639);
    nor g5025(n2201 ,n2112 ,n2136);
    dff g5026(.RN(n1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n27[4]));
    nor g5027(n5250 ,n5116 ,n5110);
    nor g5028(n2419 ,n2418 ,n2388);
    nor g5029(n6745 ,n6588 ,n6671);
    not g5030(n2479 ,n2478);
    nor g5031(n2174 ,n2114 ,n2126);
    not g5032(n6254 ,n6253);
    not g5033(n4935 ,n4934);
    nor g5034(n387 ,n232 ,n346);
    not g5035(n7398 ,n7773);
    nor g5036(n1322 ,n961 ,n642);
    nor g5037(n2066 ,n1890 ,n2004);
    or g5038(n1828 ,n1824 ,n1817);
    nor g5039(n5132 ,n5108 ,n5119);
    nor g5040(n3690 ,n3607 ,n3643);
    not g5041(n5405 ,n5404);
    nor g5042(n2460 ,n2437 ,n2447);
    not g5043(n1941 ,n1940);
    xnor g5044(n2166 ,n1968 ,n2091);
    not g5045(n7291 ,n7290);
    nor g5046(n4652 ,n4499 ,n4521);
    nor g5047(n2589 ,n2441 ,n2548);
    xor g5048(n5761 ,n5581 ,n5424);
    xnor g5049(n2736 ,n2663 ,n2575);
    nor g5050(n7120 ,n7055 ,n7091);
    not g5051(n5395 ,n5394);
    nor g5052(n5741 ,n5529 ,n5520);
    nor g5053(n7227 ,n7181 ,n7194);
    nor g5054(n5274 ,n5101 ,n5106);
    nor g5055(n6556 ,n6099 ,n6418);
    not g5056(n47 ,n19[0]);
    not g5057(n410 ,n409);
    nor g5058(n7246 ,n7215 ,n7224);
    nor g5059(n1483 ,n783 ,n1099);
    or g5060(n7660 ,n7591 ,n7590);
    xnor g5061(n3897 ,n7799 ,n7811);
    not g5062(n7416 ,n7796);
    nor g5063(n4454 ,n4413 ,n4410);
    not g5064(n5985 ,n5984);
    xnor g5065(n2406 ,n2392 ,n2378);
    not g5066(n716 ,n1841);
    xnor g5067(n6295 ,n6002 ,n5978);
    nor g5068(n4359 ,n4133 ,n4147);
    nor g5069(n4042 ,n4013 ,n4008);
    xnor g5070(n5823 ,n5164 ,n5278);
    nor g5071(n5058 ,n5033 ,n5020);
    xnor g5072(n1050 ,n648 ,n846);
    not g5073(n779 ,n3[3]);
    nor g5074(n171 ,n160 ,n149);
    nor g5075(n4599 ,n4450 ,n4492);
    nor g5076(n3498 ,n3463 ,n3466);
    not g5077(n186 ,n185);
    xnor g5078(n4387 ,n4074 ,n4030);
    nor g5079(n1999 ,n1903 ,n1974);
    not g5080(n4635 ,n4634);
    xnor g5081(n7081 ,n6976 ,n6909);
    nor g5082(n3421 ,n3395 ,n3389);
    xor g5083(n7790 ,n5062 ,n5081);
    xnor g5084(n7218 ,n7159 ,n7175);
    not g5085(n3147 ,n3146);
    xnor g5086(n3457 ,n3381 ,n3365);
    xnor g5087(n6088 ,n5818 ,n5328);
    nor g5088(n6582 ,n6376 ,n6452);
    nor g5089(n2801 ,n2754 ,n2767);
    not g5090(n2101 ,n2100);
    xnor g5091(n4514 ,n4404 ,n4359);
    nor g5092(n1222 ,n816 ,n1105);
    or g5093(n7618 ,n7510 ,n7509);
    nor g5094(n2967 ,n2931 ,n2947);
    xnor g5095(n5844 ,n5579 ,n5559);
    nor g5096(n183 ,n146 ,n157);
    nor g5097(n5855 ,n5321 ,n5643);
    nor g5098(n5992 ,n5678 ,n5875);
    nor g5099(n6471 ,n6204 ,n6324);
    nor g5100(n5136 ,n5102 ,n5100);
    xnor g5101(n2963 ,n2923 ,n2880);
    xnor g5102(n3962 ,n38[6] ,n7783);
    or g5103(n7687 ,n7613 ,n7629);
    nor g5104(n1113 ,n635 ,n1023);
    or g5105(n1695 ,n1345 ,n1459);
    not g5106(n6941 ,n6940);
    xnor g5107(n2224 ,n2167 ,n2102);
    xnor g5108(n6880 ,n6715 ,n6565);
    xnor g5109(n3360 ,n3318 ,n3261);
    nor g5110(n5730 ,n5225 ,n5381);
    nor g5111(n4088 ,n4011 ,n4008);
    nor g5112(n4192 ,n4027 ,n4006);
    not g5113(n350 ,n349);
    or g5114(n5321 ,n5092 ,n5093);
    xor g5115(n6600 ,n6431 ,n6439);
    not g5116(n5413 ,n5412);
    not g5117(n6111 ,n6110);
    nor g5118(n5540 ,n5107 ,n5093);
    nor g5119(n6434 ,n6208 ,n6304);
    or g5120(n36[4] ,n7702 ,n7713);
    nor g5121(n7503 ,n7384 ,n7476);
    xor g5122(n4672 ,n4560 ,n4552);
    not g5123(n5247 ,n5246);
    or g5124(n7704 ,n7664 ,n7662);
    or g5125(n1696 ,n1346 ,n1460);
    nor g5126(n2177 ,n2151 ,n2137);
    nor g5127(n3222 ,n3045 ,n3129);
    xnor g5128(n6261 ,n5811 ,n5462);
    or g5129(n1714 ,n1564 ,n1164);
    or g5130(n1584 ,n1247 ,n1471);
    xnor g5131(n3569 ,n3531 ,n3525);
    xnor g5132(n6296 ,n6018 ,n6053);
    nor g5133(n4841 ,n4766 ,n4805);
    or g5134(n1008 ,n885 ,n917);
    nor g5135(n4798 ,n4707 ,n4754);
    xnor g5136(n2664 ,n2501 ,n2580);
    xnor g5137(n3955 ,n38[2] ,n7779);
    xnor g5138(n6806 ,n6601 ,n6487);
    not g5139(n954 ,n12[15]);
    nor g5140(n6359 ,n5949 ,n6124);
    nor g5141(n4002 ,n3998 ,n4001);
    nor g5142(n4895 ,n4747 ,n4892);
    nor g5143(n167 ,n150 ,n158);
    or g5144(n5582 ,n5101 ,n5105);
    xnor g5145(n7722 ,n3791 ,n3815);
    xnor g5146(n2977 ,n2964 ,n2969);
    nor g5147(n612 ,n574 ,n598);
    nor g5148(n5674 ,n5435 ,n5505);
    nor g5149(n5929 ,n5455 ,n5746);
    nor g5150(n2049 ,n1894 ,n2002);
    xnor g5151(n7139 ,n7036 ,n7104);
    nor g5152(n5656 ,n5366 ,n5376);
    xnor g5153(n611 ,n580 ,n595);
    xnor g5154(n4741 ,n4611 ,n4478);
    nor g5155(n1352 ,n828 ,n637);
    not g5156(n2271 ,n2270);
    nor g5157(n4634 ,n4491 ,n4582);
    or g5158(n5568 ,n5101 ,n5117);
    nor g5159(n2030 ,n1945 ,n2026);
    not g5160(n7375 ,n40[10]);
    xnor g5161(n443 ,n189 ,n378);
    or g5162(n1707 ,n1216 ,n1534);
    dff g5163(.RN(n1), .SN(1'b1), .CK(n0), .D(n1611), .Q(n12[0]));
    nor g5164(n3775 ,n3708 ,n3729);
    or g5165(n1755 ,n1393 ,n1172);
    not g5166(n5943 ,n5942);
    xnor g5167(n5930 ,n5318 ,n5324);
    dff g5168(.RN(n1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n20[7]));
    xnor g5169(n4595 ,n4394 ,n4226);
    nor g5170(n4460 ,n4315 ,n4426);
    nor g5171(n1539 ,n744 ,n641);
    xnor g5172(n3845 ,n37[1] ,n19[1]);
    not g5173(n5287 ,n5286);
    xnor g5174(n7034 ,n6915 ,n6735);
    nor g5175(n7094 ,n6973 ,n7050);
    not g5176(n2187 ,n1887);
    nor g5177(n2814 ,n2755 ,n2799);
    xor g5178(n3452 ,n3388 ,n3417);
    not g5179(n276 ,n275);
    nor g5180(n3272 ,n3202 ,n3220);
    not g5181(n3610 ,n39[0]);
    nor g5182(n7060 ,n6959 ,n7007);
    or g5183(n5323 ,n5093 ,n5113);
    xnor g5184(n6499 ,n6293 ,n6001);
    nor g5185(n6688 ,n6421 ,n6502);
    nor g5186(n368 ,n197 ,n292);
    nor g5187(n108 ,n103 ,n106);
    nor g5188(n4357 ,n4246 ,n4266);
    nor g5189(n1419 ,n878 ,n638);
    not g5190(n886 ,n28[3]);
    nor g5191(n2583 ,n2498 ,n2561);
    xnor g5192(n3958 ,n7786 ,n7771);
    not g5193(n3520 ,n3519);
    xnor g5194(n1574 ,n25[0] ,n641);
    xnor g5195(n1972 ,n1948 ,n1938);
    nor g5196(n6212 ,n5586 ,n6060);
    not g5197(n5181 ,n5180);
    xnor g5198(n7798 ,n7289 ,n7310);
    or g5199(n998 ,n35[5] ,n35[6]);
    or g5200(n1766 ,n1404 ,n1547);
    nor g5201(n1156 ,n1100 ,n1076);
    xnor g5202(n2083 ,n1967 ,n1983);
    not g5203(n2132 ,n2131);
    xnor g5204(n6073 ,n5837 ,n5757);
    xnor g5205(n4392 ,n4152 ,n4056);
    not g5206(n246 ,n245);
    not g5207(n676 ,n36[12]);
    nor g5208(n2745 ,n2665 ,n2722);
    nor g5209(n1291 ,n719 ,n638);
    not g5210(n2344 ,n2343);
    xnor g5211(n3322 ,n3144 ,n3255);
    nor g5212(n1391 ,n931 ,n1101);
    nor g5213(n3158 ,n2994 ,n3066);
    xnor g5214(n2322 ,n2267 ,n2243);
    xnor g5215(n505 ,n440 ,n401);
    xnor g5216(n4770 ,n4684 ,n4690);
    xor g5217(n7740 ,n7779 ,n7802);
    dff g5218(.RN(n1), .SN(1'b1), .CK(n0), .D(n1740), .Q(n30[2]));
    nor g5219(n3055 ,n2994 ,n3037);
    xnor g5220(n2470 ,n2436 ,n21[2]);
    nor g5221(n3974 ,n3945 ,n3973);
    not g5222(n4465 ,n4464);
    nor g5223(n7307 ,n7275 ,n7292);
    not g5224(n2804 ,n2803);
    or g5225(n1083 ,n987 ,n1015);
    dff g5226(.RN(n1), .SN(1'b1), .CK(n0), .D(n1683), .Q(n34[4]));
    xnor g5227(n6735 ,n6490 ,n6391);
    or g5228(n4263 ,n4021 ,n4028);
    xnor g5229(n2139 ,n2071 ,n1970);
    nor g5230(n5917 ,n5521 ,n5587);
    not g5231(n7369 ,n7785);
    nor g5232(n4132 ,n4012 ,n4019);
    nor g5233(n6416 ,n6335 ,n6319);
    nor g5234(n6190 ,n5964 ,n6024);
    nor g5235(n3984 ,n3946 ,n3983);
    or g5236(n1790 ,n1429 ,n1509);
    nor g5237(n5740 ,n5285 ,n5509);
    not g5238(n2152 ,n2151);
    xnor g5239(n1975 ,n1881 ,n1950);
    nor g5240(n2960 ,n2955 ,n2944);
    not g5241(n541 ,n540);
    nor g5242(n1294 ,n923 ,n636);
    or g5243(n5549 ,n5102 ,n5103);
    nor g5244(n4918 ,n4848 ,n4877);
    not g5245(n5223 ,n5222);
    nor g5246(n6959 ,n6876 ,n6863);
    not g5247(n278 ,n277);
    nor g5248(n384 ,n313 ,n365);
    not g5249(n2367 ,n2366);
    xnor g5250(n451 ,n339 ,n393);
    xnor g5251(n7165 ,n7106 ,n7034);
    nor g5252(n2969 ,n2940 ,n2953);
    xnor g5253(n2830 ,n2803 ,n2749);
    or g5254(n1737 ,n1376 ,n1189);
    not g5255(n3698 ,n3697);
    or g5256(n986 ,n9[3] ,n9[2]);
    nor g5257(n5857 ,n5541 ,n5606);
    nor g5258(n7104 ,n6954 ,n7026);
    nor g5259(n2059 ,n1893 ,n2027);
    nor g5260(n4926 ,n4828 ,n4912);
    not g5261(n4217 ,n4216);
    xnor g5262(n5017 ,n4979 ,n4926);
    nor g5263(n1375 ,n966 ,n1105);
    nor g5264(n1869 ,n140 ,n141);
    nor g5265(n4481 ,n4338 ,n4430);
    not g5266(n887 ,n21[7]);
    not g5267(n5205 ,n5204);
    xnor g5268(n1085 ,n658 ,n662);
    nor g5269(n7214 ,n7128 ,n7183);
    xnor g5270(n7810 ,n2394 ,n2410);
    xnor g5271(n2832 ,n2735 ,n2790);
    nor g5272(n374 ,n315 ,n358);
    xnor g5273(n3889 ,n41[7] ,n7808);
    not g5274(n142 ,n141);
    nor g5275(n3080 ,n2995 ,n3032);
    dff g5276(.RN(n1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n12[14]));
    or g5277(n1758 ,n1395 ,n1494);
    nor g5278(n4993 ,n4945 ,n4961);
    xnor g5279(n5782 ,n5140 ,n5122);
    not g5280(n391 ,n390);
    nor g5281(n4202 ,n4027 ,n4022);
    nor g5282(n2716 ,n2576 ,n2662);
    xnor g5283(n3481 ,n3431 ,n3401);
    xnor g5284(n1059 ,n658 ,n880);
    xnor g5285(n3412 ,n3344 ,n3140);
    not g5286(n7425 ,n39[12]);
    dff g5287(.RN(n1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n21[7]));
    nor g5288(n6230 ,n5991 ,n5989);
    xor g5289(n4397 ,n4254 ,n4032);
    xnor g5290(n6545 ,n6297 ,n5946);
    xnor g5291(n4378 ,n4052 ,n4154);
    nor g5292(n2164 ,n2116 ,n2128);
    or g5293(n1667 ,n1218 ,n1149);
    nor g5294(n2301 ,n2118 ,n2282);
    dff g5295(.RN(n1), .SN(1'b1), .CK(n0), .D(n1612), .Q(n1837));
    nor g5296(n2559 ,n2434 ,n2517);
    nor g5297(n2347 ,n2309 ,n2321);
    nor g5298(n1103 ,n808 ,n1016);
    not g5299(n7364 ,n7806);
    not g5300(n4347 ,n4348);
    nor g5301(n390 ,n316 ,n364);
    nor g5302(n4499 ,n4316 ,n4423);
    nor g5303(n6831 ,n6676 ,n6732);
    nor g5304(n4106 ,n4008 ,n4016);
    nor g5305(n3554 ,n3521 ,n3533);
    not g5306(n722 ,n12[5]);
    not g5307(n2226 ,n1888);
    nor g5308(n3144 ,n2994 ,n3069);
    nor g5309(n2283 ,n2249 ,n2246);
    buf g5310(n15[0], n15[4]);
    nor g5311(n2527 ,n2443 ,n2519);
    not g5312(n908 ,n35[11]);
    nor g5313(n6739 ,n6554 ,n6660);
    not g5314(n4252 ,n4251);
    nor g5315(n5858 ,n5569 ,n5600);
    xnor g5316(n7837 ,n3955 ,n3950);
    nor g5317(n1495 ,n789 ,n639);
    not g5318(n4471 ,n4470);
    nor g5319(n1996 ,n1891 ,n1978);
    xnor g5320(n3531 ,n3486 ,n3389);
    nor g5321(n4335 ,n4061 ,n4225);
    nor g5322(n5867 ,n5548 ,n5657);
    xnor g5323(n7217 ,n7167 ,n7179);
    nor g5324(n4204 ,n4022 ,n4024);
    nor g5325(n4713 ,n4568 ,n4615);
    not g5326(n3596 ,n7781);
    nor g5327(n2891 ,n2855 ,n2861);
    nor g5328(n514 ,n394 ,n488);
    nor g5329(n4094 ,n4023 ,n4007);
    nor g5330(n2925 ,n2879 ,n2922);
    nor g5331(n4503 ,n4332 ,n4441);
    not g5332(n5191 ,n5190);
    xnor g5333(n61 ,n37[7] ,n19[7]);
    or g5334(n197 ,n160 ,n155);
    not g5335(n6933 ,n6932);
    or g5336(n1722 ,n1362 ,n1174);
    xnor g5337(n2105 ,n1958 ,n2031);
    nor g5338(n7557 ,n7350 ,n7478);
    xnor g5339(n3669 ,n7814 ,n7791);
    nor g5340(n7112 ,n7046 ,n7096);
    nor g5341(n7257 ,n7227 ,n7250);
    xnor g5342(n480 ,n405 ,n403);
    nor g5343(n231 ,n154 ,n153);
    xnor g5344(n39[10] ,n2971 ,n2983);
    nor g5345(n371 ,n356 ,n370);
    or g5346(n1792 ,n1203 ,n1560);
    xnor g5347(n6858 ,n6712 ,n6549);
    xnor g5348(n6707 ,n6529 ,n6569);
    nor g5349(n1413 ,n850 ,n638);
    nor g5350(n2183 ,n2120 ,n2166);
    nor g5351(n275 ,n147 ,n153);
    nor g5352(n586 ,n556 ,n569);
    nor g5353(n5966 ,n5698 ,n5888);
    dff g5354(.RN(n1), .SN(1'b1), .CK(n0), .D(n1600), .Q(n16[2]));
    nor g5355(n5610 ,n5362 ,n5134);
    nor g5356(n5013 ,n4901 ,n4977);
    xnor g5357(n7066 ,n6936 ,n6992);
    nor g5358(n5630 ,n5188 ,n5146);
    or g5359(n1003 ,n816 ,n654);
    nor g5360(n4303 ,n4210 ,n4182);
    not g5361(n5578 ,n5577);
    nor g5362(n6665 ,n6479 ,n6531);
    nor g5363(n4512 ,n4324 ,n4440);
    xnor g5364(n2156 ,n1970 ,n2074);
    xnor g5365(n7137 ,n7071 ,n7038);
    xnor g5366(n5932 ,n5751 ,n5382);
    nor g5367(n1382 ,n916 ,n1101);
    nor g5368(n4292 ,n4084 ,n4214);
    nor g5369(n4304 ,n4178 ,n4038);
    xnor g5370(n4670 ,n4600 ,n4180);
    xnor g5371(n2726 ,n2511 ,n2650);
    nor g5372(n2790 ,n2673 ,n2737);
    not g5373(n2929 ,n2928);
    not g5374(n5029 ,n5028);
    or g5375(n1841 ,n86 ,n89);
    xnor g5376(n1923 ,n1904 ,n20[1]);
    nor g5377(n3184 ,n3013 ,n3073);
    nor g5378(n3172 ,n2995 ,n3076);
    nor g5379(n310 ,n166 ,n250);
    nor g5380(n5954 ,n5715 ,n5858);
    not g5381(n7365 ,n7802);
    or g5382(n1760 ,n1399 ,n1495);
    xnor g5383(n2465 ,n2446 ,n22[3]);
    nor g5384(n1305 ,n956 ,n636);
    nor g5385(n5354 ,n5091 ,n5110);
    xnor g5386(n545 ,n483 ,n519);
    nor g5387(n177 ,n147 ,n149);
    xnor g5388(n7785 ,n5049 ,n5060);
    not g5389(n7423 ,n7790);
    xnor g5390(n6163 ,n5786 ,n5216);
    not g5391(n3143 ,n3142);
    nor g5392(n4282 ,n4200 ,n4090);
    nor g5393(n2306 ,n2204 ,n2269);
    xnor g5394(n4768 ,n4542 ,n4686);
    xnor g5395(n352 ,n273 ,n263);
    or g5396(n3034 ,n3005 ,n3002);
    not g5397(n5177 ,n5176);
    not g5398(n6268 ,n6267);
    nor g5399(n3779 ,n3720 ,n3750);
    nor g5400(n3660 ,n3619 ,n3617);
    xor g5401(n1863 ,n67 ,n72);
    xnor g5402(n1977 ,n1916 ,n1961);
    xnor g5403(n4377 ,n4162 ,n4034);
    nor g5404(n4575 ,n4398 ,n4505);
    nor g5405(n3798 ,n3755 ,n3797);
    xnor g5406(n522 ,n474 ,n497);
    nor g5407(n5935 ,n5619 ,n5844);
    nor g5408(n5009 ,n4951 ,n4982);
    nor g5409(n5900 ,n5567 ,n5648);
    not g5410(n2104 ,n2103);
    not g5411(n4171 ,n4170);
    not g5412(n5114 ,n37[0]);
    not g5413(n5477 ,n5476);
    not g5414(n6809 ,n6808);
    nor g5415(n510 ,n472 ,n486);
    nor g5416(n2975 ,n2919 ,n2962);
    nor g5417(n163 ,n145 ,n149);
    nor g5418(n3557 ,n3542 ,n3548);
    or g5419(n36[5] ,n7704 ,n7711);
    not g5420(n7354 ,n40[11]);
    nor g5421(n7559 ,n7346 ,n7477);
    nor g5422(n2877 ,n2813 ,n2840);
    nor g5423(n1184 ,n1002 ,n1104);
    xnor g5424(n6862 ,n6718 ,n6658);
    xnor g5425(n397 ,n344 ,n302);
    not g5426(n5041 ,n5040);
    nor g5427(n5910 ,n5303 ,n5655);
    nor g5428(n3137 ,n3012 ,n3068);
    nor g5429(n7023 ,n6764 ,n6948);
    not g5430(n2826 ,n2825);
    not g5431(n3728 ,n3727);
    xnor g5432(n336 ,n227 ,n253);
    not g5433(n4124 ,n4123);
    xnor g5434(n2215 ,n2157 ,n2158);
    nor g5435(n1523 ,n731 ,n641);
    nor g5436(n6749 ,n6481 ,n6696);
    not g5437(n5503 ,n5502);
    nor g5438(n4876 ,n4836 ,n4844);
    nor g5439(n5739 ,n5367 ,n5377);
    nor g5440(n3710 ,n3642 ,n3688);
    not g5441(n812 ,n27[1]);
    nor g5442(n2543 ,n2434 ,n2519);
    nor g5443(n6210 ,n6058 ,n6016);
    not g5444(n4689 ,n4688);
    xnor g5445(n2728 ,n2511 ,n2619);
    nor g5446(n3820 ,n3763 ,n3819);
    nor g5447(n7524 ,n7425 ,n7474);
    nor g5448(n4661 ,n4555 ,n4553);
    xnor g5449(n3665 ,n7816 ,n7760);
    nor g5450(n5358 ,n5112 ,n5105);
    nor g5451(n6581 ,n6375 ,n6451);
    not g5452(n1978 ,n1977);
    or g5453(n1683 ,n1336 ,n1125);
    not g5454(n958 ,n11[13]);
    not g5455(n496 ,n495);
    not g5456(n5231 ,n5230);
    nor g5457(n6211 ,n6020 ,n5970);
    not g5458(n7448 ,n38[5]);
    xnor g5459(n6531 ,n6286 ,n6065);
    nor g5460(n3987 ,n3952 ,n3986);
    nor g5461(n630 ,n590 ,n629);
    nor g5462(n3291 ,n3251 ,n3261);
    xnor g5463(n2394 ,n2366 ,n2347);
    or g5464(n1002 ,n661 ,n826);
    nor g5465(n1538 ,n792 ,n641);
    not g5466(n2707 ,n2706);
    xnor g5467(n3961 ,n38[5] ,n7782);
    nor g5468(n6563 ,n6250 ,n6437);
    nor g5469(n1190 ,n1010 ,n1104);
    xnor g5470(n6601 ,n6432 ,n6269);
    nor g5471(n3419 ,n3280 ,n3368);
    nor g5472(n2586 ,n2433 ,n2547);
    not g5473(n930 ,n11[8]);
    not g5474(n5145 ,n5144);
    nor g5475(n521 ,n509 ,n511);
    nor g5476(n3862 ,n3844 ,n3861);
    not g5477(n5044 ,n5043);
    nor g5478(n3927 ,n3880 ,n3926);
    dff g5479(.RN(n1), .SN(1'b1), .CK(n0), .D(n1723), .Q(n31[4]));
    not g5480(n709 ,n29[0]);
    xor g5481(n544 ,n508 ,n518);
    xnor g5482(n4365 ,n4058 ,n4222);
    not g5483(n813 ,n27[5]);
    nor g5484(n4659 ,n4525 ,n4523);
    not g5485(n5453 ,n5452);
    nor g5486(n2332 ,n2299 ,n2278);
    not g5487(n7363 ,n39[7]);
    xnor g5488(n6290 ,n6046 ,n6057);
    or g5489(n1602 ,n1264 ,n1481);
    nor g5490(n4345 ,n4095 ,n4099);
    nor g5491(n4766 ,n4639 ,n4706);
    or g5492(n7690 ,n7663 ,n7661);
    nor g5493(n3192 ,n3013 ,n3074);
    nor g5494(n6348 ,n5951 ,n6118);
    xor g5495(n5791 ,n5317 ,n5194);
    nor g5496(n1331 ,n969 ,n642);
    not g5497(n4457 ,n4456);
    nor g5498(n2292 ,n2247 ,n2272);
    not g5499(n6051 ,n6050);
    not g5500(n6787 ,n6786);
    nor g5501(n4880 ,n4854 ,n4849);
    not g5502(n6738 ,n6737);
    not g5503(n5752 ,n5751);
    not g5504(n3597 ,n39[14]);
    not g5505(n658 ,n36[4]);
    nor g5506(n3881 ,n3869 ,n3867);
    nor g5507(n3681 ,n3612 ,n3645);
    xnor g5508(n2468 ,n2438 ,n21[7]);
    nor g5509(n548 ,n451 ,n538);
    nor g5510(n1239 ,n857 ,n640);
    not g5511(n601 ,n600);
    nor g5512(n1266 ,n858 ,n640);
    not g5513(n1814 ,n1813);
    nor g5514(n3351 ,n3213 ,n3292);
    not g5515(n523 ,n522);
    nor g5516(n1878 ,n110 ,n111);
    nor g5517(n6024 ,n5679 ,n5923);
    nor g5518(n5282 ,n5101 ,n5111);
    xnor g5519(n1925 ,n19[5] ,n20[5]);
    nor g5520(n3363 ,n3294 ,n3348);
    not g5521(n728 ,n1849);
    xnor g5522(n455 ,n353 ,n383);
    not g5523(n6260 ,n6259);
    nor g5524(n243 ,n154 ,n151);
    not g5525(n4257 ,n4256);
    xor g5526(n2291 ,n2187 ,n2251);
    nor g5527(n7597 ,n7339 ,n7474);
    not g5528(n1896 ,n20[4]);
    nor g5529(n3682 ,n3606 ,n3647);
    not g5530(n3906 ,n3905);
    not g5531(n5415 ,n5414);
    not g5532(n5497 ,n5496);
    xnor g5533(n7237 ,n7107 ,n7205);
    nor g5534(n4893 ,n4886 ,n4869);
    dff g5535(.RN(n1), .SN(1'b1), .CK(n0), .D(n1678), .Q(n34[8]));
    nor g5536(n1547 ,n914 ,n641);
    nor g5537(n6477 ,n6195 ,n6351);
    xnor g5538(n66 ,n37[2] ,n19[2]);
    nor g5539(n6366 ,n6038 ,n6244);
    xnor g5540(n2694 ,n2627 ,n2513);
    nor g5541(n3370 ,n3281 ,n3339);
    xor g5542(n1849 ,n610 ,n620);
    xnor g5543(n2385 ,n2340 ,n2295);
    not g5544(n7080 ,n7079);
    nor g5545(n2229 ,n2079 ,n2190);
    nor g5546(n1205 ,n814 ,n1107);
    nor g5547(n4425 ,n4264 ,n4306);
    nor g5548(n3943 ,n7789 ,n7774);
    not g5549(n2099 ,n2098);
    not g5550(n5433 ,n5432);
    xnor g5551(n4923 ,n4832 ,n4888);
    dff g5552(.RN(n1), .SN(1'b1), .CK(n0), .D(n1586), .Q(n20[0]));
    not g5553(n7078 ,n7077);
    not g5554(n3750 ,n3749);
    nor g5555(n4959 ,n4888 ,n4942);
    nor g5556(n5695 ,n5387 ,n5407);
    nor g5557(n5519 ,n5115 ,n5113);
    xnor g5558(n3511 ,n3455 ,n3433);
    nor g5559(n7191 ,n7131 ,n7151);
    xnor g5560(n6094 ,n5803 ,n5256);
    nor g5561(n1306 ,n713 ,n636);
    not g5562(n7342 ,n7800);
    or g5563(n1001 ,n651 ,n649);
    nor g5564(n7092 ,n6969 ,n7064);
    not g5565(n6578 ,n6577);
    nor g5566(n1135 ,n641 ,n1054);
    xor g5567(n5803 ,n5311 ,n5432);
    nor g5568(n4336 ,n4155 ,n4053);
    not g5569(n3424 ,n3423);
    or g5570(n1825 ,n1463 ,n1820);
    nor g5571(n6672 ,n6498 ,n6571);
    nor g5572(n2184 ,n2134 ,n2147);
    xnor g5573(n2777 ,n2687 ,n2634);
    xnor g5574(n1022 ,n36[10] ,n34[10]);
    or g5575(n1795 ,n1344 ,n1510);
    xnor g5576(n7774 ,n3891 ,n3925);
    not g5577(n5359 ,n5358);
    not g5578(n6083 ,n6082);
    nor g5579(n1997 ,n1891 ,n1980);
    not g5580(n4024 ,n20[5]);
    buf g5581(n14[3], n11[3]);
    not g5582(n656 ,n36[0]);
    not g5583(n5479 ,n5478);
    not g5584(n820 ,n17[4]);
    not g5585(n5342 ,n5341);
    nor g5586(n6195 ,n5990 ,n5988);
    xnor g5587(n485 ,n398 ,n326);
    or g5588(n7614 ,n7496 ,n7495);
    or g5589(n272 ,n146 ,n155);
    nor g5590(n6191 ,n6050 ,n5976);
    nor g5591(n291 ,n167 ,n163);
    not g5592(n2438 ,n22[7]);
    nor g5593(n2529 ,n2442 ,n2519);
    not g5594(n172 ,n171);
    xnor g5595(n6981 ,n6806 ,n6850);
    not g5596(n713 ,n10[13]);
    not g5597(n699 ,n33[4]);
    xnor g5598(n3999 ,n37[3] ,n20[3]);
    nor g5599(n4114 ,n4007 ,n4009);
    xnor g5600(n6779 ,n6626 ,n6577);
    nor g5601(n7607 ,n7338 ,n7478);
    nor g5602(n2643 ,n2541 ,n2589);
    not g5603(n940 ,n25[3]);
    xnor g5604(n6595 ,n6422 ,n6485);
    not g5605(n5971 ,n5970);
    or g5606(n4134 ,n4006 ,n4010);
    xnor g5607(n6497 ,n6300 ,n5996);
    not g5608(n6991 ,n6990);
    nor g5609(n1873 ,n129 ,n128);
    nor g5610(n4709 ,n4579 ,n4621);
    dff g5611(.RN(n1), .SN(1'b1), .CK(n0), .D(n1630), .Q(n11[5]));
    xnor g5612(n4920 ,n4869 ,n4886);
    xnor g5613(n39[2] ,n2779 ,n2731);
    nor g5614(n5617 ,n5490 ,n5420);
    not g5615(n869 ,n31[0]);
    not g5616(n3911 ,n3910);
    xor g5617(n38[7] ,n39[7] ,n7839);
    nor g5618(n6748 ,n6483 ,n6666);
    not g5619(n660 ,n36[2]);
    dff g5620(.RN(n1), .SN(1'b1), .CK(n0), .D(n1623), .Q(n1833));
    or g5621(n1656 ,n1431 ,n1465);
    or g5622(n1603 ,n1271 ,n1488);
    nor g5623(n4261 ,n4012 ,n4006);
    nor g5624(n7523 ,n7383 ,n7479);
    nor g5625(n1498 ,n760 ,n639);
    not g5626(n6091 ,n6090);
    or g5627(n1631 ,n1296 ,n1232);
    xnor g5628(n3383 ,n3321 ,n3142);
    nor g5629(n6463 ,n6174 ,n6359);
    nor g5630(n4700 ,n4548 ,n4629);
    xnor g5631(n4453 ,n4357 ,n4096);
    nor g5632(n7569 ,n7441 ,n7480);
    dff g5633(.RN(n1), .SN(1'b1), .CK(n0), .D(n1591), .Q(n19[6]));
    nor g5634(n7022 ,n6900 ,n6927);
    nor g5635(n2827 ,n2762 ,n2796);
    nor g5636(n5214 ,n5107 ,n5091);
    or g5637(n1709 ,n1217 ,n1535);
    nor g5638(n466 ,n348 ,n401);
    or g5639(n3036 ,n2998 ,n3008);
    xnor g5640(n3668 ,n7788 ,n7811);
    xnor g5641(n6173 ,n5831 ,n5244);
    nor g5642(n6004 ,n5674 ,n5869);
    nor g5643(n6925 ,n6825 ,n6872);
    nor g5644(n2610 ,n2441 ,n2574);
    xnor g5645(n5824 ,n5242 ,n5158);
    not g5646(n4103 ,n4102);
    not g5647(n7714 ,n38[0]);
    not g5648(n2697 ,n2696);
    nor g5649(n7207 ,n7176 ,n7159);
    xnor g5650(n7169 ,n7110 ,n7073);
    xor g5651(n5785 ,n5346 ,n5248);
    xnor g5652(n1064 ,n809 ,n856);
    nor g5653(n4862 ,n4744 ,n4842);
    nor g5654(n6205 ,n6030 ,n6034);
    nor g5655(n3102 ,n3013 ,n3038);
    nor g5656(n1311 ,n949 ,n637);
    not g5657(n4035 ,n4034);
    not g5658(n663 ,n22[1]);
    nor g5659(n7134 ,n7051 ,n7093);
    xnor g5660(n6114 ,n5771 ,n5511);
    not g5661(n3009 ,n7741);
    nor g5662(n3162 ,n2994 ,n3068);
    nor g5663(n2572 ,n2445 ,n2521);
    nor g5664(n2373 ,n2322 ,n2357);
    nor g5665(n3836 ,n37[6] ,n19[6]);
    nor g5666(n2819 ,n2502 ,n2801);
    not g5667(n4592 ,n4591);
    xor g5668(n7742 ,n7804 ,n7781);
    xnor g5669(n4632 ,n4453 ,n4477);
    nor g5670(n3919 ,n3882 ,n3918);
    nor g5671(n6492 ,n6332 ,n6434);
    nor g5672(n3233 ,n3109 ,n3151);
    dff g5673(.RN(n1), .SN(1'b1), .CK(n0), .D(n18[0]), .Q(n15[4]));
    nor g5674(n4446 ,n4115 ,n4299);
    not g5675(n973 ,n12[9]);
    not g5676(n7345 ,n7775);
    xnor g5677(n6404 ,n6102 ,n6257);
    nor g5678(n1935 ,n1904 ,n1917);
    nor g5679(n4326 ,n4079 ,n4101);
    or g5680(n1781 ,n1420 ,n1140);
    nor g5681(n5587 ,n5254 ,n5286);
    not g5682(n145 ,n37[7]);
    not g5683(n2501 ,n2502);
    xnor g5684(n1055 ,n659 ,n865);
    nor g5685(n5063 ,n5045 ,n5060);
    nor g5686(n4306 ,n4160 ,n4170);
    nor g5687(n4355 ,n4139 ,n4111);
    nor g5688(n4212 ,n4029 ,n4021);
    nor g5689(n1517 ,n807 ,n1099);
    not g5690(n192 ,n191);
    not g5691(n6566 ,n6565);
    dff g5692(.RN(n1), .SN(1'b1), .CK(n0), .D(n1722), .Q(n31[5]));
    nor g5693(n6007 ,n5851 ,n5843);
    xnor g5694(n6624 ,n6392 ,n6253);
    xnor g5695(n4818 ,n4754 ,n4707);
    nor g5696(n7466 ,n7330 ,n7334);
    nor g5697(n2955 ,n2905 ,n2936);
    not g5698(n5409 ,n5408);
    nor g5699(n4581 ,n4461 ,n4502);
    not g5700(n696 ,n35[12]);
    not g5701(n6532 ,n6531);
    not g5702(n2970 ,n2969);
    nor g5703(n7588 ,n7377 ,n7479);
    or g5704(n2027 ,n1909 ,n1977);
    dff g5705(.RN(n1), .SN(1'b1), .CK(n0), .D(n1598), .Q(n12[6]));
    xnor g5706(n4896 ,n4822 ,n4792);
    nor g5707(n3371 ,n3306 ,n3356);
    dff g5708(.RN(n1), .SN(1'b1), .CK(n0), .D(n1767), .Q(n22[3]));
    not g5709(n7400 ,n40[0]);
    xnor g5710(n6537 ,n6292 ,n6054);
    xnor g5711(n3565 ,n3527 ,n3515);
    xnor g5712(n1020 ,n36[12] ,n34[12]);
    nor g5713(n6065 ,n5736 ,n5919);
    nor g5714(n6229 ,n5983 ,n5981);
    nor g5715(n5615 ,n5212 ,n5218);
    nor g5716(n4875 ,n4757 ,n4831);
    not g5717(n4167 ,n4166);
    not g5718(n5576 ,n5575);
    nor g5719(n1195 ,n1008 ,n1104);
    not g5720(n1891 ,n37[3]);
    nor g5721(n4774 ,n4526 ,n4739);
    not g5722(n3008 ,n7742);
    or g5723(n982 ,n35[13] ,n35[14]);
    dff g5724(.RN(n1), .SN(1'b1), .CK(n0), .D(n1732), .Q(n30[7]));
    nor g5725(n5594 ,n5222 ,n5274);
    or g5726(n1644 ,n1312 ,n1452);
    xnor g5727(n3483 ,n3397 ,n3437);
    nor g5728(n2064 ,n1902 ,n2027);
    nor g5729(n7492 ,n7405 ,n7479);
    nor g5730(n4298 ,n4192 ,n4218);
    not g5731(n2769 ,n2768);
    nor g5732(n7010 ,n6856 ,n6933);
    not g5733(n5989 ,n5988);
    not g5734(n4976 ,n4975);
    nor g5735(n5160 ,n5099 ,n5093);
    nor g5736(n3239 ,n3049 ,n3167);
    nor g5737(n4917 ,n4845 ,n4880);
    xnor g5738(n6100 ,n5848 ,n5460);
    nor g5739(n1165 ,n1102 ,n1069);
    nor g5740(n7303 ,n7283 ,n7300);
    nor g5741(n3807 ,n3760 ,n3806);
    nor g5742(n2045 ,n1891 ,n2003);
    not g5743(n653 ,n36[3]);
    nor g5744(n2953 ,n2868 ,n2938);
    not g5745(n3833 ,n19[4]);
    nor g5746(n6197 ,n5952 ,n5968);
    nor g5747(n4644 ,n4497 ,n4557);
    nor g5748(n2389 ,n2348 ,n2366);
    xor g5749(n5834 ,n5552 ,n5492);
    nor g5750(n2014 ,n1901 ,n1982);
    xnor g5751(n1071 ,n24[7] ,n35[7]);
    not g5752(n772 ,n1853);
    nor g5753(n1515 ,n755 ,n639);
    or g5754(n1641 ,n1310 ,n1568);
    xnor g5755(n3957 ,n38[3] ,n7780);
    xnor g5756(n1043 ,n872 ,n830);
    nor g5757(n4361 ,n4248 ,n4252);
    dff g5758(.RN(n1), .SN(1'b1), .CK(n0), .D(n1715), .Q(n24[2]));
    xnor g5759(n7770 ,n3888 ,n3917);
    nor g5760(n3469 ,n3451 ,n3422);
    nor g5761(n3216 ,n3055 ,n3128);
    nor g5762(n3307 ,n3144 ,n3256);
    nor g5763(n7546 ,n7412 ,n7479);
    nor g5764(n5598 ,n5232 ,n5378);
    nor g5765(n3644 ,n7804 ,n7781);
    xnor g5766(n7147 ,n7069 ,n6934);
    xnor g5767(n6984 ,n6866 ,n6907);
    not g5768(n6881 ,n6880);
    dff g5769(.RN(n1), .SN(1'b1), .CK(n0), .D(n1608), .Q(n12[2]));
    not g5770(n3828 ,n37[0]);
    nor g5771(n2421 ,n2373 ,n2420);
    nor g5772(n7271 ,n7267 ,n7226);
    not g5773(n3524 ,n3523);
    nor g5774(n7543 ,n7433 ,n7476);
    dff g5775(.RN(n1), .SN(1'b1), .CK(n0), .D(n1604), .Q(n12[4]));
    xnor g5776(n2635 ,n2510 ,n2526);
    not g5777(n781 ,n1876);
    nor g5778(n5686 ,n5203 ,n5469);
    not g5779(n6834 ,n6833);
    xnor g5780(n3727 ,n39[9] ,n3673);
    nor g5781(n6383 ,n6105 ,n6111);
    nor g5782(n221 ,n150 ,n151);
    nor g5783(n4664 ,n4540 ,n4583);
    not g5784(n5104 ,n19[6]);
    not g5785(n5365 ,n5364);
    nor g5786(n5604 ,n5214 ,n5136);
    not g5787(n6799 ,n6798);
    nor g5788(n5292 ,n5118 ,n5110);
    nor g5789(n2017 ,n1891 ,n1982);
    nor g5790(n3875 ,n7803 ,n7795);
    buf g5791(n15[1], n15[5]);
    nor g5792(n7264 ,n7249 ,n7179);
    nor g5793(n1493 ,n766 ,n639);
    nor g5794(n460 ,n388 ,n420);
    xnor g5795(n7202 ,n7140 ,n7149);
    nor g5796(n4805 ,n4738 ,n4725);
    nor g5797(n3142 ,n2994 ,n3071);
    nor g5798(n3949 ,n7778 ,n38[1]);
    nor g5799(n6305 ,n6062 ,n6221);
    not g5800(n4037 ,n4036);
    nor g5801(n1253 ,n973 ,n636);
    xor g5802(n4367 ,n4145 ,n4046);
    nor g5803(n4005 ,n3995 ,n4004);
    nor g5804(n1370 ,n869 ,n1107);
    not g5805(n6043 ,n6042);
    xnor g5806(n6330 ,n5932 ,n6066);
    not g5807(n4720 ,n4719);
    nor g5808(n5073 ,n5046 ,n5063);
    xnor g5809(n7795 ,n6974 ,n6702);
    dff g5810(.RN(n1), .SN(1'b1), .CK(n0), .D(n1734), .Q(n30[6]));
    nor g5811(n56 ,n49 ,n50);
    not g5812(n769 ,n8[1]);
    not g5813(n5512 ,n5511);
    xnor g5814(n7138 ,n7077 ,n7075);
    nor g5815(n5733 ,n5277 ,n5129);
    xnor g5816(n1084 ,n858 ,n823);
    nor g5817(n3547 ,n3479 ,n3514);
    nor g5818(n4274 ,n4212 ,n4086);
    nor g5819(n4969 ,n4943 ,n4954);
    nor g5820(n4509 ,n4327 ,n4420);
    not g5821(n79 ,n78);
    nor g5822(n4322 ,n4227 ,n4055);
    nor g5823(n1510 ,n726 ,n639);
    not g5824(n798 ,n2[1]);
    nor g5825(n5295 ,n5101 ,n5113);
    not g5826(n3415 ,n3414);
    nor g5827(n6952 ,n6905 ,n6865);
    nor g5828(n5398 ,n5116 ,n5105);
    nor g5829(n4826 ,n4597 ,n4776);
    nor g5830(n5946 ,n5718 ,n5857);
    nor g5831(n495 ,n386 ,n460);
    xnor g5832(n6407 ,n6108 ,n6106);
    nor g5833(n2673 ,n2512 ,n2631);
    not g5834(n214 ,n213);
    xnor g5835(n2160 ,n1968 ,n2095);
    dff g5836(.RN(n1), .SN(1'b1), .CK(n0), .D(n1640), .Q(n10[11]));
    xnor g5837(n6070 ,n5843 ,n5448);
    dff g5838(.RN(n1), .SN(1'b1), .CK(n0), .D(n1703), .Q(n24[7]));
    xnor g5839(n2860 ,n2827 ,n2430);
    nor g5840(n5276 ,n5101 ,n5119);
    not g5841(n962 ,n30[6]);
    nor g5842(n1225 ,n652 ,n1105);
    nor g5843(n1336 ,n662 ,n637);
    not g5844(n5094 ,n19[1]);
    xnor g5845(n6278 ,n6024 ,n6055);
    not g5846(n7142 ,n7141);
    not g5847(n3993 ,n20[0]);
    not g5848(n5053 ,n5052);
    nor g5849(n7209 ,n7119 ,n7169);
    not g5850(n5387 ,n5386);
    not g5851(n6041 ,n6040);
    nor g5852(n2403 ,n2353 ,n2397);
    or g5853(n7457 ,n26[2] ,n26[0]);
    nor g5854(n498 ,n425 ,n445);
    not g5855(n5955 ,n5954);
    xnor g5856(n5842 ,n5519 ,n5528);
    xnor g5857(n6144 ,n5802 ,n5844);
    nor g5858(n1229 ,n655 ,n634);
    not g5859(n7393 ,n41[6]);
    not g5860(n3205 ,n3204);
    nor g5861(n4441 ,n4107 ,n4289);
    xnor g5862(n3456 ,n3412 ,n3410);
    nor g5863(n1211 ,n657 ,n1101);
    nor g5864(n5962 ,n5700 ,n5922);
    nor g5865(n5753 ,n5576 ,n5296);
    nor g5866(n383 ,n312 ,n362);
    xnor g5867(n476 ,n429 ,n413);
    nor g5868(n94 ,n92 ,n93);
    nor g5869(n5081 ,n5080 ,n5064);
    nor g5870(n5850 ,n5383 ,n5752);
    nor g5871(n1407 ,n840 ,n640);
    nor g5872(n363 ,n202 ,n296);
    xnor g5873(n3321 ,n3112 ,n3264);
    nor g5874(n237 ,n160 ,n148);
    dff g5875(.RN(n1), .SN(1'b1), .CK(n0), .D(n1677), .Q(n34[9]));
    not g5876(n775 ,n1850);
    not g5877(n7389 ,n7792);
    xnor g5878(n2688 ,n2622 ,n2513);
    xnor g5879(n39[9] ,n2958 ,n2981);
    not g5880(n904 ,n12[3]);
    nor g5881(n1398 ,n953 ,n642);
    nor g5882(n6743 ,n6492 ,n6680);
    not g5883(n4629 ,n4628);
    xnor g5884(n337 ,n163 ,n167);
    nor g5885(n1234 ,n647 ,n634);
    or g5886(n2770 ,n2514 ,n2711);
    nor g5887(n1534 ,n785 ,n641);
    dff g5888(.RN(n1), .SN(1'b1), .CK(n0), .D(n1696), .Q(n33[4]));
    nor g5889(n2760 ,n2719 ,n2693);
    nor g5890(n2023 ,n1894 ,n1976);
    nor g5891(n5492 ,n5102 ,n5097);
    nor g5892(n3489 ,n3444 ,n3459);
    nor g5893(n4280 ,n4166 ,n4068);
    nor g5894(n3772 ,n3723 ,n3737);
    nor g5895(n255 ,n156 ,n155);
    nor g5896(n2044 ,n1902 ,n2003);
    nor g5897(n5958 ,n5707 ,n5902);
    nor g5898(n472 ,n406 ,n403);
    xnor g5899(n2636 ,n2514 ,n2528);
    nor g5900(n4482 ,n4333 ,n4452);
    not g5901(n4835 ,n4834);
    nor g5902(n249 ,n159 ,n149);
    not g5903(n5945 ,n5944);
    or g5904(n1659 ,n1212 ,n1144);
    nor g5905(n3525 ,n3460 ,n3497);
    not g5906(n848 ,n34[11]);
    nor g5907(n5878 ,n5308 ,n5605);
    not g5908(n6133 ,n6132);
    xnor g5909(n4611 ,n4312 ,n4466);
    xnor g5910(n7824 ,n3788 ,n3801);
    not g5911(n747 ,n2[7]);
    or g5912(n1607 ,n1270 ,n1484);
    nor g5913(n1118 ,n635 ,n1052);
    nor g5914(n2372 ,n2323 ,n2356);
    xnor g5915(n5827 ,n5368 ,n5220);
    nor g5916(n1249 ,n903 ,n637);
    not g5917(n3624 ,n7780);
    dff g5918(.RN(n1), .SN(1'b1), .CK(n0), .D(n1645), .Q(n10[6]));
    nor g5919(n7515 ,n7400 ,n7478);
    not g5920(n51 ,n19[4]);
    not g5921(n5566 ,n5565);
    nor g5922(n3198 ,n3120 ,n3152);
    not g5923(n2189 ,n2188);
    nor g5924(n6448 ,n6165 ,n6306);
    nor g5925(n5672 ,n5171 ,n5503);
    xnor g5926(n63 ,n37[1] ,n19[1]);
    nor g5927(n3282 ,n3138 ,n3215);
    nor g5928(n7046 ,n6925 ,n7002);
    nor g5929(n239 ,n145 ,n155);
    nor g5930(n1174 ,n1106 ,n1078);
    xor g5931(n4373 ,n4129 ,n4184);
    nor g5932(n515 ,n467 ,n497);
    nor g5933(n6420 ,n6198 ,n6305);
    xor g5934(n41[12] ,n7301 ,n7316);
    or g5935(n3040 ,n3011 ,n3007);
    not g5936(n5257 ,n5256);
    nor g5937(n6695 ,n6528 ,n6520);
    nor g5938(n7000 ,n6904 ,n6918);
    xor g5939(n38[3] ,n39[3] ,n7843);
    xnor g5940(n1929 ,n1904 ,n19[2]);
    not g5941(n6027 ,n6026);
    nor g5942(n5994 ,n5685 ,n5878);
    nor g5943(n6549 ,n6349 ,n6417);
    xnor g5944(n2395 ,n2365 ,n2368);
    nor g5945(n1544 ,n909 ,n641);
    nor g5946(n3699 ,n3656 ,n3681);
    nor g5947(n5288 ,n5088 ,n5111);
    nor g5948(n4803 ,n4735 ,n4734);
    not g5949(n416 ,n415);
    nor g5950(n467 ,n432 ,n417);
    nor g5951(n2992 ,n2991 ,n2952);
    or g5952(n1822 ,n1518 ,n1818);
    not g5953(n4099 ,n4098);
    not g5954(n4559 ,n4558);
    nor g5955(n3176 ,n2995 ,n3070);
    not g5956(n817 ,n24[3]);
    not g5957(n5139 ,n5138);
    nor g5958(n5853 ,n5454 ,n5745);
    nor g5959(n4567 ,n4472 ,n4486);
    or g5960(n1827 ,n1823 ,n1822);
    nor g5961(n6460 ,n6157 ,n6338);
    xnor g5962(n3376 ,n3325 ,n3342);
    or g5963(n5556 ,n5089 ,n5093);
    not g5964(n7203 ,n7202);
    xnor g5965(n6782 ,n6505 ,n6622);
    not g5966(n4021 ,n37[1]);
    xor g5967(n1851 ,n579 ,n588);
    not g5968(n5201 ,n5200);
    not g5969(n4077 ,n4076);
    nor g5970(n4649 ,n4458 ,n4559);
    nor g5971(n2416 ,n2404 ,n2415);
    nor g5972(n3910 ,n3881 ,n3909);
    xnor g5973(n39[14] ,n2959 ,n2991);
    xnor g5974(n433 ,n355 ,n267);
    xnor g5975(n4972 ,n4928 ,n4882);
    nor g5976(n1459 ,n806 ,n634);
    nor g5977(n2334 ,n2274 ,n2298);
    nor g5978(n1512 ,n730 ,n639);
    nor g5979(n2555 ,n2441 ,n2517);
    nor g5980(n223 ,n146 ,n158);
    nor g5981(n1380 ,n701 ,n1105);
    nor g5982(n6457 ,n6189 ,n6364);
    nor g5983(n3858 ,n3840 ,n3857);
    nor g5984(n2611 ,n2433 ,n2574);
    xnor g5985(n477 ,n411 ,n374);
    xnor g5986(n3891 ,n41[12] ,n7813);
    not g5987(n793 ,n3[0]);
    not g5988(n803 ,n4[4]);
    nor g5989(n4881 ,n4787 ,n4834);
    xnor g5990(n3900 ,n7796 ,n7804);
    not g5991(n587 ,n586);
    xnor g5992(n474 ,n417 ,n431);
    nor g5993(n6949 ,n6802 ,n6853);
    or g5994(n3042 ,n3003 ,n3024);
    or g5995(n3031 ,n3018 ,n3004);
    nor g5996(n2371 ,n2338 ,n2350);
    not g5997(n942 ,n35[15]);
    not g5998(n6421 ,n6420);
    nor g5999(n3941 ,n7791 ,n7776);
    xnor g6000(n2784 ,n2712 ,n2679);
    nor g6001(n5382 ,n5116 ,n5109);
    xnor g6002(n7143 ,n7070 ,n6928);
    not g6003(n3506 ,n3505);
    nor g6004(n7300 ,n7273 ,n7247);
    nor g6005(n5368 ,n5089 ,n5098);
    nor g6006(n4795 ,n4711 ,n4746);
    nor g6007(n6201 ,n6046 ,n6044);
    xor g6008(n1932 ,n20[3] ,n20[4]);
    nor g6009(n2926 ,n2896 ,n2917);
    or g6010(n1613 ,n1279 ,n1487);
    nor g6011(n1876 ,n116 ,n117);
    or g6012(n7621 ,n7511 ,n7499);
    dff g6013(.RN(n1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n28[7]));
    nor g6014(n5026 ,n4991 ,n5005);
    xnor g6015(n4684 ,n4516 ,n4353);
    xnor g6016(n2467 ,n2448 ,n22[5]);
    nor g6017(n7581 ,n7378 ,n7479);
    xor g6018(n40[10] ,n39[11] ,n7829);
    xnor g6019(n2524 ,n2502 ,n2484);
    nor g6020(n7468 ,n7331 ,n7395);
    not g6021(n4987 ,n4986);
    nor g6022(n5591 ,n5398 ,n5472);
    nor g6023(n2390 ,n2347 ,n2367);
    nor g6024(n2043 ,n1903 ,n2004);
    not g6025(n911 ,n28[12]);
    nor g6026(n2893 ,n2428 ,n2867);
    nor g6027(n1807 ,n1200 ,n1199);
    nor g6028(n6943 ,n6726 ,n6849);
    xnor g6029(n2831 ,n2661 ,n2784);
    nor g6030(n1505 ,n735 ,n639);
    not g6031(n6262 ,n6261);
    nor g6032(n2829 ,n2746 ,n2800);
    not g6033(n2357 ,n2356);
    nor g6034(n3842 ,n3826 ,n3830);
    nor g6035(n7001 ,n6943 ,n6953);
    not g6036(n670 ,n34[6]);
    not g6037(n234 ,n233);
    or g6038(n1645 ,n1314 ,n1453);
    nor g6039(n58 ,n43 ,n51);
    nor g6040(n4166 ,n4021 ,n4009);
    xnor g6041(n2133 ,n1971 ,n2094);
    nor g6042(n5158 ,n5118 ,n5117);
    nor g6043(n4214 ,n4007 ,n4025);
    or g6044(n5334 ,n5096 ,n5107);
    nor g6045(n3967 ,n3957 ,n3966);
    not g6046(n2703 ,n2702);
    dff g6047(.RN(n1), .SN(1'b1), .CK(n0), .D(n1674), .Q(n34[12]));
    nor g6048(n2254 ,n2181 ,n2235);
    nor g6049(n1320 ,n705 ,n637);
    nor g6050(n4884 ,n4809 ,n4823);
    xnor g6051(n5018 ,n4934 ,n4988);
    xnor g6052(n2841 ,n2774 ,n2700);
    not g6053(n790 ,n2[2]);
    xor g6054(n7737 ,n3570 ,n3587);
    nor g6055(n3921 ,n3876 ,n3920);
    nor g6056(n6346 ,n6100 ,n6078);
    nor g6057(n7516 ,n7419 ,n7477);
    nor g6058(n1562 ,n972 ,n1106);
    nor g6059(n5000 ,n4900 ,n4978);
    nor g6060(n2532 ,n2433 ,n2521);
    xnor g6061(n2513 ,n2491 ,n2478);
    nor g6062(n3991 ,n3959 ,n3990);
    xnor g6063(n7775 ,n3896 ,n3927);
    nor g6064(n6964 ,n6799 ,n6875);
    or g6065(n1785 ,n1426 ,n1506);
    nor g6066(n4845 ,n4634 ,n4786);
    nor g6067(n7126 ,n7039 ,n7072);
    not g6068(n3932 ,n38[4]);
    nor g6069(n1467 ,n791 ,n639);
    xor g6070(n40[9] ,n39[10] ,n7830);
    nor g6071(n1288 ,n968 ,n637);
    not g6072(n5093 ,n21[7]);
    or g6073(n5546 ,n5119 ,n5116);
    not g6074(n4864 ,n4863);
    xnor g6075(n524 ,n477 ,n485);
    xnor g6076(n6741 ,n6489 ,n6434);
    not g6077(n525 ,n524);
    nor g6078(n4639 ,n4586 ,n4590);
    not g6079(n6937 ,n6936);
    buf g6080(n14[8], n11[8]);
    xnor g6081(n2958 ,n2929 ,n2912);
    or g6082(n1733 ,n1373 ,n1167);
    or g6083(n7679 ,n7603 ,n7671);
    not g6084(n7326 ,n26[0]);
    not g6085(n4063 ,n4062);
    nor g6086(n625 ,n616 ,n624);
    nor g6087(n6192 ,n5986 ,n5978);
    nor g6088(n2459 ,n21[6] ,n21[5]);
    nor g6089(n2542 ,n2432 ,n2523);
    nor g6090(n2580 ,n2497 ,n2554);
    not g6091(n4463 ,n4462);
    not g6092(n3022 ,n40[1]);
    not g6093(n4885 ,n4884);
    not g6094(n4498 ,n4497);
    nor g6095(n6233 ,n6023 ,n5967);
    xnor g6096(n1076 ,n24[1] ,n35[1]);
    nor g6097(n5422 ,n5095 ,n5117);
    not g6098(n5957 ,n5956);
    nor g6099(n269 ,n150 ,n152);
    nor g6100(n2037 ,n1901 ,n2002);
    nor g6101(n599 ,n591 ,n584);
    not g6102(n592 ,n591);
    nor g6103(n7509 ,n7439 ,n7477);
    dff g6104(.RN(n1), .SN(1'b1), .CK(n0), .D(n1694), .Q(n24[10]));
    nor g6105(n4704 ,n4550 ,n4625);
    nor g6106(n3806 ,n3773 ,n3805);
    xnor g6107(n7763 ,n3848 ,n3851);
    xnor g6108(n5771 ,n5488 ,n5422);
    not g6109(n771 ,n1842);
    nor g6110(n6760 ,n6640 ,n6639);
    not g6111(n3852 ,n3851);
    xnor g6112(n2297 ,n2227 ,n2265);
    not g6113(n6472 ,n6471);
    not g6114(n4007 ,n37[2]);
    not g6115(n3411 ,n3410);
    nor g6116(n4182 ,n4018 ,n4009);
    not g6117(n6629 ,n6628);
    xor g6118(n40[1] ,n39[2] ,n7838);
    nor g6119(n1944 ,n1903 ,n1937);
    nor g6120(n7755 ,n3998 ,n3996);
    nor g6121(n2861 ,n2812 ,n2839);
    nor g6122(n3659 ,n3614 ,n3621);
    nor g6123(n5747 ,n5342 ,n5291);
    not g6124(n583 ,n582);
    not g6125(n4031 ,n4030);
    or g6126(n1200 ,n1091 ,n1096);
    xnor g6127(n6658 ,n6393 ,n6136);
    nor g6128(n4582 ,n4507 ,n4485);
    dff g6129(.RN(n1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n28[4]));
    xnor g6130(n4924 ,n4861 ,n4890);
    or g6131(n1183 ,n23[0] ,n1086);
    nor g6132(n7513 ,n7358 ,n7474);
    xnor g6133(n4979 ,n4921 ,n4936);
    nor g6134(n5996 ,n5705 ,n5880);
    nor g6135(n7317 ,n7316 ,n7297);
    xnor g6136(n41[7] ,n7256 ,n7270);
    not g6137(n216 ,n215);
    xnor g6138(n2216 ,n2110 ,n1884);
    not g6139(n4586 ,n4585);
    not g6140(n5283 ,n5282);
    dff g6141(.RN(n1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n26[2]));
    not g6142(n5838 ,n5837);
    or g6143(n1626 ,n1290 ,n1448);
    or g6144(n1595 ,n1257 ,n1121);
    nor g6145(n2641 ,n2544 ,n2601);
    not g6146(n2276 ,n2275);
    nor g6147(n550 ,n507 ,n528);
    not g6148(n7221 ,n7220);
    xnor g6149(n3694 ,n7802 ,n3663);
    not g6150(n2783 ,n2782);
    nor g6151(n7563 ,n7387 ,n7479);
    nor g6152(n7253 ,n7212 ,n7230);
    nor g6153(n2530 ,n2431 ,n2523);
    nor g6154(n2752 ,n2659 ,n2691);
    nor g6155(n4291 ,n4190 ,n4220);
    nor g6156(n7054 ,n7016 ,n6934);
    dff g6157(.RN(n1), .SN(1'b1), .CK(n0), .D(n1708), .Q(n32[4]));
    nor g6158(n7274 ,n7264 ,n7248);
    nor g6159(n1277 ,n955 ,n637);
    nor g6160(n1218 ,n650 ,n1101);
    xnor g6161(n4609 ,n4473 ,n4493);
    xnor g6162(n3673 ,n7810 ,n7787);
    nor g6163(n5254 ,n5101 ,n5092);
    nor g6164(n1348 ,n708 ,n637);
    xnor g6165(n7028 ,n6912 ,n6837);
    nor g6166(n3657 ,n3618 ,n3598);
    nor g6167(n2036 ,n1946 ,n2014);
    xnor g6168(n6076 ,n5799 ,n5186);
    not g6169(n6968 ,n6967);
    nor g6170(n1334 ,n846 ,n637);
    not g6171(n1904 ,n20[2]);
    not g6172(n5088 ,n22[3]);
    nor g6173(n299 ,n193 ,n255);
    nor g6174(n251 ,n159 ,n158);
    nor g6175(n7213 ,n7133 ,n7172);
    or g6176(n5532 ,n5108 ,n5105);
    dff g6177(.RN(n1), .SN(1'b1), .CK(n0), .D(n1752), .Q(n17[4]));
    dff g6178(.RN(n1), .SN(1'b1), .CK(n0), .D(n1731), .Q(n17[6]));
    nor g6179(n3133 ,n3012 ,n3069);
    xnor g6180(n6846 ,n6616 ,n6740);
    nor g6181(n1158 ,n1100 ,n1029);
    nor g6182(n1129 ,n635 ,n1056);
    not g6183(n482 ,n481);
    xnor g6184(n3337 ,n3263 ,n3162);
    nor g6185(n329 ,n276 ,n218);
    buf g6186(n13[3], n10[3]);
    xnor g6187(n2941 ,n2907 ,n2900);
    nor g6188(n6723 ,n6547 ,n6695);
    nor g6189(n1171 ,n1102 ,n1033);
    dff g6190(.RN(n1), .SN(1'b1), .CK(n0), .D(n1709), .Q(n24[4]));
    nor g6191(n5611 ,n5144 ,n5438);
    nor g6192(n5230 ,n5098 ,n5105);
    nor g6193(n320 ,n214 ,n216);
    xnor g6194(n6594 ,n6428 ,n6441);
    dff g6195(.RN(n1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n28[6]));
    nor g6196(n5064 ,n5040 ,n5054);
    not g6197(n2269 ,n2268);
    or g6198(n983 ,n35[0] ,n35[12]);
    xnor g6199(n6161 ,n5807 ,n5498);
    xnor g6200(n3533 ,n3483 ,n3399);
    not g6201(n720 ,n19[0]);
    xor g6202(n5811 ,n5549 ,n5210);
    not g6203(n6105 ,n6104);
    or g6204(n1643 ,n1313 ,n1570);
    not g6205(n928 ,n19[3]);
    not g6206(n5089 ,n37[2]);
    not g6207(n868 ,n16[1]);
    or g6208(n1651 ,n1323 ,n1552);
    not g6209(n5036 ,n5035);
    xnor g6210(n4922 ,n4787 ,n4889);
    not g6211(n6498 ,n6497);
    or g6212(n1647 ,n1316 ,n1450);
    xnor g6213(n2698 ,n2638 ,n2513);
    nor g6214(n4323 ,n4067 ,n4077);
    xor g6215(n7760 ,n4971 ,n5087);
    nor g6216(n1857 ,n146 ,n152);
    not g6217(n3538 ,n3537);
    nor g6218(n3302 ,n3161 ,n3245);
    not g6219(n3607 ,n39[6]);
    not g6220(n5947 ,n5946);
    nor g6221(n1125 ,n635 ,n1059);
    xnor g6222(n3676 ,n7813 ,n7790);
    buf g6223(n13[4], n11[4]);
    xnor g6224(n6998 ,n6847 ,n6794);
    nor g6225(n1383 ,n838 ,n1103);
    not g6226(n7035 ,n7034);
    xnor g6227(n7162 ,n7099 ,n7134);
    nor g6228(n1820 ,n1102 ,n1814);
    nor g6229(n5622 ,n5208 ,n5426);
    not g6230(n5131 ,n5130);
    xnor g6231(n7109 ,n7030 ,n7044);
    not g6232(n6258 ,n6257);
    or g6233(n1937 ,n1921 ,n1913);
    nor g6234(n2031 ,n1955 ,n2018);
    nor g6235(n7002 ,n6883 ,n6965);
    not g6236(n7419 ,n7809);
    nor g6237(n4279 ,n4150 ,n4270);
    nor g6238(n1149 ,n1100 ,n1026);
    xnor g6239(n4613 ,n4483 ,n4503);
    nor g6240(n4468 ,n4330 ,n4427);
    nor g6241(n4640 ,n4538 ,n4595);
    nor g6242(n1209 ,n818 ,n642);
    nor g6243(n1280 ,n941 ,n637);
    or g6244(n1723 ,n1363 ,n1179);
    nor g6245(n7181 ,n7097 ,n7145);
    nor g6246(n6886 ,n6836 ,n6765);
    nor g6247(n7319 ,n7296 ,n7318);
    nor g6248(n5260 ,n5118 ,n5099);
    nor g6249(n2475 ,n2448 ,n2459);
    nor g6250(n5926 ,n5551 ,n5618);
    xor g6251(n5813 ,n5538 ,n5434);
    dff g6252(.RN(n1), .SN(1'b1), .CK(n0), .D(n1596), .Q(n16[3]));
    nor g6253(n1255 ,n947 ,n637);
    nor g6254(n6988 ,n6961 ,n6942);
    nor g6255(n3705 ,n3651 ,n3684);
    nor g6256(n5144 ,n5107 ,n5103);
    nor g6257(n3046 ,n2994 ,n3032);
    nor g6258(n1916 ,n19[7] ,n20[7]);
    or g6259(n7616 ,n7498 ,n7493);
    nor g6260(n5948 ,n5670 ,n5907);
    nor g6261(n5984 ,n5686 ,n5859);
    not g6262(n725 ,n33[7]);
    xnor g6263(n2924 ,n2887 ,n2825);
    xnor g6264(n2359 ,n2326 ,n2224);
    nor g6265(n2230 ,n2168 ,n2197);
    not g6266(n943 ,n10[1]);
    nor g6267(n6973 ,n6820 ,n6890);
    nor g6268(n1108 ,n922 ,n642);
    not g6269(n777 ,n1855);
    or g6270(n7661 ,n7602 ,n7586);
    nor g6271(n6376 ,n6129 ,n6127);
    nor g6272(n3503 ,n3447 ,n3469);
    not g6273(n6184 ,n6183);
    nor g6274(n2016 ,n1902 ,n1982);
    nor g6275(n4799 ,n4685 ,n4717);
    xnor g6276(n2324 ,n2209 ,n2287);
    nor g6277(n5880 ,n5555 ,n5627);
    not g6278(n2365 ,n2364);
    nor g6279(n3058 ,n3012 ,n3040);
    nor g6280(n4844 ,n4727 ,n4790);
    not g6281(n3825 ,n37[4]);
    nor g6282(n1217 ,n646 ,n642);
    or g6283(n5309 ,n5092 ,n5097);
    nor g6284(n2176 ,n1958 ,n2160);
    xnor g6285(n4364 ,n4076 ,n4066);
    nor g6286(n5380 ,n5100 ,n5094);
    not g6287(n774 ,n5[2]);
    nor g6288(n1132 ,n639 ,n1094);
    not g6289(n6538 ,n6537);
    nor g6290(n5944 ,n5663 ,n5855);
    nor g6291(n1500 ,n805 ,n1099);
    xnor g6292(n4721 ,n4604 ,n4481);
    nor g6293(n7297 ,n7279 ,n7277);
    nor g6294(n5478 ,n5092 ,n5091);
    nor g6295(n3720 ,n3654 ,n3690);
    not g6296(n3592 ,n7803);
    nor g6297(n4990 ,n4947 ,n4964);
    not g6298(n764 ,n5[7]);
    not g6299(n97 ,n25[6]);
    or g6300(n1636 ,n1304 ,n1571);
    nor g6301(n4638 ,n4508 ,n4573);
    xnor g6302(n3070 ,n40[12] ,n7751);
    nor g6303(n1196 ,n1011 ,n1104);
    nor g6304(n3234 ,n3121 ,n3153);
    not g6305(n236 ,n235);
    xnor g6306(n6852 ,n6722 ,n6517);
    xnor g6307(n6098 ,n5821 ,n5332);
    xnor g6308(n2720 ,n2511 ,n2621);
    nor g6309(n5059 ,n5034 ,n5019);
    nor g6310(n4891 ,n4803 ,n4829);
    nor g6311(n3577 ,n3556 ,n3576);
    not g6312(n7146 ,n7145);
    or g6313(n981 ,n35[9] ,n35[10]);
    xnor g6314(n6156 ,n5824 ,n5301);
    nor g6315(n4953 ,n4878 ,n4914);
    not g6316(n6119 ,n6118);
    nor g6317(n1488 ,n797 ,n639);
    not g6318(n3730 ,n3729);
    nor g6319(n6951 ,n6906 ,n6864);
    nor g6320(n5012 ,n4925 ,n4985);
    nor g6321(n3287 ,n3102 ,n3250);
    not g6322(n860 ,n21[4]);
    not g6323(n2150 ,n2149);
    not g6324(n6857 ,n6856);
    nor g6325(n5894 ,n5311 ,n5597);
    nor g6326(n6751 ,n6586 ,n6683);
    nor g6327(n6200 ,n5958 ,n5962);
    not g6328(n898 ,n12[2]);
    xnor g6329(n2227 ,n2160 ,n1959);
    xnor g6330(n2478 ,n21[5] ,n22[5]);
    not g6331(n3396 ,n3395);
    nor g6332(n6238 ,n6047 ,n6045);
    nor g6333(n80 ,n62 ,n79);
    nor g6334(n3305 ,n3107 ,n3257);
    xnor g6335(n2511 ,n2490 ,n2469);
    nor g6336(n6487 ,n6211 ,n6344);
    not g6337(n7378 ,n7782);
    nor g6338(n5925 ,n5298 ,n5638);
    not g6339(n4157 ,n4156);
    nor g6340(n73 ,n67 ,n72);
    not g6341(n248 ,n247);
    xnor g6342(n6638 ,n6402 ,n6275);
    not g6343(n945 ,n35[10]);
    buf g6344(n37[3] ,n1834);
    xnor g6345(n4395 ,n4156 ,n4036);
    nor g6346(n5498 ,n5108 ,n5107);
    or g6347(n1762 ,n1400 ,n1544);
    nor g6348(n185 ,n159 ,n151);
    nor g6349(n3811 ,n3754 ,n3810);
    xor g6350(n7725 ,n3377 ,n3314);
    not g6351(n946 ,n35[8]);
    nor g6352(n7132 ,n7056 ,n7090);
    not g6353(n799 ,n5[5]);
    not g6354(n5489 ,n5488);
    nor g6355(n5550 ,n5114 ,n5100);
    xnor g6356(n1078 ,n813 ,n816);
    xnor g6357(n564 ,n451 ,n538);
    nor g6358(n2990 ,n2989 ,n2966);
    nor g6359(n4289 ,n4202 ,n4048);
    nor g6360(n5708 ,n5363 ,n5135);
    xor g6361(n6170 ,n5772 ,n5402);
    or g6362(n1842 ,n493 ,n633);
    xnor g6363(n7727 ,n3504 ,n3503);
    xnor g6364(n6942 ,n6781 ,n6810);
    nor g6365(n5657 ,n5506 ,n5138);
    dff g6366(.RN(n1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n29[1]));
    not g6367(n5381 ,n5380);
    not g6368(n3746 ,n3745);
    nor g6369(n4702 ,n4560 ,n4618);
    not g6370(n735 ,n5[4]);
    not g6371(n2446 ,n22[4]);
    dff g6372(.RN(n1), .SN(1'b1), .CK(n0), .D(n1681), .Q(n24[15]));
    not g6373(n3738 ,n3737);
    xnor g6374(n475 ,n304 ,n399);
    nor g6375(n5873 ,n5338 ,n5585);
    nor g6376(n2934 ,n2901 ,n2907);
    nor g6377(n4176 ,n4020 ,n4016);
    nor g6378(n6002 ,n5683 ,n5916);
    nor g6379(n295 ,n245 ,n173);
    nor g6380(n7044 ,n6923 ,n7006);
    nor g6381(n6734 ,n6550 ,n6689);
    xnor g6382(n565 ,n501 ,n522);
    not g6383(n4139 ,n4138);
    nor g6384(n6458 ,n6170 ,n6336);
    xor g6385(n7736 ,n3549 ,n3585);
    dff g6386(.RN(n1), .SN(1'b1), .CK(n0), .D(n1718), .Q(n24[1]));
    nor g6387(n2794 ,n2652 ,n2747);
    nor g6388(n7602 ,n7373 ,n7479);
    not g6389(n7374 ,n7738);
    or g6390(n1657 ,n1423 ,n1556);
    xnor g6391(n3068 ,n40[2] ,n7741);
    nor g6392(n2722 ,n2669 ,n2682);
    nor g6393(n7538 ,n7347 ,n7481);
    xnor g6394(n3539 ,n3485 ,n3449);
    not g6395(n7133 ,n7132);
    not g6396(n903 ,n12[11]);
    not g6397(n553 ,n552);
    not g6398(n838 ,n23[3]);
    nor g6399(n4617 ,n4481 ,n4566);
    nor g6400(n2818 ,n2750 ,n2804);
    nor g6401(n7150 ,n7045 ,n7121);
    nor g6402(n1327 ,n926 ,n642);
    not g6403(n6633 ,n6632);
    nor g6404(n3904 ,n3895 ,n3903);
    not g6405(n5159 ,n5158);
    not g6406(n3388 ,n3387);
    not g6407(n6240 ,n6239);
    nor g6408(n6022 ,n5702 ,n5890);
    nor g6409(n5638 ,n5258 ,n5418);
    xnor g6410(n3513 ,n3456 ,n3435);
    xnor g6411(n6788 ,n6603 ,n6511);
    nor g6412(n3132 ,n3012 ,n3066);
    xnor g6413(n4587 ,n4392 ,n4143);
    xnor g6414(n6870 ,n6708 ,n6543);
    nor g6415(n3976 ,n3948 ,n3975);
    xnor g6416(n2107 ,n1959 ,n2035);
    nor g6417(n5922 ,n5552 ,n5660);
    or g6418(n990 ,n17[2] ,n17[3]);
    nor g6419(n1232 ,n658 ,n634);
    not g6420(n454 ,n453);
    not g6421(n4728 ,n4727);
    nor g6422(n6810 ,n6605 ,n6753);
    xnor g6423(n2326 ,n2279 ,n2253);
    not g6424(n6025 ,n6024);
    not g6425(n2451 ,n21[2]);
    nor g6426(n1870 ,n137 ,n138);
    xnor g6427(n6489 ,n6333 ,n6177);
    not g6428(n6520 ,n6519);
    xnor g6429(n6783 ,n6636 ,n6634);
    nor g6430(n3218 ,n3080 ,n3184);
    dff g6431(.RN(n1), .SN(1'b1), .CK(n0), .D(n1634), .Q(n11[1]));
    nor g6432(n3084 ,n2995 ,n3038);
    xnor g6433(n6247 ,n5827 ,n5336);
    nor g6434(n3929 ,n3878 ,n3928);
    dff g6435(.RN(n1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n27[0]));
    not g6436(n677 ,n28[2]);
    xnor g6437(n2883 ,n2832 ,n2789);
    nor g6438(n3083 ,n2995 ,n3033);
    or g6439(n1612 ,n1278 ,n1486);
    or g6440(n7631 ,n7519 ,n7494);
    xnor g6441(n6432 ,n6067 ,n6005);
    xnor g6442(n3066 ,n40[4] ,n7743);
    nor g6443(n3997 ,n37[1] ,n20[1]);
    nor g6444(n6482 ,n6205 ,n6342);
    not g6445(n912 ,n11[10]);
    nor g6446(n2263 ,n2201 ,n2232);
    nor g6447(n1189 ,n1004 ,n1104);
    nor g6448(n3548 ,n3498 ,n3516);
    not g6449(n3935 ,n7781);
    or g6450(n7623 ,n7518 ,n7514);
    nor g6451(n4827 ,n4815 ,n4779);
    nor g6452(n6481 ,n6209 ,n6314);
    nor g6453(n1351 ,n865 ,n1103);
    nor g6454(n562 ,n452 ,n539);
    xnor g6455(n3566 ,n3535 ,n3519);
    buf g6456(n14[5], n10[5]);
    not g6457(n3260 ,n3259);
    nor g6458(n4333 ,n4207 ,n4205);
    or g6459(n92 ,n33[2] ,n33[0]);
    nor g6460(n4348 ,n4151 ,n4271);
    xnor g6461(n2402 ,n2386 ,n2376);
    not g6462(n5572 ,n5571);
    nor g6463(n4232 ,n4029 ,n4008);
    nor g6464(n6003 ,n5665 ,n5927);
    nor g6465(n1858 ,n53 ,n82);
    nor g6466(n6689 ,n6494 ,n6508);
    nor g6467(n7182 ,n7126 ,n7161);
    xnor g6468(n2143 ,n2073 ,n1970);
    nor g6469(n2650 ,n2566 ,n2586);
    nor g6470(n1241 ,n669 ,n640);
    nor g6471(n2987 ,n2961 ,n2986);
    nor g6472(n6438 ,n6200 ,n6302);
    nor g6473(n2251 ,n2177 ,n2234);
    xnor g6474(n2220 ,n2130 ,n2132);
    nor g6475(n1994 ,n1901 ,n1978);
    xnor g6476(n4668 ,n4556 ,n4497);
    nor g6477(n7248 ,n7223 ,n7167);
    nor g6478(n7533 ,n7453 ,n7479);
    nor g6479(n2375 ,n2337 ,n2349);
    or g6480(n1668 ,n1327 ,n1521);
    nor g6481(n3345 ,n3319 ,n3309);
    xnor g6482(n6652 ,n6413 ,n6271);
    nor g6483(n5626 ,n5272 ,n5384);
    nor g6484(n4574 ,n4510 ,n4484);
    nor g6485(n2805 ,n2716 ,n2738);
    nor g6486(n68 ,n57 ,n63);
    or g6487(n1806 ,n1381 ,n1571);
    or g6488(n1627 ,n1292 ,n1229);
    not g6489(n710 ,n12[6]);
    not g6490(n5979 ,n5978);
    not g6491(n648 ,n36[5]);
    nor g6492(n3316 ,n3163 ,n3263);
    nor g6493(n6479 ,n6214 ,n6339);
    nor g6494(n3761 ,n3703 ,n3728);
    not g6495(n2721 ,n2720);
    nor g6496(n4706 ,n4599 ,n4622);
    nor g6497(n4281 ,n4040 ,n4082);
    or g6498(n1682 ,n1334 ,n1126);
    nor g6499(n6896 ,n6833 ,n6793);
    nor g6500(n6445 ,n5994 ,n6352);
    nor g6501(n2400 ,n2377 ,n2386);
    nor g6502(n5654 ,n5122 ,n5140);
    nor g6503(n4419 ,n4128 ,n4280);
    nor g6504(n6312 ,n6114 ,n6112);
    xnor g6505(n4691 ,n4513 ,n4510);
    not g6506(n2521 ,n2520);
    nor g6507(n5164 ,n5097 ,n5113);
    not g6508(n825 ,n24[1]);
    nor g6509(n6946 ,n6841 ,n6892);
    not g6510(n4231 ,n4230);
    nor g6511(n4054 ,n4006 ,n4025);
    nor g6512(n1406 ,n907 ,n642);
    nor g6513(n2648 ,n2539 ,n2602);
    or g6514(n7653 ,n7572 ,n7566);
    nor g6515(n7510 ,n7369 ,n7479);
    nor g6516(n1875 ,n119 ,n120);
    dff g6517(.RN(n1), .SN(1'b1), .CK(n0), .D(n1610), .Q(n1838));
    nor g6518(n3200 ,n3100 ,n3176);
    nor g6519(n4619 ,n4478 ,n4578);
    nor g6520(n5286 ,n5107 ,n5116);
    nor g6521(n1533 ,n738 ,n641);
    xnor g6522(n3888 ,n7797 ,n7809);
    xnor g6523(n2267 ,n2188 ,n2241);
    xnor g6524(n1074 ,n24[3] ,n35[3]);
    not g6525(n262 ,n261);
    nor g6526(n3773 ,n3719 ,n3747);
    nor g6527(n6488 ,n6199 ,n6320);
    nor g6528(n5690 ,n5447 ,n5437);
    not g6529(n6500 ,n6499);
    xnor g6530(n7032 ,n6916 ,n6808);
    nor g6531(n2792 ,n2429 ,n2757);
    not g6532(n727 ,n1843);
    nor g6533(n5896 ,n5547 ,n5593);
    xnor g6534(n3507 ,n3454 ,n3425);
    not g6535(n5443 ,n5442);
    xnor g6536(n6860 ,n6705 ,n6630);
    not g6537(n7223 ,n7222);
    not g6538(n7415 ,n7801);
    nor g6539(n1341 ,n964 ,n1106);
    xnor g6540(n532 ,n479 ,n498);
    or g6541(n7612 ,n7492 ,n7491);
    not g6542(n5187 ,n5186);
    nor g6543(n6683 ,n6544 ,n6541);
    nor g6544(n3368 ,n3300 ,n3357);
    nor g6545(n4433 ,n4134 ,n4297);
    or g6546(n7476 ,n26[0] ,n7323);
    not g6547(n6514 ,n6513);
    xnor g6548(n6289 ,n5743 ,n5956);
    nor g6549(n4044 ,n4020 ,n4017);
    nor g6550(n7606 ,n7410 ,n7475);
    not g6551(n3870 ,n7804);
    nor g6552(n5366 ,n5099 ,n5091);
    nor g6553(n4086 ,n4019 ,n4028);
    not g6554(n4033 ,n4032);
    not g6555(n230 ,n229);
    dff g6556(.RN(n1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n27[1]));
    or g6557(n5320 ,n5099 ,n5103);
    not g6558(n6425 ,n6424);
    nor g6559(n5972 ,n5687 ,n5879);
    nor g6560(n2355 ,n2301 ,n2320);
    not g6561(n730 ,n1859);
    nor g6562(n1518 ,n716 ,n641);
    nor g6563(n4616 ,n4534 ,n4532);
    nor g6564(n6387 ,n6268 ,n6264);
    not g6565(n7178 ,n7177);
    or g6566(n1690 ,n1108 ,n1528);
    nor g6567(n2951 ,n2926 ,n2932);
    not g6568(n7372 ,n7786);
    dff g6569(.RN(n1), .SN(1'b1), .CK(n0), .D(n1663), .Q(n25[7]));
    not g6570(n5399 ,n5398);
    xnor g6571(n3335 ,n3160 ,n3245);
    xnor g6572(n7776 ,n3892 ,n3929);
    or g6573(n1653 ,n1321 ,n1454);
    not g6574(n3338 ,n3337);
    nor g6575(n281 ,n154 ,n152);
    xnor g6576(n6128 ,n5784 ,n5496);
    nor g6577(n6765 ,n6701 ,n6644);
    not g6578(n7061 ,n7060);
    nor g6579(n233 ,n154 ,n158);
    not g6580(n4189 ,n4188);
    nor g6581(n2602 ,n2441 ,n2549);
    nor g6582(n6235 ,n6041 ,n5943);
    xnor g6583(n3336 ,n3146 ,n3247);
    not g6584(n220 ,n219);
    xnor g6585(n3455 ,n3414 ,n3419);
    nor g6586(n169 ,n150 ,n157);
    or g6587(n1622 ,n1287 ,n1446);
    dff g6588(.RN(n1), .SN(1'b1), .CK(n0), .D(n1603), .Q(n16[1]));
    not g6589(n5100 ,n21[3]);
    nor g6590(n2954 ,n2913 ,n2929);
    nor g6591(n7464 ,n41[4] ,n7824);
    nor g6592(n2311 ,n2205 ,n2268);
    not g6593(n7388 ,n7729);
    nor g6594(n6567 ,n6374 ,n6450);
    nor g6595(n135 ,n124 ,n133);
    or g6596(n634 ,n643 ,n1018);
    not g6597(n6859 ,n6858);
    not g6598(n693 ,n26[0]);
    or g6599(n3037 ,n3020 ,n3015);
    nor g6600(n1363 ,n884 ,n1107);
    nor g6601(n4428 ,n4254 ,n4278);
    nor g6602(n620 ,n608 ,n619);
    or g6603(n5308 ,n5100 ,n5109);
    nor g6604(n116 ,n25[5] ,n114);
    xnor g6605(n6395 ,n6114 ,n6112);
    nor g6606(n6341 ,n6142 ,n6138);
    xnor g6607(n6271 ,n5833 ,n5524);
    not g6608(n4175 ,n4174);
    nor g6609(n7769 ,n3835 ,n3864);
    nor g6610(n6239 ,n5664 ,n6008);
    nor g6611(n5694 ,n5273 ,n5385);
    or g6612(n7664 ,n7598 ,n7597);
    not g6613(n3011 ,n40[0]);
    nor g6614(n5688 ,n5211 ,n5463);
    not g6615(n972 ,n30[4]);
    dff g6616(.RN(n1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n28[10]));
    not g6617(n7176 ,n7175);
    nor g6618(n7195 ,n7120 ,n7190);
    xnor g6619(n4861 ,n4779 ,n4815);
    not g6620(n4201 ,n4200);
    not g6621(n3618 ,n7805);
    nor g6622(n4473 ,n4318 ,n4445);
    xnor g6623(n6072 ,n5845 ,n5454);
    nor g6624(n6206 ,n5936 ,n5992);
    nor g6625(n5716 ,n5453 ,n5207);
    xor g6626(n40[2] ,n39[3] ,n7837);
    not g6627(n7328 ,n41[5]);
    xnor g6628(n2109 ,n1958 ,n2036);
    not g6629(n6029 ,n6028);
    not g6630(n5383 ,n5382);
    not g6631(n264 ,n263);
    not g6632(n917 ,n29[3]);
    nor g6633(n6592 ,n6379 ,n6443);
    not g6634(n7339 ,n39[5]);
    xnor g6635(n7839 ,n3889 ,n3915);
    xnor g6636(n1973 ,n1882 ,n1962);
    not g6637(n4027 ,n19[4]);
    nor g6638(n5879 ,n5320 ,n5599);
    not g6639(n7451 ,n7811);
    nor g6640(n5138 ,n5095 ,n5106);
    nor g6641(n5621 ,n5470 ,n5396);
    or g6642(n1649 ,n1318 ,n1456);
    or g6643(n1662 ,n1418 ,n1455);
    not g6644(n3386 ,n3385);
    xnor g6645(n2887 ,n2771 ,n2856);
    nor g6646(n5318 ,n5118 ,n5113);
    not g6647(n685 ,n36[11]);
    or g6648(n1670 ,n1371 ,n1146);
    nor g6649(n6370 ,n6266 ,n6254);
    not g6650(n6179 ,n6178);
    nor g6651(n7548 ,n7340 ,n7479);
    nor g6652(n7460 ,n41[15] ,n7817);
    nor g6653(n3840 ,n3825 ,n3833);
    not g6654(n5509 ,n5508);
    nor g6655(n535 ,n450 ,n504);
    not g6656(n7361 ,n7720);
    or g6657(n7712 ,n7646 ,n7676);
    nor g6658(n5682 ,n5399 ,n5473);
    xnor g6659(n4380 ,n4204 ,n4206);
    nor g6660(n3170 ,n2995 ,n3071);
    not g6661(n6508 ,n6507);
    nor g6662(n3635 ,n7806 ,n7783);
    nor g6663(n6314 ,n6056 ,n6235);
    dff g6664(.RN(n1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n26[0]));
    xnor g6665(n2686 ,n2514 ,n2620);
    nor g6666(n1397 ,n970 ,n1101);
    not g6667(n880 ,n32[4]);
    dff g6668(.RN(n1), .SN(1'b1), .CK(n0), .D(n1698), .Q(n24[9]));
    dff g6669(.RN(n1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n27[2]));
    xnor g6670(n6517 ,n6281 ,n6028);
    buf g6671(n13[9], n10[9]);
    not g6672(n3514 ,n3513);
    not g6673(n2273 ,n2272);
    nor g6674(n4756 ,n4652 ,n4695);
    not g6675(n933 ,n26[1]);
    nor g6676(n5216 ,n5118 ,n5109);
    nor g6677(n6958 ,n6877 ,n6862);
    xnor g6678(n6292 ,n6042 ,n5960);
    nor g6679(n3420 ,n3397 ,n3399);
    nor g6680(n2011 ,n1893 ,n1980);
    nor g6681(n3764 ,n3705 ,n3732);
    xnor g6682(n7025 ,n6856 ,n6932);
    xnor g6683(n6994 ,n6843 ,n6737);
    nor g6684(n2863 ,n2837 ,n2835);
    not g6685(n3831 ,n37[3]);
    xnor g6686(n3670 ,n7815 ,n7792);
    not g6687(n4069 ,n4068);
    not g6688(n5495 ,n5494);
    xnor g6689(n6912 ,n6628 ,n6831);
    nor g6690(n2679 ,n2515 ,n2636);
    nor g6691(n3917 ,n3872 ,n3916);
    xnor g6692(n6614 ,n6414 ,n6335);
    nor g6693(n7267 ,n7244 ,n7173);
    nor g6694(n5976 ,n5668 ,n5864);
    xnor g6695(n7088 ,n6990 ,n6996);
    nor g6696(n1168 ,n1102 ,n1038);
    nor g6697(n1206 ,n812 ,n1107);
    not g6698(n2244 ,n2243);
    dff g6699(.RN(n1), .SN(1'b1), .CK(n0), .D(n1736), .Q(n35[1]));
    nor g6700(n2234 ,n1885 ,n2195);
    not g6701(n2146 ,n2145);
    xnor g6702(n2360 ,n2324 ,n2261);
    not g6703(n6830 ,n6829);
    dff g6704(.RN(n1), .SN(1'b1), .CK(n0), .D(n1713), .Q(n24[3]));
    or g6705(n1787 ,n1425 ,n1198);
    nor g6706(n6965 ,n6826 ,n6873);
    nor g6707(n6956 ,n6788 ,n6881);
    not g6708(n4722 ,n4721);
    xnor g6709(n4973 ,n4919 ,n4904);
    or g6710(n7711 ,n7660 ,n7679);
    not g6711(n4235 ,n4234);
    nor g6712(n2103 ,n2009 ,n2063);
    nor g6713(n4318 ,n4173 ,n4187);
    nor g6714(n3774 ,n3710 ,n3726);
    nor g6715(n5256 ,n5095 ,n5107);
    not g6716(n3609 ,n7792);
    not g6717(n3706 ,n3705);
    not g6718(n7063 ,n7062);
    nor g6719(n540 ,n464 ,n513);
    not g6720(n7446 ,n39[4]);
    not g6721(n5493 ,n5492);
    nor g6722(n5928 ,n5449 ,n5750);
    xnor g6723(n7830 ,n3958 ,n3980);
    xor g6724(n5765 ,n5344 ,n5374);
    dff g6725(.RN(n1), .SN(1'b1), .CK(n0), .D(n1597), .Q(n19[4]));
    xnor g6726(n6854 ,n6721 ,n6741);
    nor g6727(n538 ,n462 ,n512);
    xor g6728(n38[6] ,n39[6] ,n7840);
    not g6729(n5002 ,n5001);
    nor g6730(n492 ,n191 ,n454);
    buf g6731(n14[14], n11[14]);
    not g6732(n1102 ,n1103);
    nor g6733(n3496 ,n3450 ,n3475);
    nor g6734(n1178 ,n1106 ,n1082);
    nor g6735(n4577 ,n4313 ,n4466);
    xnor g6736(n4410 ,n4146 ,n4132);
    nor g6737(n4886 ,n4773 ,n4825);
    xnor g6738(n6808 ,n6593 ,n6436);
    not g6739(n3107 ,n3106);
    nor g6740(n5915 ,n5302 ,n5640);
    nor g6741(n2633 ,n2555 ,n2609);
    nor g6742(n3059 ,n3012 ,n3031);
    or g6743(n3033 ,n3022 ,n3014);
    xnor g6744(n6938 ,n6778 ,n6839);
    xnor g6745(n6068 ,n5839 ,n5755);
    not g6746(n5004 ,n5003);
    xnor g6747(n1063 ,n813 ,n831);
    xnor g6748(n4983 ,n4930 ,n4863);
    nor g6749(n385 ,n303 ,n344);
    nor g6750(n2041 ,n1892 ,n2003);
    nor g6751(n6351 ,n6172 ,n6230);
    nor g6752(n489 ,n384 ,n447);
    nor g6753(n2938 ,n2787 ,n2911);
    nor g6754(n6583 ,n6377 ,n6453);
    dff g6755(.RN(n1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n22[0]));
    dff g6756(.RN(n1), .SN(1'b1), .CK(n0), .D(n1583), .Q(n12[13]));
    xnor g6757(n2153 ,n1971 ,n2072);
    not g6758(n4089 ,n4088);
    not g6759(n701 ,n30[1]);
    nor g6760(n4991 ,n4893 ,n4966);
    not g6761(n3005 ,n40[4]);
    not g6762(n5983 ,n5982);
    nor g6763(n60 ,n44 ,n48);
    not g6764(n7392 ,n41[4]);
    nor g6765(n4653 ,n4415 ,n4601);
    nor g6766(n3156 ,n2994 ,n3073);
    dff g6767(.RN(n1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n28[1]));
    nor g6768(n6473 ,n6202 ,n6357);
    or g6769(n7684 ,n7620 ,n7618);
    not g6770(n5300 ,n5299);
    xnor g6771(n2803 ,n2515 ,n2711);
    nor g6772(n3879 ,n7806 ,n41[5]);
    nor g6773(n3989 ,n3956 ,n3988);
    not g6774(n5319 ,n5318);
    not g6775(n3744 ,n3743);
    xnor g6776(n2908 ,n2859 ,n2833);
    xnor g6777(n6251 ,n5773 ,n5156);
    not g6778(n3867 ,n41[4]);
    not g6779(n6832 ,n6831);
    nor g6780(n4796 ,n4530 ,n4719);
    not g6781(n6613 ,n6612);
    nor g6782(n6835 ,n6604 ,n6734);
    xnor g6783(n1041 ,n875 ,n834);
    dff g6784(.RN(n1), .SN(1'b1), .CK(n0), .D(n1638), .Q(n10[13]));
    nor g6785(n6303 ,n6247 ,n6080);
    nor g6786(n1335 ,n718 ,n642);
    nor g6787(n1567 ,n685 ,n634);
    nor g6788(n5212 ,n5108 ,n5092);
    xnor g6789(n1843 ,n499 ,n632);
    nor g6790(n5851 ,n5448 ,n5749);
    nor g6791(n5919 ,n5331 ,n5635);
    nor g6792(n3166 ,n3012 ,n3072);
    nor g6793(n5244 ,n5097 ,n5106);
    nor g6794(n7514 ,n7420 ,n7477);
    xnor g6795(n2277 ,n2219 ,n2147);
    nor g6796(n191 ,n145 ,n151);
    xnor g6797(n617 ,n602 ,n593);
    nor g6798(n1417 ,n863 ,n638);
    not g6799(n3866 ,n7796);
    nor g6800(n5513 ,n5096 ,n5094);
    or g6801(n36[15] ,n7697 ,n7709);
    nor g6802(n2558 ,n2442 ,n2517);
    nor g6803(n119 ,n25[6] ,n117);
    nor g6804(n7114 ,n7028 ,n7073);
    not g6805(n2434 ,n7763);
    nor g6806(n7048 ,n7023 ,n7008);
    nor g6807(n2062 ,n1892 ,n2027);
    nor g6808(n3856 ,n3838 ,n3855);
    or g6809(n5294 ,n5112 ,n5109);
    nor g6810(n3646 ,n7805 ,n7782);
    nor g6811(n2880 ,n2819 ,n2849);
    nor g6812(n2820 ,n2501 ,n2802);
    nor g6813(n3471 ,n3401 ,n3431);
    nor g6814(n364 ,n278 ,n283);
    nor g6815(n5078 ,n5077 ,n5067);
    nor g6816(n6009 ,n5610 ,n5841);
    not g6817(n7357 ,n7717);
    nor g6818(n2361 ,n2345 ,n2343);
    not g6819(n2844 ,n2843);
    not g6820(n2175 ,n2174);
    dff g6821(.RN(n1), .SN(1'b1), .CK(n0), .D(n1695), .Q(n33[5]));
    xnor g6822(n7803 ,n2216 ,n2170);
    xnor g6823(n2670 ,n2501 ,n2579);
    xnor g6824(n7073 ,n6985 ,n6860);
    xnor g6825(n370 ,n217 ,n275);
    xnor g6826(n6714 ,n6130 ,n6535);
    nor g6827(n4466 ,n4311 ,n4418);
    or g6828(n7643 ,n7501 ,n7553);
    not g6829(n5329 ,n5328);
    not g6830(n4057 ,n4056);
    xnor g6831(n5052 ,n5016 ,n4993);
    not g6832(n2890 ,n2889);
    nor g6833(n5729 ,n5175 ,n5459);
    or g6834(n1650 ,n1298 ,n1551);
    or g6835(n1598 ,n1260 ,n1115);
    not g6836(n5167 ,n5166);
    xnor g6837(n6778 ,n6646 ,n6652);
    nor g6838(n7520 ,n7428 ,n7474);
    not g6839(n4545 ,n4544);
    dff g6840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1660), .Q(n10[2]));
    not g6841(n2006 ,n2005);
    nor g6842(n2414 ,n2396 ,n2413);
    nor g6843(n227 ,n145 ,n158);
    dff g6844(.RN(n1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n33[7]));
    not g6845(n323 ,n322);
    nor g6846(n2896 ,n2788 ,n2866);
    xor g6847(n2424 ,n2453 ,n2471);
    or g6848(n7658 ,n7585 ,n7584);
    nor g6849(n3179 ,n2995 ,n3068);
    nor g6850(n6904 ,n6617 ,n6786);
    not g6851(n4866 ,n4865);
    not g6852(n865 ,n32[6]);
    not g6853(n894 ,n24[12]);
    xor g6854(n6406 ,n6165 ,n6150);
    nor g6855(n7284 ,n7269 ,n7201);
    nor g6856(n4662 ,n4547 ,n4588);
    xnor g6857(n6936 ,n6782 ,n6656);
    nor g6858(n4342 ,n4031 ,n4075);
    nor g6859(n2053 ,n1902 ,n2002);
    not g6860(n2656 ,n2655);
    xnor g6861(n7108 ,n7064 ,n6969);
    xnor g6862(n6868 ,n6716 ,n6531);
    nor g6863(n1281 ,n854 ,n637);
    not g6864(n3252 ,n3251);
    nor g6865(n5755 ,n5574 ,n5516);
    nor g6866(n2652 ,n2558 ,n2607);
    xnor g6867(n7800 ,n7309 ,n7314);
    nor g6868(n3441 ,n3410 ,n3412);
    not g6869(n753 ,n6[5]);
    xnor g6870(n2637 ,n2512 ,n2527);
    nor g6871(n5612 ,n5194 ,n5240);
    dff g6872(.RN(n1), .SN(1'b1), .CK(n0), .D(n1729), .Q(n23[6]));
    xnor g6873(n7255 ,n7173 ,n7226);
    nor g6874(n4690 ,n4577 ,n4619);
    nor g6875(n6729 ,n6438 ,n6673);
    nor g6876(n3776 ,n3721 ,n3749);
    not g6877(n6139 ,n6138);
    xnor g6878(n2658 ,n2502 ,n2583);
    nor g6879(n588 ,n563 ,n568);
    xnor g6880(n1040 ,n886 ,n669);
    buf g6881(n14[12], n11[12]);
    nor g6882(n1166 ,n1102 ,n1039);
    nor g6883(n382 ,n310 ,n363);
    nor g6884(n4426 ,n4103 ,n4304);
    nor g6885(n5075 ,n5074 ,n5058);
    nor g6886(n1550 ,n953 ,n1100);
    not g6887(n6659 ,n6658);
    nor g6888(n3971 ,n3944 ,n3970);
    nor g6889(n5166 ,n5095 ,n5089);
    or g6890(n1757 ,n1396 ,n1542);
    not g6891(n5461 ,n5460);
    or g6892(n1823 ,n1017 ,n1821);
    nor g6893(n4064 ,n4027 ,n4007);
    or g6894(n7325 ,n7391 ,n26[2]);
    nor g6895(n1819 ,n1104 ,n1815);
    or g6896(n1680 ,n1333 ,n1124);
    nor g6897(n1525 ,n752 ,n641);
    nor g6898(n7310 ,n7303 ,n7281);
    nor g6899(n595 ,n560 ,n571);
    nor g6900(n7512 ,n7363 ,n7474);
    nor g6901(n3197 ,n3114 ,n3140);
    nor g6902(n5874 ,n5572 ,n5624);
    nor g6903(n4602 ,n4334 ,n4455);
    nor g6904(n3582 ,n3563 ,n3581);
    nor g6905(n3923 ,n3871 ,n3922);
    nor g6906(n4750 ,n4543 ,n4686);
    xnor g6907(n3504 ,n3465 ,n3463);
    nor g6908(n1347 ,n971 ,n636);
    nor g6909(n5444 ,n5090 ,n5109);
    nor g6910(n245 ,n147 ,n155);
    xnor g6911(n4583 ,n4393 ,n4214);
    nor g6912(n2681 ,n2513 ,n2637);
    nor g6913(n6547 ,n6370 ,n6462);
    nor g6914(n2454 ,n21[7] ,n22[7]);
    not g6915(n702 ,n11[2]);
    nor g6916(n3656 ,n3623 ,n3615);
    nor g6917(n4941 ,n4884 ,n4898);
    xnor g6918(n6980 ,n6864 ,n6905);
    xor g6919(n41[14] ,n7288 ,n7320);
    nor g6920(n6691 ,n6476 ,n6514);
    nor g6921(n5442 ,n5114 ,n5103);
    nor g6922(n4650 ,n4495 ,n4519);
    nor g6923(n82 ,n61 ,n81);
    xnor g6924(n3790 ,n3739 ,n3712);
    nor g6925(n6225 ,n5953 ,n5969);
    not g6926(n7335 ,n7819);
    nor g6927(n3983 ,n3960 ,n3982);
    nor g6928(n6194 ,n5982 ,n5980);
    nor g6929(n4108 ,n4020 ,n4010);
    not g6930(n4494 ,n4493);
    xnor g6931(n2775 ,n2513 ,n2728);
    nor g6932(n7206 ,n7191 ,n7189);
    buf g6933(n14[9], n11[9]);
    xnor g6934(n3323 ,n3156 ,n3216);
    or g6935(n1743 ,n1383 ,n1169);
    not g6936(n2264 ,n2263);
    not g6937(n321 ,n320);
    not g6938(n5574 ,n5573);
    not g6939(n4215 ,n4214);
    nor g6940(n1338 ,n909 ,n642);
    not g6941(n4759 ,n4758);
    nor g6942(n6204 ,n6032 ,n5984);
    dff g6943(.RN(n1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n16[8]));
    not g6944(n872 ,n28[6]);
    not g6945(n5937 ,n5936);
    not g6946(n5465 ,n5464);
    dff g6947(.RN(n1), .SN(1'b1), .CK(n0), .D(n1652), .Q(n35[11]));
    xnor g6948(n62 ,n37[6] ,n19[6]);
    not g6949(n866 ,n16[4]);
    not g6950(n408 ,n407);
    xnor g6951(n6146 ,n5796 ,n5206);
    not g6952(n190 ,n189);
    not g6953(n6097 ,n6096);
    nor g6954(n5032 ,n4968 ,n4996);
    not g6955(n420 ,n419);
    nor g6956(n5872 ,n5293 ,n5646);
    nor g6957(n2577 ,n2499 ,n2570);
    not g6958(n7387 ,n7788);
    dff g6959(.RN(n1), .SN(1'b1), .CK(n0), .D(n1705), .Q(n24[6]));
    xnor g6960(n4906 ,n4819 ,n4766);
    nor g6961(n3408 ,n3297 ,n3364);
    nor g6962(n6389 ,n6014 ,n6210);
    not g6963(n5840 ,n5839);
    nor g6964(n2578 ,n2488 ,n2557);
    nor g6965(n3801 ,n3764 ,n3800);
    dff g6966(.RN(n1), .SN(1'b1), .CK(n0), .D(n1621), .Q(n1834));
    not g6967(n2485 ,n22[0]);
    xnor g6968(n3675 ,n7809 ,n7786);
    dff g6969(.RN(n1), .SN(1'b1), .CK(n0), .D(n1714), .Q(n32[1]));
    not g6970(n7286 ,n7285);
    nor g6971(n4697 ,n4564 ,n4620);
    nor g6972(n1450 ,n846 ,n634);
    nor g6973(n6231 ,n5937 ,n5993);
    xnor g6974(n2382 ,n2344 ,n2345);
    dff g6975(.RN(n1), .SN(1'b1), .CK(n0), .D(n1691), .Q(n33[0]));
    not g6976(n6101 ,n6100);
    not g6977(n1016 ,n1015);
    xnor g6978(n6916 ,n6841 ,n6827);
    nor g6979(n3516 ,n3503 ,n3493);
    not g6980(n5931 ,n5930);
    nor g6981(n3853 ,n3848 ,n3852);
    nor g6982(n4196 ,n4029 ,n4006);
    not g6983(n6506 ,n6505);
    nor g6984(n6052 ,n5731 ,n5913);
    nor g6985(n3583 ,n3558 ,n3582);
    nor g6986(n2645 ,n2572 ,n2615);
    buf g6987(n37[2] ,n1833);
    not g6988(n657 ,n35[7]);
    nor g6989(n3228 ,n3047 ,n3166);
    nor g6990(n6833 ,n6668 ,n6731);
    not g6991(n896 ,n12[1]);
    nor g6992(n5416 ,n5112 ,n5111);
    not g6993(n6099 ,n6098);
    not g6994(n5095 ,n22[4]);
    not g6995(n5758 ,n5757);
    nor g6996(n2917 ,n2870 ,n2893);
    nor g6997(n1447 ,n828 ,n634);
    nor g6998(n1337 ,n847 ,n636);
    not g6999(n5525 ,n5524);
    not g7000(n224 ,n223);
    not g7001(n280 ,n279);
    not g7002(n6877 ,n6876);
    nor g7003(n6367 ,n6095 ,n6245);
    or g7004(n7652 ,n7571 ,n7567);
    not g7005(n4149 ,n4148);
    nor g7006(n3138 ,n2994 ,n3075);
    not g7007(n6801 ,n6800);
    xnor g7008(n2852 ,n2778 ,n2429);
    not g7009(n5129 ,n5128);
    or g7010(n1713 ,n1208 ,n1536);
    buf g7011(n15[2], n15[6]);
    or g7012(n1772 ,n1411 ,n1135);
    not g7013(n5110 ,n19[4]);
    nor g7014(n4949 ,n4833 ,n4907);
    not g7015(n6861 ,n6860);
    dff g7016(.RN(n1), .SN(1'b1), .CK(n0), .D(n1682), .Q(n34[5]));
    nor g7017(n5659 ,n5196 ,n5496);
    xor g7018(n1861 ,n65 ,n76);
    nor g7019(n5553 ,n5108 ,n5110);
    not g7020(n5153 ,n5152);
    nor g7021(n3876 ,n7810 ,n7798);
    nor g7022(n1146 ,n1100 ,n1037);
    xnor g7023(n2270 ,n2210 ,n2174);
    nor g7024(n207 ,n160 ,n152);
    nor g7025(n2309 ,n2221 ,n2271);
    nor g7026(n1230 ,n659 ,n634);
    nor g7027(n1945 ,n1901 ,n1937);
    nor g7028(n2310 ,n2248 ,n2273);
    nor g7029(n1813 ,n992 ,n1692);
    nor g7030(n4511 ,n4340 ,n4417);
    xnor g7031(n6275 ,n5826 ,n5388);
    nor g7032(n4951 ,n4827 ,n4910);
    not g7033(n2519 ,n2518);
    nor g7034(n4849 ,n4635 ,n4785);
    nor g7035(n4677 ,n4511 ,n4657);
    nor g7036(n1238 ,n835 ,n638);
    nor g7037(n1877 ,n113 ,n114);
    not g7038(n681 ,n21[0]);
    nor g7039(n2071 ,n1997 ,n2042);
    nor g7040(n3765 ,n3702 ,n3735);
    nor g7041(n7270 ,n7239 ,n7231);
    xnor g7042(n6800 ,n6600 ,n6509);
    xnor g7043(n6648 ,n6406 ,n6082);
    nor g7044(n6203 ,n6028 ,n6026);
    not g7045(n3740 ,n3739);
    nor g7046(n1424 ,n859 ,n642);
    nor g7047(n4986 ,n4894 ,n4965);
    nor g7048(n5386 ,n5088 ,n5089);
    nor g7049(n3647 ,n39[13] ,n7814);
    nor g7050(n607 ,n596 ,n581);
    nor g7051(n5184 ,n5088 ,n5110);
    nor g7052(n6310 ,n6001 ,n6225);
    not g7053(n750 ,n3[5]);
    xnor g7054(n3431 ,n3328 ,n3363);
    not g7055(n6188 ,n6187);
    xnor g7056(n7809 ,n2382 ,n2408);
    nor g7057(n113 ,n25[4] ,n111);
    not g7058(n759 ,n2[6]);
    xnor g7059(n4675 ,n4538 ,n4595);
    nor g7060(n6611 ,n6430 ,n6509);
    nor g7061(n3093 ,n3012 ,n3034);
    not g7062(n2449 ,n21[3]);
    buf g7063(n13[10], n10[10]);
    xnor g7064(n2700 ,n2649 ,n2513);
    not g7065(n841 ,n34[13]);
    nor g7066(n4663 ,n4541 ,n4584);
    not g7067(n6331 ,n6330);
    not g7068(n5055 ,n5054);
    xor g7069(n6175 ,n5804 ,n5392);
    nor g7070(n4964 ,n4917 ,n4946);
    xnor g7071(n4610 ,n4398 ,n4505);
    not g7072(n6645 ,n6644);
    nor g7073(n6342 ,n6063 ,n6237);
    xnor g7074(n3385 ,n3343 ,n3150);
    not g7075(n2081 ,n2080);
    nor g7076(n5436 ,n5098 ,n5094);
    or g7077(n7630 ,n7531 ,n7527);
    nor g7078(n4752 ,n4664 ,n4692);
    nor g7079(n7228 ,n7198 ,n7147);
    nor g7080(n1445 ,n848 ,n634);
    nor g7081(n6892 ,n6828 ,n6809);
    or g7082(n1638 ,n1306 ,n1565);
    xnor g7083(n6410 ,n6104 ,n6110);
    nor g7084(n426 ,n325 ,n376);
    or g7085(n1182 ,n17[0] ,n1089);
    nor g7086(n547 ,n535 ,n543);
    not g7087(n4786 ,n4785);
    not g7088(n5099 ,n37[7]);
    nor g7089(n3578 ,n3561 ,n3577);
    nor g7090(n5735 ,n5237 ,n5425);
    not g7091(n724 ,n28[15]);
    xnor g7092(n1026 ,n677 ,n833);
    nor g7093(n6468 ,n6166 ,n6346);
    not g7094(n7417 ,n40[12]);
    xnor g7095(n7222 ,n7163 ,n7143);
    nor g7096(n3348 ,n3227 ,n3278);
    not g7097(n3827 ,n37[2]);
    nor g7098(n4247 ,n4012 ,n4020);
    nor g7099(n3347 ,n3228 ,n3304);
    not g7100(n905 ,n1834);
    xnor g7101(n7141 ,n7067 ,n7085);
    nor g7102(n369 ,n212 ,n297);
    nor g7103(n3372 ,n3240 ,n3337);
    nor g7104(n5669 ,n5215 ,n5137);
    nor g7105(n6922 ,n6837 ,n6903);
    not g7106(n2154 ,n2153);
    or g7107(n5317 ,n5119 ,n5100);
    not g7108(n4095 ,n4094);
    nor g7109(n1212 ,n821 ,n1101);
    nor g7110(n560 ,n516 ,n531);
    not g7111(n3721 ,n3720);
    nor g7112(n5877 ,n5317 ,n5612);
    xnor g7113(n4400 ,n4240 ,n4261);
    nor g7114(n5472 ,n5096 ,n5104);
    not g7115(n6536 ,n6535);
    not g7116(n2680 ,n2679);
    xnor g7117(n503 ,n443 ,n438);
    xnor g7118(n7192 ,n7145 ,n7097);
    nor g7119(n88 ,n83 ,n87);
    nor g7120(n2979 ,n2935 ,n2978);
    nor g7121(n2051 ,n1894 ,n2003);
    nor g7122(n1427 ,n888 ,n642);
    not g7123(n3141 ,n3140);
    not g7124(n4782 ,n4781);
    nor g7125(n1246 ,n691 ,n637);
    nor g7126(n4320 ,n4085 ,n4215);
    not g7127(n7359 ,n7816);
    xnor g7128(n2944 ,n2903 ,n2866);
    or g7129(n1620 ,n1286 ,n1445);
    buf g7130(n37[4] ,n1835);
    xor g7131(n5784 ,n5343 ,n5196);
    nor g7132(n1342 ,n942 ,n1101);
    not g7133(n4399 ,n4398);
    nor g7134(n1105 ,n18[2] ,n999);
    dff g7135(.RN(n1), .SN(1'b1), .CK(n0), .D(n1628), .Q(n1831));
    or g7136(n5310 ,n5095 ,n5119);
    xnor g7137(n1056 ,n655 ,n688);
    or g7138(n1752 ,n1223 ,n1194);
    nor g7139(n209 ,n146 ,n149);
    nor g7140(n1946 ,n1893 ,n1937);
    xnor g7141(n6523 ,n6301 ,n6056);
    not g7142(n3590 ,n39[9]);
    nor g7143(n4098 ,n4027 ,n4021);
    not g7144(n1816 ,n1815);
    or g7145(n1093 ,n983 ,n982);
    nor g7146(n551 ,n496 ,n524);
    xnor g7147(n3453 ,n3391 ,n3316);
    nor g7148(n4058 ,n4027 ,n4020);
    not g7149(n2384 ,n2383);
    nor g7150(n1524 ,n771 ,n641);
    nor g7151(n5677 ,n5401 ,n5361);
    not g7152(n751 ,n1862);
    nor g7153(n1145 ,n1100 ,n1025);
    nor g7154(n4030 ,n4014 ,n4022);
    nor g7155(n2260 ,n2241 ,n2188);
    nor g7156(n3226 ,n3081 ,n3192);
    not g7157(n712 ,n19[2]);
    nor g7158(n1176 ,n1106 ,n1081);
    buf g7159(n14[7], n10[7]);
    nor g7160(n4228 ,n4022 ,n4016);
    nor g7161(n2585 ,n2443 ,n2547);
    xor g7162(n7738 ,n3565 ,n3589);
    xnor g7163(n3463 ,n3378 ,n3158);
    not g7164(n883 ,n32[0]);
    or g7165(n1731 ,n1221 ,n1193);
    nor g7166(n1408 ,n934 ,n642);
    not g7167(n5227 ,n5226);
    not g7168(n2450 ,n21[4]);
    xnor g7169(n3749 ,n39[7] ,n3674);
    xnor g7170(n4792 ,n4675 ,n4598);
    xnor g7171(n5072 ,n5054 ,n5040);
    nor g7172(n4449 ,n4181 ,n4347);
    nor g7173(n5280 ,n5114 ,n5093);
    nor g7174(n1221 ,n819 ,n1105);
    not g7175(n5173 ,n5172);
    buf g7176(n13[6], n11[6]);
    nor g7177(n543 ,n491 ,n514);
    xnor g7178(n3794 ,n3729 ,n3707);
    not g7179(n704 ,n26[2]);
    dff g7180(.RN(n1), .SN(1'b1), .CK(n0), .D(n1746), .Q(n29[5]));
    or g7181(n4120 ,n4020 ,n4009);
    nor g7182(n4141 ,n4006 ,n4024);
    not g7183(n815 ,n24[7]);
    xnor g7184(n4607 ,n4468 ,n4511);
    or g7185(n1587 ,n1249 ,n1130);
    not g7186(n238 ,n237);
    xnor g7187(n2392 ,n2359 ,n2313);
    not g7188(n7174 ,n7173);
    not g7189(n6125 ,n6124);
    nor g7190(n1340 ,n635 ,n1062);
    nor g7191(n5870 ,n5323 ,n5650);
    nor g7192(n378 ,n309 ,n361);
    or g7193(n2547 ,n2508 ,n2522);
    xnor g7194(n7220 ,n7162 ,n7165);
    nor g7195(n5616 ,n5236 ,n5424);
    nor g7196(n5528 ,n5115 ,n5114);
    nor g7197(n3352 ,n3212 ,n3293);
    nor g7198(n6380 ,n6103 ,n6258);
    nor g7199(n3214 ,n3093 ,n3194);
    nor g7200(n2797 ,n2730 ,n2756);
    xnor g7201(n2162 ,n1968 ,n2075);
    nor g7202(n3154 ,n2994 ,n3076);
    xor g7203(n7110 ,n7029 ,n7045);
    not g7204(n3861 ,n3860);
    not g7205(n126 ,n33[5]);
    not g7206(n5371 ,n5370);
    nor g7207(n3468 ,n3393 ,n3425);
    nor g7208(n6684 ,n6543 ,n6542);
    not g7209(n4874 ,n4873);
    nor g7210(n4340 ,n4191 ,n4221);
    not g7211(n906 ,n11[6]);
    xnor g7212(n3893 ,n7802 ,n7794);
    nor g7213(n1514 ,n757 ,n639);
    nor g7214(n5901 ,n5351 ,n5642);
    xor g7215(n4390 ,n4255 ,n4186);
    nor g7216(n5891 ,n5333 ,n5611);
    nor g7217(n6755 ,n6659 ,n6686);
    xnor g7218(n4558 ,n4371 ,n4042);
    not g7219(n7244 ,n7243);
    xor g7220(n7752 ,n7814 ,n7791);
    xnor g7221(n67 ,n37[3] ,n19[3]);
    xor g7222(n7729 ,n3552 ,n3571);
    not g7223(n4549 ,n4548);
    xnor g7224(n335 ,n175 ,n235);
    or g7225(n1689 ,n1329 ,n1122);
    or g7226(n36[7] ,n7684 ,n7710);
    nor g7227(n5642 ,n5174 ,n5458);
    nor g7228(n6907 ,n6771 ,n6814);
    not g7229(n176 ,n175);
    not g7230(n70 ,n69);
    nor g7231(n7055 ,n6996 ,n6991);
    nor g7232(n365 ,n294 ,n330);
    or g7233(n36[6] ,n7683 ,n7706);
    nor g7234(n7605 ,n7360 ,n7476);
    or g7235(n1712 ,n1276 ,n1163);
    not g7236(n6079 ,n6078);
    or g7237(n36[11] ,n7682 ,n7690);
    nor g7238(n2484 ,n2443 ,n2477);
    nor g7239(n487 ,n457 ,n444);
    nor g7240(n141 ,n126 ,n139);
    nor g7241(n3841 ,n3827 ,n3824);
    nor g7242(n2076 ,n2021 ,n2064);
    nor g7243(n1139 ,n641 ,n1044);
    nor g7244(n7666 ,n7473 ,n7483);
    not g7245(n4259 ,n4258);
    nor g7246(n2531 ,n2431 ,n2519);
    nor g7247(n5856 ,n5537 ,n5615);
    nor g7248(n3579 ,n3554 ,n3578);
    not g7249(n2785 ,n2784);
    nor g7250(n1160 ,n1102 ,n1063);
    xnor g7251(n6104 ,n5787 ,n5297);
    nor g7252(n574 ,n540 ,n552);
    nor g7253(n1109 ,n635 ,n1042);
    not g7254(n103 ,n25[2]);
    dff g7255(.RN(n1), .SN(1'b1), .CK(n0), .D(n1673), .Q(n25[2]));
    nor g7256(n4966 ,n4913 ,n4939);
    not g7257(n2523 ,n2522);
    not g7258(n873 ,n32[1]);
    nor g7259(n6371 ,n6248 ,n6081);
    nor g7260(n2058 ,n1903 ,n2002);
    nor g7261(n7473 ,n7333 ,n7394);
    nor g7262(n5134 ,n5118 ,n5111);
    not g7263(n3019 ,n40[14]);
    or g7264(n4140 ,n4008 ,n4009);
    nor g7265(n2851 ,n2751 ,n2828);
    nor g7266(n4988 ,n4941 ,n4969);
    xnor g7267(n6798 ,n6598 ,n6513);
    not g7268(n5133 ,n5132);
    nor g7269(n7050 ,n6936 ,n6992);
    xnor g7270(n6178 ,n5761 ,n5236);
    nor g7271(n2492 ,n2461 ,n2473);
    nor g7272(n3544 ,n3492 ,n3512);
    nor g7273(n1376 ,n972 ,n1105);
    nor g7274(n1287 ,n912 ,n637);
    not g7275(n5051 ,n5050);
    nor g7276(n5624 ,n5400 ,n5360);
    nor g7277(n3050 ,n2994 ,n3036);
    not g7278(n5123 ,n5122);
    xnor g7279(n6866 ,n6707 ,n6587);
    or g7280(n1014 ,n684 ,n706);
    nor g7281(n3805 ,n3771 ,n3804);
    not g7282(n5421 ,n5420);
    nor g7283(n3060 ,n3012 ,n3030);
    nor g7284(n1879 ,n107 ,n108);
    xnor g7285(n353 ,n181 ,n185);
    nor g7286(n2495 ,n2472 ,n2465);
    nor g7287(n2606 ,n2442 ,n2574);
    nor g7288(n5600 ,n5204 ,n5120);
    nor g7289(n5676 ,n5491 ,n5421);
    not g7290(n778 ,n3[2]);
    dff g7291(.RN(n1), .SN(1'b1), .CK(n0), .D(n1759), .Q(n28[14]));
    xnor g7292(n7820 ,n3792 ,n3817);
    nor g7293(n3581 ,n3528 ,n3580);
    xnor g7294(n3963 ,n7788 ,n7773);
    nor g7295(n5629 ,n5368 ,n5220);
    nor g7296(n7545 ,n7449 ,n7476);
    not g7297(n3616 ,n7814);
    nor g7298(n5720 ,n5257 ,n5433);
    not g7299(n4681 ,n4680);
    not g7300(n6089 ,n6088);
    nor g7301(n1324 ,n895 ,n642);
    not g7302(n250 ,n249);
    nor g7303(n3693 ,n3664 ,n3649);
    buf g7304(n13[5], n11[5]);
    nor g7305(n5689 ,n5123 ,n5141);
    nor g7306(n5718 ,n5461 ,n5179);
    nor g7307(n1405 ,n668 ,n638);
    dff g7308(.RN(n1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n28[15]));
    nor g7309(n1257 ,n957 ,n637);
    xor g7310(n6189 ,n5776 ,n5348);
    xnor g7311(n6930 ,n6783 ,n6739);
    not g7312(n7413 ,n7721);
    dff g7313(.RN(n1), .SN(1'b1), .CK(n0), .D(n1655), .Q(n35[9]));
    xnor g7314(n6282 ,n6034 ,n6030);
    not g7315(n5431 ,n5430);
    nor g7316(n7508 ,n7436 ,n7475);
    not g7317(n5215 ,n5214);
    nor g7318(n5636 ,n5234 ,n5466);
    nor g7319(n6020 ,n5697 ,n5925);
    nor g7320(n4911 ,n4866 ,n4868);
    nor g7321(n2038 ,n1891 ,n2004);
    or g7322(n1658 ,n1211 ,n1143);
    not g7323(n5473 ,n5472);
    not g7324(n5147 ,n5146);
    nor g7325(n5938 ,n5680 ,n5921);
    nor g7326(n6752 ,n6650 ,n6648);
    nor g7327(n5671 ,n5213 ,n5219);
    nor g7328(n1185 ,n1013 ,n1104);
    nor g7329(n3418 ,n3302 ,n3370);
    nor g7330(n5025 ,n4993 ,n5008);
    nor g7331(n5743 ,n5325 ,n5319);
    xnor g7332(n6928 ,n6777 ,n6821);
    nor g7333(n5180 ,n5095 ,n5099);
    not g7334(n7414 ,n40[9]);
    nor g7335(n5039 ,n5001 ,n5028);
    nor g7336(n5980 ,n5725 ,n5867);
    xnor g7337(n4628 ,n4377 ,n4512);
    nor g7338(n5120 ,n5102 ,n5091);
    nor g7339(n6343 ,n6255 ,n6251);
    nor g7340(n4746 ,n4591 ,n4682);
    nor g7341(n205 ,n147 ,n148);
    not g7342(n252 ,n251);
    nor g7343(n2621 ,n2534 ,n2587);
    xnor g7344(n6124 ,n5763 ,n5470);
    nor g7345(n2231 ,n2078 ,n2191);
    nor g7346(n7211 ,n7175 ,n7160);
    xor g7347(n4560 ,n4390 ,n4172);
    nor g7348(n69 ,n52 ,n68);
    not g7349(n2440 ,n21[0]);
    nor g7350(n2013 ,n1891 ,n1974);
    xnor g7351(n4604 ,n4464 ,n4456);
    nor g7352(n6775 ,n6560 ,n6661);
    nor g7353(n5999 ,n5693 ,n5873);
    nor g7354(n3274 ,n3199 ,n3223);
    not g7355(n691 ,n12[12]);
    nor g7356(n1274 ,n694 ,n638);
    not g7357(n5107 ,n37[4]);
    nor g7358(n1540 ,n768 ,n641);
    nor g7359(n5068 ,n5043 ,n5053);
    dff g7360(.RN(n1), .SN(1'b1), .CK(n0), .D(n1647), .Q(n10[5]));
    or g7361(n7486 ,n7464 ,n7480);
    nor g7362(n1390 ,n674 ,n1103);
    nor g7363(n4948 ,n4853 ,n4905);
    nor g7364(n1453 ,n670 ,n634);
    nor g7365(n4330 ,n4169 ,n4235);
    nor g7366(n3101 ,n3012 ,n3029);
    nor g7367(n4615 ,n4475 ,n4581);
    nor g7368(n4794 ,n4632 ,n4758);
    nor g7369(n1548 ,n697 ,n641);
    not g7370(n5349 ,n5348);
    nor g7371(n4912 ,n4851 ,n4874);
    nor g7372(n5590 ,n5386 ,n5406);
    not g7373(n6653 ,n6652);
    xnor g7374(n4667 ,n4585 ,n4589);
    xnor g7375(n3340 ,n3116 ,n3218);
    nor g7376(n5705 ,n5187 ,n5391);
    nor g7377(n1197 ,n1014 ,n1104);
    xor g7378(n2426 ,n2510 ,n2635);
    nor g7379(n7496 ,n7393 ,n7481);
    not g7380(n6121 ,n6120);
    nor g7381(n1871 ,n134 ,n135);
    not g7382(n780 ,n5[6]);
    or g7383(n1739 ,n1377 ,n1184);
    xnor g7384(n5049 ,n5021 ,n4986);
    nor g7385(n1283 ,n976 ,n637);
    nor g7386(n598 ,n572 ,n588);
    dff g7387(.RN(n1), .SN(1'b1), .CK(n0), .D(n1686), .Q(n24[13]));
    nor g7388(n2957 ,n2862 ,n2925);
    or g7389(n36[0] ,n7687 ,n7685);
    xnor g7390(n7835 ,n3964 ,n3968);
    not g7391(n6530 ,n6529);
    xnor g7392(n6718 ,n6495 ,n6539);
    not g7393(n2788 ,n2428);
    not g7394(n6264 ,n6263);
    nor g7395(n5583 ,n5197 ,n5497);
    xnor g7396(n6596 ,n6241 ,n6488);
    xor g7397(n334 ,n271 ,n187);
    nor g7398(n2528 ,n2443 ,n2521);
    nor g7399(n5710 ,n5125 ,n5475);
    xnor g7400(n6513 ,n6279 ,n5972);
    nor g7401(n7471 ,n7328 ,n7337);
    nor g7402(n461 ,n305 ,n399);
    nor g7403(n7127 ,n7061 ,n7101);
    xnor g7404(n5070 ,n5050 ,n5035);
    nor g7405(n2756 ,n2704 ,n2689);
    or g7406(n4254 ,n4019 ,n4010);
    not g7407(n6643 ,n6642);
    xnor g7408(n2520 ,n2423 ,n2493);
    xnor g7409(n1039 ,n890 ,n664);
    xnor g7410(n5843 ,n5515 ,n5573);
    nor g7411(n6374 ,n6115 ,n6113);
    nor g7412(n6317 ,n6128 ,n6126);
    nor g7413(n4762 ,n4661 ,n4702);
    not g7414(n680 ,n36[10]);
    xnor g7415(n2343 ,n2290 ,n2270);
    or g7416(n1623 ,n1289 ,n1491);
    nor g7417(n2759 ,n2709 ,n2703);
    nor g7418(n5336 ,n5107 ,n5090);
    nor g7419(n4569 ,n4412 ,n4477);
    nor g7420(n3497 ,n3449 ,n3478);
    or g7421(n1005 ,n819 ,n821);
    nor g7422(n2984 ,n2983 ,n2968);
    xnor g7423(n4834 ,n4714 ,n4764);
    not g7424(n789 ,n6[6]);
    nor g7425(n5577 ,n5095 ,n5113);
    nor g7426(n7116 ,n7095 ,n7087);
    not g7427(n7383 ,n7778);
    not g7428(n5355 ,n5354);
    nor g7429(n187 ,n147 ,n158);
    not g7430(n3430 ,n3429);
    not g7431(n3752 ,n3751);
    nor g7432(n4224 ,n4022 ,n4025);
    nor g7433(n3990 ,n3947 ,n3989);
    nor g7434(n3808 ,n3776 ,n3807);
    nor g7435(n2639 ,n2538 ,n2617);
    nor g7436(n3263 ,n3058 ,n3173);
    not g7437(n4025 ,n20[1]);
    xnor g7438(n2084 ,n1959 ,n2007);
    nor g7439(n6967 ,n6756 ,n6889);
    nor g7440(n5625 ,n5412 ,n5154);
    not g7441(n5411 ,n5410);
    xnor g7442(n4548 ,n4397 ,n4232);
    or g7443(n7694 ,n7630 ,n7621);
    xnor g7444(n2318 ,n2247 ,n2272);
    not g7445(n969 ,n25[2]);
    nor g7446(n1301 ,n939 ,n636);
    not g7447(n7037 ,n7036);
    xnor g7448(n5809 ,n5268 ,n5246);
    not g7449(n1839 ,n1840);
    nor g7450(n6889 ,n6762 ,n6840);
    not g7451(n4079 ,n4078);
    dff g7452(.RN(n1), .SN(1'b1), .CK(n0), .D(n1627), .Q(n11[7]));
    nor g7453(n4452 ,n4117 ,n4308);
    nor g7454(n4846 ,n4728 ,n4789);
    or g7455(n7700 ,n7652 ,n7649);
    xnor g7456(n1691 ,n635 ,n33[0]);
    xnor g7457(n4781 ,n4669 ,n4524);
    nor g7458(n2561 ,n2441 ,n2525);
    nor g7459(n6306 ,n6150 ,n6082);
    nor g7460(n306 ,n248 ,n188);
    nor g7461(n2848 ,n2767 ,n2809);
    nor g7462(n2313 ,n2186 ,n2284);
    not g7463(n5267 ,n5266);
    nor g7464(n3210 ,n3090 ,n3185);
    nor g7465(n1458 ,n804 ,n634);
    not g7466(n4989 ,n4988);
    not g7467(n3020 ,n40[6]);
    nor g7468(n1343 ,n725 ,n636);
    xnor g7469(n347 ,n269 ,n259);
    xnor g7470(n4554 ,n4379 ,n4114);
    or g7471(n1748 ,n1388 ,n1153);
    nor g7472(n4230 ,n4006 ,n4017);
    not g7473(n2300 ,n2299);
    or g7474(n5759 ,n5353 ,n5316);
    or g7475(n5547 ,n5099 ,n5098);
    nor g7476(n7573 ,n7431 ,n7474);
    nor g7477(n128 ,n33[1] ,n33[0]);
    nor g7478(n7250 ,n7220 ,n7178);
    xnor g7479(n3672 ,n7803 ,n7780);
    xnor g7480(n2906 ,n2860 ,n2845);
    xnor g7481(n6263 ,n5781 ,n5557);
    not g7482(n4016 ,n20[7]);
    nor g7483(n3446 ,n3398 ,n3400);
    not g7484(n3203 ,n3202);
    not g7485(n3824 ,n19[2]);
    or g7486(n1720 ,n1360 ,n1180);
    nor g7487(n5608 ,n5176 ,n5244);
    nor g7488(n4621 ,n4482 ,n4580);
    nor g7489(n626 ,n613 ,n625);
    nor g7490(n322 ,n264 ,n274);
    xnor g7491(n6426 ,n6068 ,n6059);
    nor g7492(n7490 ,n7403 ,n7480);
    or g7493(n984 ,n35[4] ,n35[11]);
    xnor g7494(n6598 ,n6486 ,n6475);
    xnor g7495(n6721 ,n6497 ,n6571);
    nor g7496(n7549 ,n7450 ,n7475);
    nor g7497(n6732 ,n6581 ,n6674);
    xnor g7498(n7079 ,n6981 ,n6940);
    nor g7499(n4960 ,n4891 ,n4948);
    xnor g7500(n6527 ,n6290 ,n6044);
    or g7501(n5533 ,n5102 ,n5090);
    nor g7502(n1555 ,n907 ,n1100);
    nor g7503(n3640 ,n39[9] ,n7810);
    not g7504(n4461 ,n4460);
    not g7505(n5143 ,n5142);
    xnor g7506(n3065 ,n40[3] ,n7742);
    xnor g7507(n396 ,n346 ,n231);
    nor g7508(n4618 ,n4554 ,n4552);
    not g7509(n6143 ,n6142);
    nor g7510(n4712 ,n4571 ,n4617);
    nor g7511(n458 ,n385 ,n424);
    xnor g7512(n2776 ,n2659 ,n2729);
    nor g7513(n5662 ,n5485 ,n5183);
    not g7514(n2748 ,n2747);
    nor g7515(n2404 ,n2378 ,n2393);
    not g7516(n5505 ,n5504);
    nor g7517(n7231 ,n7157 ,n7203);
    not g7518(n4352 ,n4351);
    or g7519(n7648 ,n7562 ,n7561);
    nor g7520(n1532 ,n775 ,n641);
    not g7521(n3617 ,n7788);
    not g7522(n3704 ,n3703);
    buf g7523(n13[12], n10[12]);
    or g7524(n2003 ,n1966 ,n1973);
    xnor g7525(n2172 ,n1970 ,n2085);
    nor g7526(n5246 ,n5096 ,n5102);
    xnor g7527(n6116 ,n5789 ,n5120);
    not g7528(n874 ,n21[2]);
    xnor g7529(n4605 ,n4458 ,n4476);
    nor g7530(n7599 ,n7398 ,n7475);
    or g7531(n7626 ,n7523 ,n7522);
    xnor g7532(n3733 ,n39[2] ,n3672);
    nor g7533(n1360 ,n867 ,n1107);
    not g7534(n737 ,n6[0]);
    xnor g7535(n2671 ,n2501 ,n2584);
    xnor g7536(n2702 ,n2644 ,n2513);
    nor g7537(n1403 ,n900 ,n642);
    nor g7538(n5394 ,n5095 ,n5092);
    not g7539(n6129 ,n6128);
    or g7540(n2002 ,n1965 ,n1979);
    not g7541(n3003 ,n40[13]);
    xnor g7542(n2247 ,n2079 ,n2207);
    not g7543(n4537 ,n4536);
    nor g7544(n6340 ,n5996 ,n6217);
    nor g7545(n3106 ,n3013 ,n3039);
    not g7546(n910 ,n19[4]);
    nor g7547(n4267 ,n4018 ,n4010);
    nor g7548(n4034 ,n4011 ,n4019);
    xnor g7549(n526 ,n476 ,n384);
    nor g7550(n1516 ,n769 ,n1099);
    nor g7551(n2897 ,n2817 ,n2876);
    nor g7552(n225 ,n154 ,n149);
    not g7553(n2029 ,n2028);
    nor g7554(n7530 ,n7409 ,n7480);
    nor g7555(n1142 ,n641 ,n1084);
    not g7556(n3153 ,n3152);
    nor g7557(n4334 ,n4211 ,n4183);
    nor g7558(n2749 ,n2633 ,n2725);
    xnor g7559(n3332 ,n3148 ,n3206);
    nor g7560(n6697 ,n6131 ,n6536);
    nor g7561(n319 ,n224 ,n226);
    or g7562(n7678 ,n7589 ,n7670);
    xnor g7563(n2708 ,n2515 ,n2648);
    nor g7564(n7009 ,n6857 ,n6932);
    nor g7565(n4745 ,n4592 ,n4683);
    not g7566(n3258 ,n3257);
    or g7567(n1634 ,n1301 ,n1234);
    not g7568(n914 ,n24[10]);
    not g7569(n2840 ,n2839);
    nor g7570(n4178 ,n4023 ,n4008);
    not g7571(n674 ,n23[1]);
    nor g7572(n4162 ,n4020 ,n4024);
    not g7573(n5499 ,n5498);
    nor g7574(n5488 ,n5092 ,n5090);
    not g7575(n5527 ,n5526);
    xor g7576(n40[12] ,n39[13] ,n7827);
    not g7577(n7368 ,n39[9]);
    not g7578(n2124 ,n2123);
    not g7579(n5189 ,n5188);
    not g7580(n48 ,n19[5]);
    xnor g7581(n4787 ,n4671 ,n4563);
    nor g7582(n6898 ,n6642 ,n6824);
    xnor g7583(n2268 ,n2218 ,n2136);
    nor g7584(n1323 ,n696 ,n1101);
    xnor g7585(n6168 ,n5812 ,n5526);
    nor g7586(n4451 ,n4097 ,n4358);
    xnor g7587(n3465 ,n3361 ,n3418);
    nor g7588(n4731 ,n4658 ,n4698);
    or g7589(n1609 ,n1273 ,n1119);
    nor g7590(n6677 ,n6474 ,n6521);
    nor g7591(n6554 ,n6249 ,n6436);
    xnor g7592(n1965 ,n1954 ,n1925);
    nor g7593(n2825 ,n2743 ,n2792);
    or g7594(n1669 ,n1328 ,n1522);
    xnor g7595(n3890 ,n7798 ,n7810);
    not g7596(n402 ,n401);
    not g7597(n4952 ,n4951);
    nor g7598(n3714 ,n3657 ,n3687);
    not g7599(n6623 ,n6622);
    nor g7600(n2653 ,n2565 ,n2608);
    nor g7601(n4068 ,n4008 ,n4025);
    not g7602(n2751 ,n2430);
    or g7603(n7686 ,n7624 ,n7622);
    nor g7604(n7778 ,n4279 ,n4348);
    nor g7605(n3477 ,n3415 ,n3434);
    nor g7606(n7572 ,n7447 ,n7479);
    nor g7607(n5893 ,n5289 ,n5631);
    not g7608(n4213 ,n4212);
    not g7609(n1908 ,n19[2]);
    or g7610(n1671 ,n1330 ,n1541);
    not g7611(n3016 ,n40[2]);
    not g7612(n42 ,n19[2]);
    nor g7613(n4052 ,n4019 ,n4025);
    nor g7614(n2642 ,n2542 ,n2618);
    xnor g7615(n6335 ,n5809 ,n6060);
    nor g7616(n6750 ,n6652 ,n6646);
    dff g7617(.RN(n1), .SN(1'b1), .CK(n0), .D(n1648), .Q(n35[14]));
    not g7618(n2842 ,n2841);
    not g7619(n947 ,n12[8]);
    nor g7620(n4343 ,n4165 ,n4065);
    nor g7621(n3230 ,n3059 ,n3170);
    not g7622(n2441 ,n7764);
    nor g7623(n1292 ,n929 ,n636);
    not g7624(n153 ,n19[1]);
    xnor g7625(n7828 ,n3963 ,n3984);
    not g7626(n188 ,n187);
    or g7627(n7683 ,n7614 ,n7612);
    nor g7628(n3168 ,n2995 ,n3072);
    nor g7629(n4852 ,n4705 ,n4812);
    nor g7630(n4110 ,n4013 ,n4020);
    not g7631(n5541 ,n5540);
    or g7632(n997 ,n808 ,n18[1]);
    nor g7633(n1443 ,n841 ,n634);
    not g7634(n822 ,n24[5]);
    not g7635(n845 ,n22[2]);
    nor g7636(n5890 ,n5310 ,n5651);
    xnor g7637(n2932 ,n2885 ,n2855);
    not g7638(n2921 ,n2920);
    nor g7639(n2198 ,n2145 ,n2150);
    nor g7640(n1330 ,n940 ,n642);
    xnor g7641(n1034 ,n871 ,n845);
    nor g7642(n5592 ,n5394 ,n5230);
    nor g7643(n2983 ,n2950 ,n2982);
    nor g7644(n1388 ,n897 ,n1101);
    nor g7645(n5618 ,n5446 ,n5436);
    nor g7646(n4992 ,n4949 ,n4959);
    nor g7647(n5170 ,n5102 ,n5116);
    nor g7648(n7525 ,n7330 ,n7481);
    xnor g7649(n3331 ,n3154 ,n3259);
    xnor g7650(n1046 ,n690 ,n822);
    not g7651(n664 ,n22[7]);
    nor g7652(n5511 ,n5103 ,n5110);
    nor g7653(n3461 ,n3387 ,n3429);
    not g7654(n6496 ,n6495);
    nor g7655(n3965 ,n3950 ,n3955);
    nor g7656(n6812 ,n6592 ,n6752);
    nor g7657(n1094 ,n986 ,n994);
    nor g7658(n3654 ,n3626 ,n3595);
    nor g7659(n7526 ,n7404 ,n7474);
    nor g7660(n570 ,n519 ,n558);
    not g7661(n3023 ,n40[10]);
    nor g7662(n6770 ,n6506 ,n6623);
    nor g7663(n493 ,n192 ,n453);
    xnor g7664(n64 ,n37[4] ,n19[4]);
    xnor g7665(n6940 ,n6779 ,n6840);
    not g7666(n5516 ,n5515);
    not g7667(n921 ,n11[11]);
    xnor g7668(n4793 ,n4668 ,n4688);
    nor g7669(n2800 ,n2727 ,n2758);
    nor g7670(n4050 ,n4027 ,n4019);
    nor g7671(n4301 ,n4056 ,n4152);
    nor g7672(n4775 ,n4713 ,n4749);
    dff g7673(.RN(n1), .SN(1'b1), .CK(n0), .D(n1656), .Q(n10[3]));
    xnor g7674(n7832 ,n3953 ,n3976);
    not g7675(n4738 ,n4737);
    not g7676(n3629 ,n39[7]);
    not g7677(n4223 ,n4222);
    xnor g7678(n2902 ,n2868 ,n2786);
    not g7679(n875 ,n31[5]);
    nor g7680(n5640 ,n5158 ,n5242);
    nor g7681(n4074 ,n4011 ,n4020);
    nor g7682(n4754 ,n4656 ,n4696);
    or g7683(n1578 ,n1239 ,n1517);
    or g7684(n5312 ,n5091 ,n5105);
    nor g7685(n7521 ,n7424 ,n7481);
    not g7686(n2142 ,n2141);
    nor g7687(n6198 ,n5954 ,n5946);
    xnor g7688(n4729 ,n4608 ,n4475);
    xnor g7689(n7118 ,n7025 ,n7000);
    xor g7690(n7834 ,n3961 ,n3971);
    or g7691(n1583 ,n1244 ,n1111);
    not g7692(n5195 ,n5194);
    not g7693(n683 ,n36[13]);
    nor g7694(n5968 ,n5730 ,n5883);
    not g7695(n3713 ,n3712);
    nor g7696(n3722 ,n3660 ,n3689);
    nor g7697(n2305 ,n2263 ,n2285);
    not g7698(n170 ,n169);
    not g7699(n4051 ,n4050);
    not g7700(n6931 ,n6930);
    nor g7701(n5861 ,n5334 ,n5617);
    xnor g7702(n6074 ,n5829 ,n5170);
    not g7703(n7384 ,n7735);
    nor g7704(n3873 ,n7802 ,n7794);
    buf g7705(n428 ,n328);
    nor g7706(n5613 ,n5278 ,n5164);
    nor g7707(n3857 ,n3846 ,n3856);
    not g7708(n899 ,n10[4]);
    nor g7709(n1866 ,n57 ,n55);
    xnor g7710(n2168 ,n1968 ,n2097);
    nor g7711(n181 ,n156 ,n157);
    nor g7712(n6950 ,n6908 ,n6866);
    not g7713(n4405 ,n4404);
    not g7714(n971 ,n33[3]);
    nor g7715(n2962 ,n2916 ,n2957);
    nor g7716(n6207 ,n6005 ,n6017);
    nor g7717(n3278 ,n3118 ,n3205);
    xnor g7718(n3956 ,n7790 ,n7775);
    xnor g7719(n7815 ,n2381 ,n2420);
    xnor g7720(n7756 ,n4001 ,n3998);
    not g7721(n2242 ,n2241);
    xnor g7722(n5776 ,n5480 ,n5150);
    nor g7723(n2573 ,n2431 ,n2525);
    xnor g7724(n5846 ,n5513 ,n5522);
    nor g7725(n2731 ,n2551 ,n2670);
    not g7726(n242 ,n241);
    nor g7727(n6054 ,n5721 ,n5871);
    nor g7728(n4997 ,n4924 ,n4984);
    nor g7729(n7462 ,n41[14] ,n7818);
    xnor g7730(n2151 ,n1972 ,n2070);
    not g7731(n3139 ,n3138);
    not g7732(n852 ,n20[0]);
    xnor g7733(n4612 ,n4176 ,n4470);
    dff g7734(.RN(n1), .SN(1'b1), .CK(n0), .D(n1676), .Q(n25[1]));
    xnor g7735(n1073 ,n24[4] ,n35[4]);
    dff g7736(.RN(n1), .SN(1'b1), .CK(n0), .D(n1711), .Q(n34[11]));
    not g7737(n4525 ,n4524);
    nor g7738(n6469 ,n6216 ,n6326);
    not g7739(n6276 ,n6275);
    nor g7740(n7059 ,n7021 ,n7011);
    nor g7741(n500 ,n435 ,n481);
    or g7742(n1624 ,n1288 ,n1447);
    xnor g7743(n2472 ,n2446 ,n21[4]);
    nor g7744(n5168 ,n5116 ,n5094);
    nor g7745(n283 ,n169 ,n239);
    xnor g7746(n3784 ,n3745 ,n3697);
    not g7747(n3394 ,n3393);
    nor g7748(n5200 ,n5107 ,n5100);
    not g7749(n1922 ,n1921);
    xnor g7750(n3725 ,n39[13] ,n3669);
    nor g7751(n3860 ,n3842 ,n3859);
    nor g7752(n134 ,n33[3] ,n132);
    nor g7753(n4004 ,n4000 ,n4003);
    xor g7754(n40[8] ,n39[9] ,n7831);
    nor g7755(n6442 ,n6218 ,n6340);
    not g7756(n956 ,n10[14]);
    nor g7757(n5704 ,n5423 ,n5489);
    nor g7758(n1444 ,n667 ,n634);
    or g7759(n1761 ,n1401 ,n1496);
    nor g7760(n7311 ,n7310 ,n7282);
    not g7761(n3123 ,n3122);
    xnor g7762(n4715 ,n4530 ,n4636);
    not g7763(n4015 ,n19[1]);
    xnor g7764(n1087 ,n864 ,n827);
    nor g7765(n4297 ,n4050 ,n4188);
    not g7766(n804 ,n1868);
    not g7767(n4356 ,n4355);
    not g7768(n5316 ,n5315);
    nor g7769(n4908 ,n4843 ,n4862);
    nor g7770(n6302 ,n5998 ,n6223);
    xnor g7771(n4723 ,n4605 ,n4558);
    xnor g7772(n609 ,n582 ,n577);
    nor g7773(n6466 ,n6276 ,n6343);
    not g7774(n960 ,n29[5]);
    not g7775(n5211 ,n5210);
    nor g7776(n5008 ,n4952 ,n4981);
    or g7777(n1754 ,n1392 ,n1156);
    not g7778(n7426 ,n7716);
    not g7779(n6164 ,n6163);
    nor g7780(n1344 ,n681 ,n640);
    xnor g7781(n3535 ,n3481 ,n3438);
    nor g7782(n1251 ,n925 ,n636);
    nor g7783(n5384 ,n5119 ,n5103);
    nor g7784(n4273 ,n4030 ,n4074);
    xnor g7785(n7258 ,n7217 ,n7222);
    not g7786(n3119 ,n3118);
    nor g7787(n3277 ,n3198 ,n3266);
    xnor g7788(n6974 ,n6620 ,n6884);
    nor g7789(n2503 ,n2481 ,n2492);
    nor g7790(n6558 ,n6470 ,n6422);
    nor g7791(n5906 ,n5532 ,n5591);
    nor g7792(n7472 ,n7332 ,n7397);
    nor g7793(n427 ,n324 ,n377);
    xnor g7794(n4565 ,n4402 ,n4216);
    nor g7795(n6357 ,n6159 ,n6233);
    or g7796(n7624 ,n7521 ,n7520);
    not g7797(n3736 ,n3735);
    nor g7798(n7208 ,n7099 ,n7166);
    nor g7799(n1464 ,n851 ,n634);
    nor g7800(n6208 ,n5940 ,n5944);
    nor g7801(n2474 ,n2446 ,n2456);
    nor g7802(n6345 ,n6267 ,n6263);
    not g7803(n7390 ,n7723);
    nor g7804(n7570 ,n7406 ,n7481);
    not g7805(n667 ,n34[12]);
    nor g7806(n6388 ,n6101 ,n6079);
    nor g7807(n3687 ,n3628 ,n3646);
    not g7808(n3767 ,n3766);
    xnor g7809(n7816 ,n2339 ,n2422);
    or g7810(n4145 ,n4006 ,n4026);
    nor g7811(n2228 ,n2084 ,n2192);
    nor g7812(n1130 ,n635 ,n1035);
    nor g7813(n3574 ,n3543 ,n3573);
    nor g7814(n1303 ,n707 ,n636);
    nor g7815(n4284 ,n4046 ,n4194);
    nor g7816(n3760 ,n3718 ,n3748);
    or g7817(n5538 ,n5102 ,n5098);
    xnor g7818(n6436 ,n6070 ,n5749);
    not g7819(n3402 ,n3401);
    not g7820(n5435 ,n5434);
    nor g7821(n3709 ,n3652 ,n3691);
    or g7822(n5518 ,n5107 ,n5097);
    nor g7823(n7026 ,n7020 ,n6950);
    nor g7824(n3253 ,n3046 ,n3126);
    xnor g7825(n4375 ,n4086 ,n4212);
    not g7826(n7299 ,n7298);
    nor g7827(n7456 ,n41[13] ,n7819);
    dff g7828(.RN(n1), .SN(1'b1), .CK(n0), .D(n1720), .Q(n31[6]));
    nor g7829(n6681 ,n6569 ,n6530);
    nor g7830(n1267 ,n904 ,n636);
    not g7831(n2665 ,n2664);
    nor g7832(n1319 ,n837 ,n637);
    xnor g7833(n4733 ,n4609 ,n4593);
    nor g7834(n304 ,n210 ,n208);
    nor g7835(n3501 ,n3441 ,n3472);
    nor g7836(n1531 ,n728 ,n641);
    or g7837(n641 ,n18[2] ,n997);
    not g7838(n5531 ,n5530);
    nor g7839(n6320 ,n6004 ,n6236);
    nor g7840(n1017 ,n644 ,n18[0]);
    xnor g7841(n6150 ,n5813 ,n5504);
    not g7842(n2314 ,n2313);
    nor g7843(n6953 ,n6805 ,n6855);
    nor g7844(n1566 ,n676 ,n634);
    not g7845(n5558 ,n5557);
    not g7846(n843 ,n22[6]);
    nor g7847(n555 ,n508 ,n529);
    nor g7848(n3977 ,n3953 ,n3976);
    nor g7849(n1461 ,n800 ,n634);
    nor g7850(n1275 ,n927 ,n636);
    not g7851(n881 ,n31[3]);
    not g7852(n3015 ,n7745);
    nor g7853(n1339 ,n894 ,n642);
    not g7854(n3522 ,n3521);
    nor g7855(n5079 ,n5068 ,n5078);
    xnor g7856(n6067 ,n5835 ,n5747);
    nor g7857(n6012 ,n5756 ,n5839);
    not g7858(n888 ,n28[0]);
    nor g7859(n5313 ,n5095 ,n5114);
    xnor g7860(n6626 ,n6409 ,n6263);
    nor g7861(n4315 ,n4179 ,n4039);
    nor g7862(n7594 ,n7411 ,n7479);
    xor g7863(n7746 ,n7808 ,n7785);
    xnor g7864(n1065 ,n811 ,n838);
    nor g7865(n3126 ,n3012 ,n3073);
    nor g7866(n6577 ,n6358 ,n6457);
    not g7867(n7362 ,n7777);
    nor g7868(n491 ,n408 ,n455);
    buf g7869(n13[1], n10[1]);
    not g7870(n5155 ,n5154);
    dff g7871(.RN(n1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n20[4]));
    nor g7872(n7670 ,n7468 ,n7485);
    not g7873(n603 ,n602);
    not g7874(n5391 ,n5390);
    not g7875(n4547 ,n4546);
    not g7876(n2110 ,n2109);
    nor g7877(n7298 ,n7271 ,n7266);
    nor g7878(n1568 ,n680 ,n634);
    xnor g7879(n4001 ,n37[1] ,n20[1]);
    xnor g7880(n2710 ,n2515 ,n2623);
    xnor g7881(n1968 ,n1949 ,n1928);
    or g7882(n1741 ,n1222 ,n1190);
    or g7883(n7619 ,n7507 ,n7506);
    nor g7884(n6559 ,n6469 ,n6423);
    not g7885(n533 ,n532);
    nor g7886(n4170 ,n4019 ,n4026);
    nor g7887(n4804 ,n4666 ,n4741);
    nor g7888(n6841 ,n6682 ,n6745);
    nor g7889(n5606 ,n5460 ,n5178);
    nor g7890(n1110 ,n635 ,n1020);
    not g7891(n4147 ,n4146);
    not g7892(n916 ,n29[7]);
    xnor g7893(n3743 ,n39[5] ,n3678);
    xnor g7894(n7068 ,n6930 ,n7019);
    nor g7895(n2763 ,n2664 ,n2723);
    nor g7896(n201 ,n154 ,n155);
    or g7897(n4244 ,n4006 ,n4028);
    nor g7898(n2676 ,n2501 ,n2655);
    not g7899(n166 ,n165);
    nor g7900(n2180 ,n2080 ,n2141);
    xnor g7901(n3334 ,n3220 ,n3202);
    nor g7902(n2596 ,n2442 ,n2547);
    nor g7903(n7846 ,n3886 ,n3885);
    nor g7904(n5412 ,n5117 ,n5093);
    nor g7905(n215 ,n145 ,n153);
    xnor g7906(n3381 ,n3320 ,n3222);
    nor g7907(n301 ,n233 ,n171);
    nor g7908(n7235 ,n7187 ,n7197);
    not g7909(n723 ,n10[8]);
    nor g7910(n5234 ,n5099 ,n5100);
    nor g7911(n4307 ,n4172 ,n4186);
    not g7912(n2717 ,n2427);
    or g7913(n1576 ,n1237 ,n1467);
    xnor g7914(n6642 ,n6408 ,n6482);
    xnor g7915(n3505 ,n3452 ,n3429);
    nor g7916(n2874 ,n2810 ,n2834);
    dff g7917(.RN(n1), .SN(1'b1), .CK(n0), .D(n1675), .Q(n34[10]));
    not g7918(n112 ,n111);
    xnor g7919(n3549 ,n3511 ,n3491);
    not g7920(n5748 ,n5747);
    not g7921(n3105 ,n3104);
    xnor g7922(n7783 ,n4972 ,n4990);
    not g7923(n157 ,n19[5]);
    or g7924(n4264 ,n4018 ,n4016);
    nor g7925(n4751 ,n4651 ,n4689);
    nor g7926(n6377 ,n6141 ,n6135);
    nor g7927(n987 ,n643 ,n18[0]);
    xnor g7928(n3785 ,n3743 ,n3714);
    nor g7929(n2490 ,n2460 ,n2475);
    nor g7930(n5912 ,n5309 ,n5614);
    xnor g7931(n1964 ,n1942 ,n1940);
    nor g7932(n2892 ,n2873 ,n2869);
    nor g7933(n4474 ,n4328 ,n4435);
    nor g7934(n1426 ,n885 ,n638);
    or g7935(n7698 ,n7648 ,n7647);
    nor g7936(n2497 ,n2433 ,n2477);
    not g7937(n1100 ,n1101);
    xnor g7938(n6843 ,n6618 ,n6774);
    nor g7939(n4620 ,n4546 ,n4587);
    not g7940(n412 ,n411);
    nor g7941(n3292 ,n3267 ,n3226);
    nor g7942(n449 ,n311 ,n423);
    nor g7943(n5933 ,n5853 ,n5845);
    nor g7944(n1991 ,n1902 ,n1976);
    xnor g7945(n3069 ,n40[10] ,n7749);
    nor g7946(n3689 ,n3634 ,n3639);
    nor g7947(n5242 ,n5098 ,n5113);
    nor g7948(n5392 ,n5093 ,n5109);
    xor g7949(n7791 ,n5048 ,n5083);
    nor g7950(n490 ,n380 ,n446);
    xnor g7951(n4518 ,n4382 ,n4050);
    nor g7952(n3051 ,n2994 ,n3029);
    not g7953(n6494 ,n6493);
    not g7954(n5275 ,n5274);
    nor g7955(n4797 ,n4708 ,n4755);
    not g7956(n5207 ,n5206);
    nor g7957(n4472 ,n4339 ,n4421);
    nor g7958(n6373 ,n6109 ,n6107);
    nor g7959(n5024 ,n4953 ,n5006);
    nor g7960(n3474 ,n3402 ,n3432);
    not g7961(n4916 ,n4915);
    not g7962(n5243 ,n5242);
    nor g7963(n1569 ,n675 ,n634);
    nor g7964(n1918 ,n1897 ,n1907);
    or g7965(n1678 ,n1281 ,n1570);
    not g7966(n330 ,n329);
    xnor g7967(n3482 ,n3359 ,n3440);
    not g7968(n5209 ,n5208);
    nor g7969(n5304 ,n5115 ,n5110);
    not g7970(n2995 ,n7757);
    nor g7971(n3308 ,n3145 ,n3255);
    not g7972(n4718 ,n4717);
    not g7973(n3969 ,n3968);
    nor g7974(n2876 ,n2838 ,n2836);
    not g7975(n6572 ,n6571);
    nor g7976(n6679 ,n6570 ,n6529);
    xnor g7977(n3071 ,n40[11] ,n7750);
    not g7978(n7360 ,n7737);
    nor g7979(n5559 ,n5101 ,n5094);
    xnor g7980(n2778 ,n2698 ,n2697);
    xnor g7981(n395 ,n349 ,n322);
    nor g7982(n1472 ,n742 ,n639);
    not g7983(n4011 ,n19[6]);
    not g7984(n3213 ,n3212);
    xnor g7985(n546 ,n503 ,n449);
    xnor g7986(n3964 ,n38[4] ,n7781);
    xnor g7987(n3485 ,n3427 ,n3383);
    nor g7988(n6848 ,n6628 ,n6831);
    not g7989(n5975 ,n5974);
    nor g7990(n7189 ,n7063 ,n7141);
    nor g7991(n7537 ,n7434 ,n7474);
    nor g7992(n3448 ,n3381 ,n3379);
    not g7993(n3594 ,n7815);
    nor g7994(n1362 ,n875 ,n1107);
    nor g7995(n4164 ,n4023 ,n4006);
    nor g7996(n1245 ,n690 ,n640);
    not g7997(n2888 ,n2887);
    xor g7998(n5786 ,n5545 ,n5192);
    nor g7999(n5644 ,n5190 ,n5354);
    not g8000(n2298 ,n2297);
    xnor g8001(n3567 ,n3533 ,n3521);
    not g8002(n824 ,n35[4]);
    nor g8003(n5154 ,n5093 ,n5094);
    or g8004(n2206 ,n1971 ,n2156);
    nor g8005(n2088 ,n1992 ,n2039);
    not g8006(n829 ,n23[2]);
    nor g8007(n4200 ,n4011 ,n4022);
    xnor g8008(n39[0] ,n2502 ,n2524);
    nor g8009(n3922 ,n3897 ,n3921);
    nor g8010(n1437 ,n830 ,n640);
    nor g8011(n1439 ,n704 ,n638);
    nor g8012(n2939 ,n2899 ,n2908);
    nor g8013(n2473 ,n2436 ,n2455);
    not g8014(n6807 ,n6806);
    nor g8015(n4889 ,n4810 ,n4826);
    not g8016(n7455 ,n39[11]);
    nor g8017(n3440 ,n3279 ,n3403);
    nor g8018(n2068 ,n1987 ,n2041);
    not g8019(n6035 ,n6034);
    or g8020(n1660 ,n1320 ,n1464);
    buf g8021(n37[7] ,n1838);
    not g8022(n949 ,n10[9]);
    xnor g8023(n5760 ,n5412 ,n5154);
    nor g8024(n3098 ,n2994 ,n3042);
    nor g8025(n2249 ,n2194 ,n2237);
    not g8026(n7072 ,n7071);
    nor g8027(n3800 ,n3758 ,n3799);
    xnor g8028(n6281 ,n6026 ,n6064);
    dff g8029(.RN(n1), .SN(1'b1), .CK(n0), .D(n1614), .Q(n11[15]));
    not g8030(n5599 ,n5260);
    nor g8031(n5864 ,n5305 ,n5613);
    nor g8032(n5372 ,n5088 ,n5109);
    nor g8033(n6316 ,n6102 ,n6257);
    not g8034(n6270 ,n6269);
    nor g8035(n3181 ,n2995 ,n3069);
    nor g8036(n129 ,n125 ,n122);
    dff g8037(.RN(n1), .SN(1'b1), .CK(n0), .D(n1801), .Q(n20[5]));
    nor g8038(n1318 ,n899 ,n636);
    nor g8039(n1984 ,n1892 ,n1980);
    or g8040(n7650 ,n7565 ,n7564);
    xnor g8041(n1079 ,n809 ,n820);
    nor g8042(n4431 ,n4081 ,n4354);
    nor g8043(n5884 ,n5534 ,n5634);
    nor g8044(n6815 ,n6591 ,n6767);
    not g8045(n7429 ,n39[14]);
    not g8046(n452 ,n451);
    dff g8047(.RN(n1), .SN(1'b1), .CK(n0), .D(n1721), .Q(n24[0]));
    xnor g8048(n6069 ,n5842 ,n5270);
    nor g8049(n519 ,n468 ,n494);
    nor g8050(n7582 ,n7413 ,n7480);
    xnor g8051(n4522 ,n4368 ,n4060);
    not g8052(n2140 ,n2139);
    nor g8053(n1433 ,n908 ,n1101);
    nor g8054(n7006 ,n6909 ,n6964);
    not g8055(n697 ,n24[9]);
    nor g8056(n7761 ,n3839 ,n3837);
    nor g8057(n1561 ,n966 ,n1106);
    not g8058(n857 ,n16[6]);
    not g8059(n652 ,n17[2]);
    nor g8060(n7115 ,n7077 ,n7075);
    nor g8061(n2875 ,n2745 ,n2857);
    nor g8062(n279 ,n156 ,n151);
    xnor g8063(n4719 ,n4613 ,n4536);
    xnor g8064(n4822 ,n4741 ,n4665);
    or g8065(n1744 ,n1382 ,n1148);
    not g8066(n5225 ,n5224);
    nor g8067(n4445 ,n4255 ,n4307);
    xor g8068(n2290 ,n2221 ,n2250);
    nor g8069(n5290 ,n5088 ,n5113);
    nor g8070(n2605 ,n2432 ,n2547);
    nor g8071(n6804 ,n6608 ,n6725);
    nor g8072(n6227 ,n5987 ,n5979);
    nor g8073(n5603 ,n5456 ,n5416);
    nor g8074(n6221 ,n5955 ,n5947);
    nor g8075(n381 ,n306 ,n359);
    xnor g8076(n2239 ,n1972 ,n2156);
    xor g8077(n7730 ,n3551 ,n3573);
    not g8078(n4144 ,n4143);
    not g8079(n5141 ,n5140);
    not g8080(n2512 ,n2513);
    buf g8081(n14[0], n11[0]);
    nor g8082(n4003 ,n3997 ,n4002);
    nor g8083(n3136 ,n3012 ,n3065);
    not g8084(n4049 ,n4048);
    nor g8085(n4082 ,n4015 ,n4018);
    nor g8086(n2158 ,n2104 ,n2122);
    nor g8087(n549 ,n437 ,n534);
    xnor g8088(n3553 ,n3513 ,n3479);
    xnor g8089(n7720 ,n3789 ,n3811);
    not g8090(n976 ,n11[12]);
    nor g8091(n6382 ,n6091 ,n6260);
    not g8092(n821 ,n35[6]);
    or g8093(n2549 ,n2506 ,n2520);
    nor g8094(n6829 ,n6675 ,n6729);
    nor g8095(n3905 ,n3875 ,n3904);
    not g8096(n5333 ,n5332);
    xnor g8097(n3766 ,n7779 ,n3694);
    nor g8098(n2181 ,n2162 ,n2143);
    dff g8099(.RN(n1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n21[6]));
    or g8100(n1719 ,n1358 ,n1565);
    nor g8101(n5084 ,n5047 ,n5083);
    not g8102(n6879 ,n6878);
    not g8103(n2435 ,n21[1]);
    or g8104(n7487 ,n7461 ,n7480);
    dff g8105(.RN(n1), .SN(1'b1), .CK(n0), .D(n1573), .Q(n34[0]));
    nor g8106(n3587 ,n3529 ,n3586);
    not g8107(n3221 ,n3220);
    not g8108(n3151 ,n3150);
    not g8109(n717 ,n1831);
    xnor g8110(n6786 ,n6594 ,n6567);
    not g8111(n7428 ,n39[8]);
    not g8112(n2678 ,n2677);
    nor g8113(n5698 ,n5409 ,n5283);
    nor g8114(n7574 ,n7422 ,n7476);
    not g8115(n5953 ,n5952);
    nor g8116(n3859 ,n3847 ,n3858);
    not g8117(n919 ,n10[6]);
    nor g8118(n7587 ,n7359 ,n7477);
    nor g8119(n229 ,n145 ,n148);
    not g8120(n6627 ,n6626);
    or g8121(n1746 ,n1386 ,n1152);
    xor g8122(n7739 ,n7778 ,n7801);
    not g8123(n4897 ,n4896);
    or g8124(n1640 ,n1308 ,n1567);
    not g8125(n922 ,n24[11]);
    xnor g8126(n4536 ,n4380 ,n4116);
    dff g8127(.RN(n1), .SN(1'b1), .CK(n0), .D(n1728), .Q(n31[1]));
    dff g8128(.RN(n1), .SN(1'b1), .CK(n0), .D(n1589), .Q(n12[10]));
    not g8129(n5279 ,n5278);
    nor g8130(n4168 ,n4029 ,n4007);
    nor g8131(n1304 ,n950 ,n636);
    xnor g8132(n579 ,n552 ,n540);
    or g8133(n996 ,n35[2] ,n35[3]);
    xnor g8134(n7797 ,n7287 ,n7300);
    not g8135(n6546 ,n6545);
    not g8136(n842 ,n17[0]);
    nor g8137(n7093 ,n7019 ,n7057);
    not g8138(n944 ,n25[4]);
    nor g8139(n7113 ,n7038 ,n7071);
    nor g8140(n6960 ,n6803 ,n6852);
    nor g8141(n3130 ,n3012 ,n3071);
    nor g8142(n1326 ,n851 ,n637);
    nor g8143(n5458 ,n5103 ,n5113);
    nor g8144(n2008 ,n1892 ,n1976);
endmodule
