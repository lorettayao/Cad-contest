module top(n0, n1, n2, n3, n4, n7, n8, n5, n6, n9, n11, n12, n13, n10);
    input n0, n1, n2, n3, n4, n5, n6;
    input [1:0] n7;
    input [7:0] n8;
    output [7:0] n9, n10;
    output n11, n12, n13;
    wire n0, n1, n2, n3, n4, n5, n6;
    wire [1:0] n7;
    wire [7:0] n8;
    wire [7:0] n9, n10;
    wire n11, n12, n13;
    wire n14, n15, n16, n17, n18, n19, n20, n21;
    wire n22, n23, n24, n25, n26, n27, n28, n29;
    wire n30, n31, n32, n33, n34, n35, n36, n37;
    wire n38, n39, n40, n41, n42, n43, n44, n45;
    wire n46, n47, n48, n49, n50, n51, n52, n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171;
    buf g0(n10[0], n9[0]);
    buf g1(n10[1], n9[1]);
    buf g2(n10[2], n9[2]);
    buf g3(n10[3], n9[3]);
    buf g4(n10[4], n9[4]);
    buf g5(n10[5], n9[5]);
    buf g6(n10[6], n9[6]);
    buf g7(n10[7], n9[7]);
    dff g8(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n171), .Q(n12));
    dff g9(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n170), .Q(n13));
    or g10(n171 ,n169 ,n168);
    nor g11(n170 ,n169 ,n167);
    or g12(n168 ,n30 ,n166);
    nor g13(n167 ,n29 ,n165);
    nor g14(n166 ,n164 ,n163);
    nor g15(n165 ,n164 ,n162);
    or g16(n163 ,n143 ,n161);
    dff g17(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n160), .Q(n11));
    or g18(n162 ,n129 ,n159);
    or g19(n161 ,n112 ,n157);
    or g20(n160 ,n153 ,n158);
    or g21(n159 ,n127 ,n156);
    or g22(n158 ,n50 ,n154);
    or g23(n157 ,n118 ,n155);
    or g24(n156 ,n125 ,n150);
    dff g25(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n144), .Q(n9[1]));
    dff g26(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n152), .Q(n9[3]));
    dff g27(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n145), .Q(n9[0]));
    dff g28(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n147), .Q(n9[6]));
    dff g29(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n149), .Q(n9[4]));
    dff g30(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n151), .Q(n9[2]));
    dff g31(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n148), .Q(n9[7]));
    dff g32(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n146), .Q(n9[5]));
    or g33(n155 ,n137 ,n138);
    nor g34(n154 ,n54 ,n142);
    nor g35(n153 ,n42 ,n140);
    or g36(n152 ,n49 ,n122);
    or g37(n151 ,n45 ,n128);
    or g38(n150 ,n131 ,n133);
    or g39(n149 ,n46 ,n124);
    or g40(n148 ,n52 ,n139);
    or g41(n147 ,n44 ,n135);
    or g42(n146 ,n47 ,n136);
    or g43(n145 ,n53 ,n141);
    or g44(n144 ,n48 ,n126);
    or g45(n143 ,n117 ,n113);
    not g46(n142 ,n141);
    not g47(n140 ,n139);
    or g48(n138 ,n115 ,n114);
    or g49(n137 ,n111 ,n116);
    nor g50(n136 ,n134 ,n130);
    nor g51(n135 ,n134 ,n132);
    or g52(n133 ,n132 ,n119);
    or g53(n131 ,n123 ,n130);
    or g54(n129 ,n121 ,n120);
    nor g55(n128 ,n134 ,n127);
    nor g56(n126 ,n134 ,n125);
    nor g57(n124 ,n134 ,n123);
    nor g58(n122 ,n134 ,n121);
    nor g59(n141 ,n134 ,n120);
    nor g60(n139 ,n134 ,n119);
    not g61(n118 ,n120);
    not g62(n117 ,n127);
    not g63(n116 ,n130);
    not g64(n115 ,n132);
    not g65(n114 ,n119);
    not g66(n113 ,n121);
    not g67(n112 ,n125);
    not g68(n111 ,n123);
    nor g69(n120 ,n95 ,n110);
    nor g70(n127 ,n97 ,n109);
    nor g71(n130 ,n99 ,n107);
    nor g72(n132 ,n96 ,n106);
    nor g73(n119 ,n102 ,n105);
    nor g74(n121 ,n98 ,n104);
    nor g75(n125 ,n100 ,n103);
    nor g76(n123 ,n101 ,n108);
    or g77(n110 ,n78 ,n93);
    or g78(n109 ,n72 ,n91);
    or g79(n108 ,n71 ,n90);
    or g80(n107 ,n69 ,n88);
    or g81(n106 ,n85 ,n89);
    or g82(n105 ,n62 ,n87);
    or g83(n104 ,n64 ,n86);
    or g84(n103 ,n81 ,n94);
    or g85(n102 ,n34 ,n66);
    or g86(n101 ,n33 ,n74);
    or g87(n100 ,n36 ,n83);
    or g88(n99 ,n35 ,n59);
    or g89(n98 ,n31 ,n65);
    or g90(n97 ,n39 ,n76);
    or g91(n96 ,n32 ,n67);
    or g92(n95 ,n38 ,n61);
    nor g93(n94 ,n77 ,n92);
    nor g94(n93 ,n82 ,n92);
    nor g95(n91 ,n80 ,n92);
    nor g96(n90 ,n63 ,n92);
    nor g97(n89 ,n68 ,n92);
    nor g98(n88 ,n70 ,n92);
    nor g99(n87 ,n84 ,n92);
    nor g100(n86 ,n73 ,n92);
    nor g101(n85 ,n84 ,n79);
    nor g102(n83 ,n82 ,n75);
    nor g103(n81 ,n80 ,n79);
    nor g104(n78 ,n77 ,n79);
    nor g105(n76 ,n77 ,n75);
    nor g106(n74 ,n73 ,n75);
    nor g107(n72 ,n73 ,n79);
    nor g108(n71 ,n70 ,n79);
    nor g109(n69 ,n68 ,n79);
    nor g110(n67 ,n70 ,n75);
    nor g111(n66 ,n68 ,n75);
    nor g112(n65 ,n80 ,n75);
    nor g113(n64 ,n63 ,n79);
    nor g114(n62 ,n60 ,n79);
    nor g115(n61 ,n60 ,n75);
    nor g116(n59 ,n63 ,n75);
    or g117(n92 ,n4 ,n58);
    or g118(n79 ,n4 ,n55);
    or g119(n75 ,n4 ,n57);
    nor g120(n58 ,n56 ,n43);
    or g121(n57 ,n56 ,n41);
    or g122(n55 ,n56 ,n54);
    nor g123(n53 ,n82 ,n51);
    nor g124(n52 ,n84 ,n51);
    nor g125(n50 ,n20 ,n51);
    nor g126(n49 ,n73 ,n51);
    nor g127(n48 ,n77 ,n51);
    nor g128(n47 ,n70 ,n51);
    nor g129(n46 ,n63 ,n51);
    nor g130(n45 ,n80 ,n51);
    nor g131(n44 ,n68 ,n51);
    nor g132(n43 ,n42 ,n40);
    not g133(n41 ,n40);
    not g134(n54 ,n42);
    nor g135(n39 ,n37 ,n27);
    nor g136(n38 ,n37 ,n28);
    nor g137(n36 ,n37 ,n22);
    nor g138(n35 ,n37 ,n24);
    nor g139(n34 ,n37 ,n19);
    nor g140(n42 ,n17 ,n7[1]);
    or g141(n134 ,n169 ,n164);
    nor g142(n33 ,n37 ,n15);
    nor g143(n32 ,n37 ,n18);
    nor g144(n31 ,n37 ,n23);
    nor g145(n30 ,n14 ,n2);
    nor g146(n29 ,n16 ,n2);
    nor g147(n40 ,n21 ,n7[0]);
    or g148(n60 ,n25 ,n26);
    or g149(n51 ,n169 ,n2);
    not g150(n28 ,n8[0]);
    not g151(n27 ,n8[2]);
    not g152(n26 ,n6);
    not g153(n25 ,n5);
    not g154(n84 ,n9[7]);
    not g155(n82 ,n9[0]);
    not g156(n56 ,n3);
    not g157(n73 ,n9[3]);
    not g158(n77 ,n9[1]);
    not g159(n169 ,n1);
    not g160(n70 ,n9[5]);
    not g161(n80 ,n9[2]);
    not g162(n37 ,n4);
    not g163(n24 ,n8[5]);
    not g164(n23 ,n8[3]);
    not g165(n22 ,n8[1]);
    not g166(n21 ,n7[1]);
    not g167(n20 ,n11);
    not g168(n19 ,n8[7]);
    not g169(n18 ,n8[6]);
    not g170(n17 ,n7[0]);
    not g171(n16 ,n13);
    not g172(n15 ,n8[4]);
    not g173(n14 ,n12);
    not g174(n164 ,n2);
    not g175(n68 ,n9[6]);
    not g176(n63 ,n9[4]);
endmodule
