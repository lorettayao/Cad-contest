module top(n0, n1, n2, n3, n4, n5);
    input n0, n1;
    input [127:0] n2;
    output [63:0] n3, n4, n5;
    wire n0, n1;
    wire [127:0] n2;
    wire [63:0] n3, n4, n5;
    wire [2:0] n6;
    wire [15:0] n7;
    wire [7:0] n8;
    wire n9, n10, n11, n12, n13, n14, n15, n16;
    wire n17, n18, n19, n20, n21, n22, n23, n24;
    wire n25, n26, n27, n28, n29, n30, n31, n32;
    wire n33, n34, n35, n36, n37, n38, n39, n40;
    wire n41, n42, n43, n44, n45, n46, n47, n48;
    wire n49, n50, n51, n52, n53, n54, n55, n56;
    wire n57, n58, n59, n60, n61, n62, n63, n64;
    wire n65, n66, n67, n68, n69, n70, n71, n72;
    wire n73, n74, n75, n76, n77, n78, n79, n80;
    wire n81, n82, n83, n84, n85, n86, n87, n88;
    wire n89, n90, n91, n92, n93, n94, n95, n96;
    wire n97, n98, n99, n100, n101, n102, n103, n104;
    wire n105, n106, n107, n108, n109, n110, n111, n112;
    wire n113, n114, n115, n116, n117, n118, n119, n120;
    wire n121, n122, n123, n124, n125, n126, n127, n128;
    wire n129, n130, n131, n132, n133, n134, n135, n136;
    wire n137, n138, n139, n140, n141, n142, n143, n144;
    wire n145, n146, n147, n148, n149, n150, n151, n152;
    wire n153, n154, n155, n156, n157, n158, n159, n160;
    wire n161, n162, n163, n164, n165, n166, n167, n168;
    wire n169, n170, n171, n172, n173, n174, n175, n176;
    wire n177, n178, n179, n180, n181, n182, n183, n184;
    wire n185, n186, n187, n188, n189, n190, n191, n192;
    wire n193, n194, n195, n196, n197, n198, n199, n200;
    wire n201, n202, n203, n204, n205, n206, n207, n208;
    wire n209, n210, n211, n212, n213, n214, n215, n216;
    wire n217, n218, n219, n220, n221, n222, n223, n224;
    wire n225, n226, n227, n228, n229, n230, n231, n232;
    wire n233, n234, n235, n236, n237, n238, n239, n240;
    wire n241, n242, n243, n244, n245, n246, n247, n248;
    wire n249, n250, n251, n252, n253, n254, n255, n256;
    wire n257, n258, n259, n260, n261, n262, n263, n264;
    wire n265, n266, n267, n268, n269, n270, n271, n272;
    wire n273, n274, n275, n276, n277, n278, n279, n280;
    wire n281, n282, n283, n284, n285, n286, n287, n288;
    wire n289, n290, n291, n292, n293, n294, n295, n296;
    wire n297, n298, n299, n300, n301, n302, n303, n304;
    wire n305, n306, n307, n308, n309, n310, n311, n312;
    wire n313, n314, n315, n316, n317, n318, n319, n320;
    wire n321, n322, n323, n324, n325, n326, n327, n328;
    wire n329, n330, n331, n332, n333, n334, n335, n336;
    wire n337, n338, n339, n340, n341, n342, n343, n344;
    wire n345, n346, n347, n348, n349, n350, n351, n352;
    wire n353, n354, n355, n356, n357, n358, n359, n360;
    wire n361, n362, n363, n364, n365, n366, n367, n368;
    wire n369, n370, n371, n372, n373, n374, n375, n376;
    wire n377, n378, n379, n380, n381, n382, n383, n384;
    wire n385, n386, n387, n388, n389, n390, n391, n392;
    wire n393, n394, n395, n396, n397, n398, n399, n400;
    wire n401, n402, n403, n404, n405, n406, n407, n408;
    wire n409, n410, n411, n412, n413, n414, n415, n416;
    wire n417, n418, n419, n420, n421, n422, n423, n424;
    wire n425, n426, n427, n428, n429, n430, n431, n432;
    wire n433, n434, n435, n436, n437, n438, n439, n440;
    wire n441, n442, n443, n444, n445, n446, n447, n448;
    wire n449, n450, n451, n452, n453, n454, n455, n456;
    wire n457, n458, n459, n460, n461, n462, n463, n464;
    wire n465, n466, n467, n468, n469, n470, n471, n472;
    wire n473, n474, n475, n476, n477, n478, n479, n480;
    wire n481, n482, n483, n484, n485, n486, n487, n488;
    wire n489, n490, n491, n492, n493, n494, n495, n496;
    wire n497, n498, n499, n500, n501, n502, n503, n504;
    wire n505, n506, n507, n508, n509, n510, n511, n512;
    wire n513, n514, n515, n516, n517, n518, n519, n520;
    wire n521, n522, n523, n524, n525, n526, n527, n528;
    wire n529, n530, n531, n532, n533, n534, n535, n536;
    wire n537, n538, n539, n540, n541, n542, n543, n544;
    wire n545, n546, n547, n548, n549, n550, n551, n552;
    wire n553, n554, n555, n556, n557, n558, n559, n560;
    wire n561, n562, n563, n564, n565, n566, n567, n568;
    wire n569, n570, n571, n572, n573, n574, n575, n576;
    wire n577, n578, n579, n580, n581, n582, n583, n584;
    wire n585, n586, n587, n588, n589, n590, n591, n592;
    wire n593, n594, n595, n596, n597, n598, n599, n600;
    wire n601, n602, n603, n604, n605, n606, n607, n608;
    wire n609, n610, n611, n612, n613, n614, n615, n616;
    wire n617, n618, n619, n620, n621, n622, n623, n624;
    wire n625, n626, n627, n628, n629, n630, n631, n632;
    wire n633, n634, n635, n636, n637, n638, n639, n640;
    wire n641, n642, n643, n644, n645, n646, n647, n648;
    wire n649, n650, n651, n652, n653, n654, n655, n656;
    wire n657, n658, n659, n660, n661, n662, n663, n664;
    wire n665, n666, n667, n668, n669, n670, n671, n672;
    wire n673, n674, n675, n676, n677, n678, n679, n680;
    wire n681, n682, n683, n684, n685, n686, n687, n688;
    wire n689, n690, n691, n692, n693, n694, n695, n696;
    wire n697, n698, n699, n700, n701, n702, n703, n704;
    wire n705, n706, n707, n708, n709, n710, n711, n712;
    wire n713, n714, n715, n716, n717, n718, n719, n720;
    wire n721, n722, n723, n724, n725, n726, n727, n728;
    wire n729, n730, n731, n732, n733, n734, n735, n736;
    wire n737, n738, n739, n740, n741, n742, n743, n744;
    wire n745, n746, n747, n748, n749, n750, n751, n752;
    wire n753, n754, n755, n756, n757, n758, n759, n760;
    wire n761, n762, n763, n764, n765, n766, n767, n768;
    wire n769, n770, n771, n772, n773, n774, n775, n776;
    wire n777, n778, n779, n780, n781, n782, n783, n784;
    wire n785, n786, n787, n788, n789, n790, n791, n792;
    wire n793, n794, n795, n796, n797, n798, n799, n800;
    wire n801, n802, n803, n804, n805, n806, n807, n808;
    wire n809, n810, n811, n812, n813, n814, n815, n816;
    wire n817, n818, n819, n820, n821, n822, n823, n824;
    wire n825, n826, n827, n828, n829, n830, n831, n832;
    wire n833, n834, n835, n836, n837, n838, n839, n840;
    wire n841, n842, n843, n844, n845, n846, n847, n848;
    wire n849, n850, n851, n852, n853, n854, n855, n856;
    wire n857, n858, n859, n860, n861, n862, n863, n864;
    wire n865, n866, n867, n868, n869, n870, n871, n872;
    wire n873, n874, n875, n876, n877, n878, n879, n880;
    wire n881, n882, n883, n884, n885, n886, n887, n888;
    wire n889, n890, n891, n892, n893, n894, n895, n896;
    wire n897, n898, n899, n900, n901, n902, n903, n904;
    wire n905, n906, n907, n908, n909, n910, n911, n912;
    wire n913, n914, n915, n916, n917, n918, n919, n920;
    wire n921, n922, n923, n924, n925, n926, n927, n928;
    wire n929, n930, n931, n932, n933, n934, n935, n936;
    wire n937, n938, n939, n940, n941, n942, n943, n944;
    wire n945, n946, n947, n948, n949, n950, n951, n952;
    wire n953, n954, n955, n956, n957, n958, n959, n960;
    wire n961, n962, n963, n964, n965, n966, n967, n968;
    wire n969, n970, n971, n972, n973, n974, n975, n976;
    wire n977, n978, n979, n980, n981, n982, n983, n984;
    wire n985, n986, n987, n988, n989, n990, n991, n992;
    wire n993, n994, n995, n996, n997, n998, n999, n1000;
    wire n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008;
    wire n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016;
    wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
    wire n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
    wire n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
    wire n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
    wire n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056;
    wire n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064;
    wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
    wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
    wire n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088;
    wire n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096;
    wire n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104;
    wire n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112;
    wire n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120;
    wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
    wire n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136;
    wire n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
    wire n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152;
    wire n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160;
    wire n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168;
    wire n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176;
    wire n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184;
    wire n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192;
    wire n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200;
    wire n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208;
    wire n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216;
    wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
    wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
    wire n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240;
    wire n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248;
    wire n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256;
    wire n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264;
    wire n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
    wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
    wire n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288;
    wire n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296;
    wire n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304;
    wire n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312;
    wire n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320;
    wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
    wire n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
    wire n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344;
    wire n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352;
    wire n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360;
    wire n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368;
    wire n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376;
    wire n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384;
    wire n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392;
    wire n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400;
    wire n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408;
    wire n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416;
    wire n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424;
    wire n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432;
    wire n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440;
    wire n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448;
    wire n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456;
    wire n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464;
    wire n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472;
    wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480;
    wire n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488;
    wire n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496;
    wire n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504;
    wire n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512;
    wire n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520;
    wire n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528;
    wire n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536;
    wire n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544;
    wire n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552;
    wire n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560;
    wire n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568;
    wire n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576;
    wire n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584;
    wire n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592;
    wire n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600;
    wire n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608;
    wire n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616;
    wire n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624;
    wire n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632;
    wire n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640;
    wire n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648;
    wire n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656;
    wire n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664;
    wire n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672;
    wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
    wire n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688;
    wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
    wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
    wire n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712;
    wire n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720;
    wire n1721, n1722, n1723, n1724, n1725;
    buf g0(n5[16], 1'b0);
    buf g1(n5[17], 1'b0);
    buf g2(n5[18], 1'b0);
    buf g3(n5[19], 1'b0);
    buf g4(n5[20], 1'b0);
    buf g5(n5[21], 1'b0);
    buf g6(n5[22], 1'b0);
    buf g7(n5[23], 1'b0);
    buf g8(n5[24], 1'b0);
    buf g9(n5[25], 1'b0);
    buf g10(n5[26], 1'b0);
    buf g11(n5[27], 1'b0);
    buf g12(n5[28], 1'b0);
    buf g13(n5[29], 1'b0);
    buf g14(n5[30], 1'b0);
    buf g15(n5[31], 1'b0);
    buf g16(n5[32], 1'b0);
    buf g17(n5[33], 1'b0);
    buf g18(n5[34], 1'b0);
    buf g19(n5[35], 1'b0);
    buf g20(n5[36], 1'b0);
    buf g21(n5[37], 1'b0);
    buf g22(n5[38], 1'b0);
    buf g23(n5[39], 1'b0);
    buf g24(n5[40], 1'b0);
    buf g25(n5[41], 1'b0);
    buf g26(n5[42], 1'b0);
    buf g27(n5[43], 1'b0);
    buf g28(n5[44], 1'b0);
    buf g29(n5[45], 1'b0);
    buf g30(n5[46], 1'b0);
    buf g31(n5[47], 1'b0);
    buf g32(n5[48], 1'b0);
    buf g33(n5[49], 1'b0);
    buf g34(n5[50], 1'b0);
    buf g35(n5[51], 1'b0);
    buf g36(n5[52], 1'b0);
    buf g37(n5[53], 1'b0);
    buf g38(n5[54], 1'b0);
    buf g39(n5[55], 1'b0);
    buf g40(n5[56], 1'b0);
    buf g41(n5[57], 1'b0);
    buf g42(n5[58], 1'b0);
    buf g43(n5[59], 1'b0);
    buf g44(n5[60], 1'b0);
    buf g45(n5[61], 1'b0);
    buf g46(n5[62], 1'b0);
    buf g47(n5[63], 1'b0);
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1303), .Q(n5[0]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1302), .Q(n5[1]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1301), .Q(n5[2]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1300), .Q(n5[3]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1299), .Q(n5[4]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1298), .Q(n5[5]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1297), .Q(n5[6]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1296), .Q(n5[7]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1294), .Q(n5[8]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1295), .Q(n5[9]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1293), .Q(n5[10]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1292), .Q(n5[11]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1291), .Q(n5[12]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1290), .Q(n5[13]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1289), .Q(n5[14]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1288), .Q(n5[15]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1410), .Q(n3[0]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1409), .Q(n3[1]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1408), .Q(n3[2]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1407), .Q(n3[3]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1406), .Q(n3[4]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1405), .Q(n3[5]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1403), .Q(n3[6]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1404), .Q(n3[7]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1402), .Q(n3[8]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1401), .Q(n3[9]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1400), .Q(n3[10]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1413), .Q(n3[11]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1399), .Q(n3[12]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1414), .Q(n3[13]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1412), .Q(n3[14]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1411), .Q(n3[15]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1149), .Q(n3[16]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1148), .Q(n3[17]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1147), .Q(n3[18]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1146), .Q(n3[19]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1145), .Q(n3[20]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1144), .Q(n3[21]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1143), .Q(n3[22]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1142), .Q(n3[23]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1141), .Q(n3[24]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1140), .Q(n3[25]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1139), .Q(n3[26]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1138), .Q(n3[27]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1137), .Q(n3[28]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1136), .Q(n3[29]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1135), .Q(n3[30]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1158), .Q(n3[31]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1159), .Q(n3[32]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1160), .Q(n3[33]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1161), .Q(n3[34]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1162), .Q(n3[35]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1163), .Q(n3[36]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1164), .Q(n3[37]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1165), .Q(n3[38]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1166), .Q(n3[39]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1167), .Q(n3[40]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1169), .Q(n3[41]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1170), .Q(n3[42]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1171), .Q(n3[43]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1172), .Q(n3[44]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1173), .Q(n3[45]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1174), .Q(n3[46]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1116), .Q(n3[47]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1115), .Q(n3[48]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1114), .Q(n3[49]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1113), .Q(n3[50]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1111), .Q(n3[51]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1110), .Q(n3[52]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1109), .Q(n3[53]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1108), .Q(n3[54]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1107), .Q(n3[55]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1106), .Q(n3[56]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1105), .Q(n3[57]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1104), .Q(n3[58]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1103), .Q(n3[59]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1102), .Q(n3[60]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1101), .Q(n3[61]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1100), .Q(n3[62]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1099), .Q(n3[63]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1098), .Q(n6[0]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1096), .Q(n6[1]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1095), .Q(n6[2]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1416), .Q(n4[0]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1430), .Q(n4[1]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1429), .Q(n4[2]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1428), .Q(n4[3]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1427), .Q(n4[4]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1426), .Q(n4[5]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1425), .Q(n4[6]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1424), .Q(n4[7]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1423), .Q(n4[8]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1422), .Q(n4[9]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1421), .Q(n4[10]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1420), .Q(n4[11]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1419), .Q(n4[12]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1418), .Q(n4[13]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1417), .Q(n4[14]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1431), .Q(n4[15]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1334), .Q(n4[16]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1333), .Q(n4[17]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1332), .Q(n4[18]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1330), .Q(n4[19]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1329), .Q(n4[20]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1328), .Q(n4[21]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1327), .Q(n4[22]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1326), .Q(n4[23]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1324), .Q(n4[24]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1323), .Q(n4[25]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1322), .Q(n4[26]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1321), .Q(n4[27]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1320), .Q(n4[28]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1319), .Q(n4[29]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1318), .Q(n4[30]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1317), .Q(n4[31]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1316), .Q(n4[32]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1314), .Q(n4[33]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1313), .Q(n4[34]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1311), .Q(n4[35]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1310), .Q(n4[36]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1309), .Q(n4[37]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1307), .Q(n4[38]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1306), .Q(n4[39]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1305), .Q(n4[40]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1304), .Q(n4[41]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1367), .Q(n4[42]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1366), .Q(n4[43]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1365), .Q(n4[44]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1364), .Q(n4[45]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1363), .Q(n4[46]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1361), .Q(n4[47]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1359), .Q(n4[48]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1358), .Q(n4[49]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1357), .Q(n4[50]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1356), .Q(n4[51]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1355), .Q(n4[52]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1354), .Q(n4[53]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1353), .Q(n4[54]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1352), .Q(n4[55]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1350), .Q(n4[56]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1349), .Q(n4[57]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1348), .Q(n4[58]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1347), .Q(n4[59]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1346), .Q(n4[60]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1345), .Q(n4[61]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1343), .Q(n4[62]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1342), .Q(n4[63]));
    or g195(n1431 ,n920 ,n1384);
    or g196(n1430 ,n1046 ,n1398);
    or g197(n1429 ,n1029 ,n1397);
    or g198(n1428 ,n1053 ,n1396);
    or g199(n1427 ,n1056 ,n1395);
    or g200(n1426 ,n939 ,n1394);
    or g201(n1425 ,n937 ,n1393);
    or g202(n1424 ,n936 ,n1392);
    or g203(n1423 ,n999 ,n1391);
    or g204(n1422 ,n932 ,n1390);
    or g205(n1421 ,n929 ,n1389);
    or g206(n1420 ,n926 ,n1388);
    or g207(n1419 ,n923 ,n1387);
    or g208(n1418 ,n897 ,n1386);
    or g209(n1417 ,n921 ,n1385);
    or g210(n1416 ,n924 ,n1415);
    or g211(n1415 ,n1216 ,n1383);
    or g212(n1414 ,n1269 ,n1351);
    or g213(n1413 ,n1283 ,n1362);
    or g214(n1412 ,n1030 ,n1344);
    or g215(n1411 ,n935 ,n1341);
    or g216(n1410 ,n1052 ,n1340);
    or g217(n1409 ,n976 ,n1339);
    or g218(n1408 ,n1244 ,n1338);
    or g219(n1407 ,n1240 ,n1337);
    or g220(n1406 ,n1235 ,n1336);
    or g221(n1405 ,n1231 ,n1335);
    or g222(n1404 ,n1219 ,n1325);
    or g223(n1403 ,n917 ,n1331);
    or g224(n1402 ,n1211 ,n1315);
    or g225(n1401 ,n1202 ,n1312);
    or g226(n1400 ,n903 ,n1308);
    or g227(n1399 ,n1027 ,n1360);
    or g228(n1398 ,n1256 ,n1382);
    or g229(n1397 ,n1255 ,n1381);
    or g230(n1396 ,n1253 ,n1380);
    or g231(n1395 ,n1252 ,n1379);
    or g232(n1394 ,n1251 ,n1378);
    or g233(n1393 ,n1248 ,n1377);
    or g234(n1392 ,n1245 ,n1376);
    or g235(n1391 ,n1243 ,n1375);
    or g236(n1390 ,n1241 ,n1374);
    or g237(n1389 ,n1239 ,n1373);
    or g238(n1388 ,n1238 ,n1372);
    or g239(n1387 ,n1236 ,n1371);
    or g240(n1386 ,n1233 ,n1370);
    or g241(n1385 ,n1230 ,n1369);
    or g242(n1384 ,n1229 ,n1368);
    nor g243(n1383 ,n505 ,n1191);
    nor g244(n1382 ,n498 ,n1190);
    nor g245(n1381 ,n508 ,n1189);
    nor g246(n1380 ,n510 ,n1188);
    nor g247(n1379 ,n509 ,n1187);
    nor g248(n1378 ,n497 ,n1186);
    nor g249(n1377 ,n511 ,n1185);
    nor g250(n1376 ,n507 ,n1184);
    nor g251(n1375 ,n501 ,n1183);
    nor g252(n1374 ,n503 ,n1182);
    nor g253(n1373 ,n496 ,n1181);
    nor g254(n1372 ,n500 ,n1180);
    nor g255(n1371 ,n499 ,n1179);
    nor g256(n1370 ,n506 ,n1178);
    nor g257(n1369 ,n504 ,n1177);
    nor g258(n1368 ,n502 ,n1176);
    or g259(n1367 ,n916 ,n1281);
    or g260(n1366 ,n1039 ,n1280);
    or g261(n1365 ,n980 ,n1279);
    or g262(n1364 ,n1037 ,n1278);
    or g263(n1363 ,n1009 ,n1276);
    or g264(n1362 ,n979 ,n1277);
    or g265(n1361 ,n1036 ,n1275);
    or g266(n1360 ,n1274 ,n1270);
    or g267(n1359 ,n1035 ,n1284);
    or g268(n1358 ,n1032 ,n1273);
    or g269(n1357 ,n1033 ,n1272);
    or g270(n1356 ,n1040 ,n1271);
    or g271(n1355 ,n938 ,n1232);
    or g272(n1354 ,n1026 ,n1268);
    or g273(n1353 ,n930 ,n1267);
    or g274(n1352 ,n1054 ,n1266);
    or g275(n1351 ,n934 ,n1265);
    or g276(n1350 ,n1057 ,n1209);
    or g277(n1349 ,n909 ,n1263);
    or g278(n1348 ,n1004 ,n1262);
    or g279(n1347 ,n1038 ,n1261);
    or g280(n1346 ,n1055 ,n1259);
    or g281(n1345 ,n892 ,n1287);
    or g282(n1344 ,n1264 ,n1260);
    or g283(n1343 ,n922 ,n1285);
    or g284(n1342 ,n1048 ,n1250);
    or g285(n1341 ,n1286 ,n1258);
    or g286(n1340 ,n1254 ,n1249);
    or g287(n1339 ,n1247 ,n1246);
    or g288(n1338 ,n933 ,n1242);
    or g289(n1337 ,n925 ,n1237);
    or g290(n1336 ,n907 ,n1234);
    or g291(n1335 ,n919 ,n1227);
    or g292(n1334 ,n918 ,n1228);
    or g293(n1333 ,n931 ,n1226);
    or g294(n1332 ,n1023 ,n1224);
    or g295(n1331 ,n1225 ,n1222);
    or g296(n1330 ,n1028 ,n1223);
    or g297(n1329 ,n1042 ,n1221);
    or g298(n1328 ,n1031 ,n1220);
    or g299(n1327 ,n915 ,n1218);
    or g300(n1326 ,n1034 ,n1217);
    or g301(n1325 ,n912 ,n1215);
    or g302(n1324 ,n913 ,n1257);
    or g303(n1323 ,n1045 ,n1214);
    or g304(n1322 ,n1044 ,n1213);
    or g305(n1321 ,n1050 ,n1212);
    or g306(n1320 ,n1051 ,n1210);
    or g307(n1319 ,n1043 ,n1208);
    or g308(n1318 ,n927 ,n1206);
    or g309(n1317 ,n1047 ,n1205);
    or g310(n1316 ,n902 ,n1204);
    or g311(n1315 ,n904 ,n1207);
    or g312(n1314 ,n911 ,n1203);
    or g313(n1313 ,n900 ,n1201);
    or g314(n1312 ,n901 ,n1199);
    or g315(n1311 ,n1041 ,n1200);
    or g316(n1310 ,n1049 ,n1198);
    or g317(n1309 ,n898 ,n1196);
    or g318(n1308 ,n1195 ,n1193);
    or g319(n1307 ,n899 ,n1197);
    or g320(n1306 ,n905 ,n1194);
    or g321(n1305 ,n910 ,n1192);
    or g322(n1304 ,n914 ,n1282);
    xor g323(n1303 ,n1119 ,n960);
    xor g324(n1302 ,n1133 ,n975);
    xor g325(n1301 ,n1120 ,n961);
    xor g326(n1300 ,n1121 ,n962);
    xor g327(n1299 ,n1122 ,n963);
    xor g328(n1298 ,n1123 ,n964);
    xor g329(n1297 ,n1124 ,n965);
    xor g330(n1296 ,n1125 ,n966);
    xor g331(n1295 ,n1127 ,n968);
    xor g332(n1294 ,n1126 ,n967);
    xor g333(n1293 ,n1128 ,n969);
    xor g334(n1292 ,n1129 ,n970);
    xor g335(n1291 ,n1130 ,n971);
    xor g336(n1290 ,n1131 ,n972);
    xor g337(n1289 ,n1132 ,n973);
    xor g338(n1288 ,n1118 ,n974);
    nor g339(n1287 ,n760 ,n495);
    nor g340(n1286 ,n502 ,n1151);
    nor g341(n1285 ,n778 ,n495);
    nor g342(n1284 ,n693 ,n495);
    nor g343(n1283 ,n653 ,n1157);
    nor g344(n1282 ,n682 ,n495);
    nor g345(n1281 ,n716 ,n495);
    nor g346(n1280 ,n743 ,n495);
    nor g347(n1279 ,n786 ,n495);
    nor g348(n1278 ,n686 ,n495);
    nor g349(n1277 ,n500 ,n1153);
    nor g350(n1276 ,n744 ,n495);
    nor g351(n1275 ,n721 ,n495);
    nor g352(n1274 ,n499 ,n1087);
    nor g353(n1273 ,n755 ,n495);
    nor g354(n1272 ,n732 ,n495);
    nor g355(n1271 ,n711 ,n495);
    nor g356(n1270 ,n667 ,n1156);
    nor g357(n1269 ,n655 ,n1155);
    nor g358(n1268 ,n723 ,n495);
    nor g359(n1267 ,n688 ,n495);
    nor g360(n1266 ,n730 ,n495);
    nor g361(n1265 ,n506 ,n1097);
    nor g362(n1264 ,n504 ,n1065);
    nor g363(n1263 ,n775 ,n495);
    nor g364(n1262 ,n758 ,n495);
    nor g365(n1261 ,n756 ,n495);
    nor g366(n1260 ,n662 ,n1070);
    nor g367(n1259 ,n678 ,n495);
    nor g368(n1258 ,n672 ,n1150);
    nor g369(n1257 ,n703 ,n495);
    nor g370(n1256 ,n647 ,n1092);
    nor g371(n1255 ,n668 ,n1152);
    nor g372(n1254 ,n505 ,n1090);
    nor g373(n1253 ,n648 ,n1091);
    nor g374(n1252 ,n671 ,n1089);
    nor g375(n1251 ,n650 ,n1086);
    nor g376(n1250 ,n772 ,n495);
    nor g377(n1249 ,n665 ,n1088);
    nor g378(n1248 ,n669 ,n1085);
    nor g379(n1247 ,n498 ,n1083);
    nor g380(n1246 ,n660 ,n1084);
    nor g381(n1245 ,n664 ,n1112);
    nor g382(n1244 ,n645 ,n1081);
    nor g383(n1243 ,n652 ,n1168);
    nor g384(n1242 ,n508 ,n1134);
    nor g385(n1241 ,n657 ,n1080);
    nor g386(n1240 ,n646 ,n1078);
    nor g387(n1239 ,n659 ,n1079);
    nor g388(n1238 ,n651 ,n1077);
    nor g389(n1237 ,n510 ,n1076);
    nor g390(n1236 ,n675 ,n1075);
    nor g391(n1235 ,n649 ,n1074);
    nor g392(n1234 ,n509 ,n1060);
    nor g393(n1233 ,n673 ,n1073);
    nor g394(n1232 ,n699 ,n495);
    nor g395(n1231 ,n654 ,n1069);
    nor g396(n1230 ,n670 ,n1072);
    nor g397(n1229 ,n663 ,n1068);
    nor g398(n1228 ,n720 ,n495);
    nor g399(n1227 ,n497 ,n1067);
    nor g400(n1226 ,n783 ,n495);
    nor g401(n1225 ,n511 ,n1154);
    nor g402(n1224 ,n725 ,n495);
    nor g403(n1223 ,n784 ,n495);
    nor g404(n1222 ,n656 ,n1064);
    nor g405(n1221 ,n729 ,n495);
    nor g406(n1220 ,n731 ,n495);
    nor g407(n1219 ,n674 ,n1066);
    nor g408(n1218 ,n761 ,n495);
    nor g409(n1217 ,n701 ,n495);
    nor g410(n1216 ,n644 ,n1093);
    nor g411(n1215 ,n507 ,n1062);
    nor g412(n1214 ,n782 ,n495);
    nor g413(n1213 ,n739 ,n495);
    nor g414(n1212 ,n780 ,n495);
    nor g415(n1211 ,n658 ,n1061);
    nor g416(n1210 ,n707 ,n495);
    nor g417(n1209 ,n750 ,n495);
    nor g418(n1208 ,n728 ,n495);
    nor g419(n1207 ,n501 ,n1082);
    nor g420(n1206 ,n702 ,n495);
    nor g421(n1205 ,n691 ,n495);
    nor g422(n1204 ,n712 ,n495);
    nor g423(n1203 ,n694 ,n495);
    nor g424(n1202 ,n666 ,n1059);
    nor g425(n1201 ,n736 ,n495);
    nor g426(n1200 ,n717 ,n495);
    nor g427(n1199 ,n503 ,n1094);
    nor g428(n1198 ,n741 ,n495);
    nor g429(n1197 ,n684 ,n495);
    nor g430(n1196 ,n765 ,n495);
    nor g431(n1195 ,n496 ,n1071);
    nor g432(n1194 ,n771 ,n495);
    nor g433(n1193 ,n661 ,n1063);
    nor g434(n1192 ,n715 ,n495);
    nor g435(n1191 ,n874 ,n1175);
    nor g436(n1190 ,n881 ,n1175);
    nor g437(n1189 ,n880 ,n1175);
    nor g438(n1188 ,n890 ,n1175);
    nor g439(n1187 ,n894 ,n1175);
    nor g440(n1186 ,n882 ,n1175);
    nor g441(n1185 ,n876 ,n1175);
    nor g442(n1184 ,n878 ,n1175);
    nor g443(n1183 ,n875 ,n1175);
    nor g444(n1182 ,n873 ,n1175);
    nor g445(n1181 ,n872 ,n1175);
    nor g446(n1180 ,n871 ,n1175);
    nor g447(n1179 ,n870 ,n1175);
    nor g448(n1178 ,n868 ,n1175);
    nor g449(n1177 ,n864 ,n1175);
    nor g450(n1176 ,n867 ,n1175);
    or g451(n1174 ,n825 ,n928);
    or g452(n1173 ,n826 ,n991);
    or g453(n1172 ,n813 ,n992);
    or g454(n1171 ,n831 ,n993);
    or g455(n1170 ,n832 ,n994);
    or g456(n1169 ,n833 ,n995);
    nor g457(n1168 ,n948 ,n940);
    or g458(n1167 ,n834 ,n996);
    or g459(n1166 ,n835 ,n997);
    or g460(n1165 ,n836 ,n998);
    or g461(n1164 ,n837 ,n1000);
    or g462(n1163 ,n838 ,n1001);
    or g463(n1162 ,n839 ,n1002);
    or g464(n1161 ,n840 ,n1005);
    or g465(n1160 ,n841 ,n1006);
    or g466(n1159 ,n842 ,n1007);
    or g467(n1158 ,n843 ,n1008);
    nor g468(n1157 ,n944 ,n942);
    nor g469(n1156 ,n957 ,n942);
    nor g470(n1155 ,n949 ,n942);
    nor g471(n1154 ,n795 ,n866);
    nor g472(n1153 ,n795 ,n889);
    nor g473(n1152 ,n946 ,n940);
    nor g474(n1151 ,n795 ,n888);
    nor g475(n1150 ,n952 ,n942);
    or g476(n1149 ,n845 ,n1025);
    or g477(n1148 ,n858 ,n1024);
    or g478(n1147 ,n857 ,n1022);
    or g479(n1146 ,n856 ,n1021);
    or g480(n1145 ,n855 ,n1020);
    or g481(n1144 ,n854 ,n1019);
    or g482(n1143 ,n853 ,n1018);
    or g483(n1142 ,n852 ,n1017);
    or g484(n1141 ,n851 ,n1016);
    or g485(n1140 ,n850 ,n1015);
    or g486(n1139 ,n849 ,n1014);
    or g487(n1138 ,n847 ,n1013);
    or g488(n1137 ,n846 ,n1011);
    or g489(n1136 ,n859 ,n1010);
    or g490(n1135 ,n844 ,n1058);
    nor g491(n1134 ,n795 ,n886);
    nor g492(n1133 ,n498 ,n943);
    nor g493(n1132 ,n504 ,n943);
    nor g494(n1131 ,n506 ,n943);
    nor g495(n1130 ,n499 ,n943);
    nor g496(n1129 ,n500 ,n943);
    nor g497(n1128 ,n496 ,n943);
    nor g498(n1127 ,n503 ,n943);
    nor g499(n1126 ,n501 ,n943);
    nor g500(n1125 ,n507 ,n943);
    nor g501(n1124 ,n511 ,n943);
    nor g502(n1123 ,n497 ,n943);
    nor g503(n1122 ,n509 ,n943);
    nor g504(n1121 ,n510 ,n943);
    nor g505(n1120 ,n508 ,n943);
    nor g506(n1119 ,n505 ,n943);
    nor g507(n1118 ,n502 ,n943);
    nor g508(n1175 ,n940 ,n941);
    not g509(n495 ,n1117);
    or g510(n1116 ,n824 ,n990);
    or g511(n1115 ,n823 ,n989);
    or g512(n1114 ,n822 ,n988);
    or g513(n1113 ,n848 ,n1003);
    nor g514(n1112 ,n953 ,n940);
    or g515(n1111 ,n820 ,n987);
    or g516(n1110 ,n819 ,n986);
    or g517(n1109 ,n818 ,n985);
    or g518(n1108 ,n821 ,n984);
    or g519(n1107 ,n816 ,n983);
    or g520(n1106 ,n815 ,n1012);
    or g521(n1105 ,n814 ,n982);
    or g522(n1104 ,n809 ,n896);
    or g523(n1103 ,n827 ,n981);
    or g524(n1102 ,n812 ,n908);
    or g525(n1101 ,n817 ,n906);
    or g526(n1100 ,n810 ,n978);
    or g527(n1099 ,n811 ,n977);
    nor g528(n1098 ,n1 ,n895);
    nor g529(n1097 ,n795 ,n883);
    nor g530(n1096 ,n1 ,n861);
    nor g531(n1095 ,n1 ,n860);
    nor g532(n1094 ,n795 ,n862);
    nor g533(n1093 ,n945 ,n940);
    nor g534(n1092 ,n951 ,n940);
    nor g535(n1091 ,n959 ,n940);
    nor g536(n1090 ,n795 ,n879);
    nor g537(n1089 ,n947 ,n940);
    nor g538(n1088 ,n945 ,n942);
    nor g539(n1087 ,n795 ,n891);
    nor g540(n1086 ,n954 ,n940);
    nor g541(n1085 ,n955 ,n940);
    nor g542(n1084 ,n951 ,n942);
    nor g543(n1083 ,n795 ,n877);
    nor g544(n1082 ,n795 ,n893);
    nor g545(n1081 ,n946 ,n942);
    nor g546(n1080 ,n958 ,n940);
    nor g547(n1079 ,n950 ,n940);
    nor g548(n1078 ,n959 ,n942);
    nor g549(n1077 ,n944 ,n940);
    nor g550(n1076 ,n795 ,n885);
    nor g551(n1075 ,n957 ,n940);
    nor g552(n1074 ,n947 ,n942);
    nor g553(n1073 ,n949 ,n940);
    nor g554(n1072 ,n956 ,n940);
    nor g555(n1071 ,n795 ,n869);
    nor g556(n1070 ,n956 ,n942);
    nor g557(n1069 ,n954 ,n942);
    nor g558(n1068 ,n952 ,n940);
    nor g559(n1067 ,n795 ,n884);
    nor g560(n1066 ,n953 ,n942);
    nor g561(n1065 ,n795 ,n887);
    nor g562(n1064 ,n955 ,n942);
    nor g563(n1063 ,n950 ,n942);
    nor g564(n1062 ,n795 ,n865);
    nor g565(n1061 ,n948 ,n942);
    nor g566(n1060 ,n795 ,n863);
    nor g567(n1059 ,n958 ,n942);
    or g568(n1117 ,n829 ,n940);
    nor g569(n1058 ,n614 ,n491);
    nor g570(n1057 ,n539 ,n491);
    nor g571(n1056 ,n532 ,n494);
    nor g572(n1055 ,n543 ,n494);
    nor g573(n1054 ,n537 ,n491);
    nor g574(n1053 ,n583 ,n492);
    nor g575(n1052 ,n563 ,n494);
    nor g576(n1051 ,n590 ,n491);
    nor g577(n1050 ,n519 ,n491);
    nor g578(n1049 ,n591 ,n491);
    nor g579(n1048 ,n569 ,n494);
    nor g580(n1047 ,n606 ,n491);
    nor g581(n1046 ,n615 ,n492);
    nor g582(n1045 ,n581 ,n491);
    nor g583(n1044 ,n593 ,n491);
    nor g584(n1043 ,n558 ,n494);
    nor g585(n1042 ,n624 ,n494);
    nor g586(n1041 ,n525 ,n494);
    nor g587(n1040 ,n560 ,n491);
    nor g588(n1039 ,n582 ,n494);
    nor g589(n1038 ,n586 ,n494);
    nor g590(n1037 ,n520 ,n494);
    nor g591(n1036 ,n538 ,n491);
    nor g592(n1035 ,n616 ,n494);
    nor g593(n1034 ,n630 ,n494);
    nor g594(n1033 ,n574 ,n494);
    nor g595(n1032 ,n613 ,n494);
    nor g596(n1031 ,n622 ,n491);
    nor g597(n1030 ,n553 ,n492);
    nor g598(n1029 ,n623 ,n491);
    nor g599(n1028 ,n551 ,n491);
    nor g600(n1027 ,n526 ,n492);
    nor g601(n1026 ,n545 ,n492);
    nor g602(n1025 ,n518 ,n492);
    nor g603(n1024 ,n554 ,n492);
    nor g604(n1023 ,n595 ,n492);
    nor g605(n1022 ,n603 ,n492);
    nor g606(n1021 ,n544 ,n491);
    nor g607(n1020 ,n542 ,n491);
    nor g608(n1019 ,n605 ,n491);
    nor g609(n1018 ,n598 ,n491);
    nor g610(n1017 ,n562 ,n492);
    nor g611(n1016 ,n524 ,n492);
    nor g612(n1015 ,n625 ,n492);
    nor g613(n1014 ,n632 ,n492);
    nor g614(n1013 ,n609 ,n491);
    nor g615(n1012 ,n533 ,n491);
    nor g616(n1011 ,n627 ,n492);
    nor g617(n1010 ,n637 ,n492);
    nor g618(n1009 ,n604 ,n491);
    nor g619(n1008 ,n570 ,n491);
    nor g620(n1007 ,n635 ,n491);
    nor g621(n1006 ,n588 ,n494);
    nor g622(n1005 ,n529 ,n494);
    nor g623(n1004 ,n619 ,n491);
    nor g624(n1003 ,n514 ,n494);
    nor g625(n1002 ,n528 ,n494);
    nor g626(n1001 ,n579 ,n494);
    nor g627(n1000 ,n620 ,n491);
    nor g628(n999 ,n573 ,n492);
    nor g629(n998 ,n600 ,n491);
    nor g630(n997 ,n568 ,n491);
    nor g631(n996 ,n597 ,n491);
    nor g632(n995 ,n602 ,n492);
    nor g633(n994 ,n594 ,n494);
    nor g634(n993 ,n631 ,n491);
    nor g635(n992 ,n572 ,n491);
    nor g636(n991 ,n522 ,n494);
    nor g637(n990 ,n521 ,n492);
    nor g638(n989 ,n629 ,n491);
    nor g639(n988 ,n584 ,n494);
    nor g640(n987 ,n585 ,n494);
    nor g641(n986 ,n557 ,n494);
    nor g642(n985 ,n547 ,n491);
    nor g643(n984 ,n626 ,n494);
    nor g644(n983 ,n628 ,n494);
    nor g645(n982 ,n540 ,n494);
    nor g646(n981 ,n589 ,n494);
    nor g647(n980 ,n515 ,n494);
    nor g648(n979 ,n548 ,n491);
    nor g649(n978 ,n587 ,n494);
    nor g650(n977 ,n549 ,n494);
    nor g651(n976 ,n535 ,n492);
    nor g652(n975 ,n738 ,n830);
    nor g653(n974 ,n768 ,n830);
    nor g654(n973 ,n705 ,n830);
    nor g655(n972 ,n713 ,n830);
    nor g656(n971 ,n767 ,n830);
    nor g657(n970 ,n773 ,n830);
    nor g658(n969 ,n718 ,n830);
    nor g659(n968 ,n727 ,n830);
    nor g660(n967 ,n698 ,n830);
    nor g661(n966 ,n770 ,n830);
    nor g662(n965 ,n697 ,n830);
    nor g663(n964 ,n726 ,n830);
    nor g664(n963 ,n781 ,n830);
    nor g665(n962 ,n706 ,n830);
    nor g666(n961 ,n695 ,n830);
    nor g667(n960 ,n681 ,n830);
    not g668(n941 ,n942);
    nor g669(n939 ,n575 ,n491);
    nor g670(n938 ,n556 ,n491);
    nor g671(n937 ,n611 ,n492);
    nor g672(n936 ,n571 ,n492);
    nor g673(n935 ,n566 ,n491);
    nor g674(n934 ,n607 ,n492);
    nor g675(n933 ,n567 ,n492);
    nor g676(n932 ,n634 ,n494);
    nor g677(n931 ,n552 ,n494);
    nor g678(n930 ,n536 ,n491);
    nor g679(n929 ,n612 ,n491);
    nor g680(n928 ,n565 ,n494);
    nor g681(n927 ,n530 ,n494);
    nor g682(n926 ,n576 ,n494);
    nor g683(n925 ,n617 ,n494);
    nor g684(n924 ,n592 ,n492);
    nor g685(n923 ,n601 ,n494);
    nor g686(n922 ,n559 ,n492);
    nor g687(n921 ,n513 ,n494);
    nor g688(n920 ,n527 ,n491);
    nor g689(n919 ,n578 ,n491);
    nor g690(n918 ,n618 ,n494);
    nor g691(n917 ,n555 ,n492);
    nor g692(n916 ,n561 ,n494);
    nor g693(n915 ,n633 ,n491);
    nor g694(n914 ,n550 ,n492);
    nor g695(n913 ,n636 ,n494);
    nor g696(n912 ,n608 ,n494);
    nor g697(n911 ,n639 ,n491);
    nor g698(n910 ,n599 ,n491);
    nor g699(n909 ,n523 ,n491);
    nor g700(n908 ,n640 ,n492);
    nor g701(n907 ,n610 ,n491);
    nor g702(n906 ,n541 ,n491);
    nor g703(n905 ,n621 ,n494);
    nor g704(n904 ,n534 ,n492);
    nor g705(n903 ,n577 ,n494);
    nor g706(n902 ,n546 ,n492);
    nor g707(n901 ,n638 ,n491);
    nor g708(n900 ,n531 ,n491);
    nor g709(n899 ,n517 ,n492);
    nor g710(n898 ,n596 ,n492);
    nor g711(n897 ,n580 ,n494);
    nor g712(n896 ,n516 ,n494);
    nor g713(n895 ,n807 ,n803);
    nor g714(n894 ,n4[4] ,n828);
    nor g715(n893 ,n3[8] ,n828);
    nor g716(n892 ,n564 ,n494);
    nor g717(n891 ,n3[12] ,n828);
    nor g718(n890 ,n4[3] ,n828);
    nor g719(n889 ,n3[11] ,n828);
    nor g720(n888 ,n3[15] ,n828);
    nor g721(n887 ,n3[14] ,n828);
    nor g722(n886 ,n3[2] ,n828);
    nor g723(n885 ,n3[3] ,n828);
    nor g724(n884 ,n3[5] ,n828);
    nor g725(n883 ,n3[13] ,n828);
    nor g726(n882 ,n4[5] ,n828);
    nor g727(n881 ,n4[1] ,n828);
    nor g728(n880 ,n4[2] ,n828);
    nor g729(n879 ,n3[0] ,n828);
    nor g730(n878 ,n4[7] ,n828);
    nor g731(n877 ,n3[1] ,n828);
    nor g732(n876 ,n4[6] ,n828);
    nor g733(n875 ,n4[8] ,n828);
    nor g734(n874 ,n4[0] ,n828);
    nor g735(n873 ,n4[9] ,n828);
    nor g736(n872 ,n4[10] ,n828);
    nor g737(n871 ,n4[11] ,n828);
    nor g738(n870 ,n4[12] ,n828);
    nor g739(n869 ,n3[10] ,n828);
    nor g740(n868 ,n4[13] ,n828);
    nor g741(n867 ,n4[15] ,n828);
    nor g742(n866 ,n3[6] ,n828);
    nor g743(n865 ,n3[7] ,n828);
    nor g744(n864 ,n4[14] ,n828);
    nor g745(n863 ,n3[4] ,n828);
    nor g746(n862 ,n3[9] ,n828);
    nor g747(n861 ,n806 ,n804);
    nor g748(n860 ,n805 ,n802);
    nor g749(n959 ,n7[3] ,n828);
    nor g750(n958 ,n7[9] ,n828);
    nor g751(n957 ,n7[12] ,n828);
    nor g752(n956 ,n7[14] ,n828);
    nor g753(n955 ,n7[6] ,n828);
    nor g754(n954 ,n7[5] ,n828);
    nor g755(n953 ,n7[7] ,n828);
    nor g756(n952 ,n7[15] ,n828);
    nor g757(n951 ,n7[1] ,n828);
    nor g758(n950 ,n7[10] ,n828);
    nor g759(n949 ,n7[13] ,n828);
    nor g760(n948 ,n7[8] ,n828);
    nor g761(n947 ,n7[4] ,n828);
    nor g762(n946 ,n7[2] ,n828);
    nor g763(n945 ,n7[0] ,n828);
    nor g764(n944 ,n7[11] ,n828);
    nor g765(n943 ,n800 ,n493);
    nor g766(n942 ,n794 ,n829);
    nor g767(n940 ,n1 ,n808);
    nor g768(n859 ,n757 ,n794);
    nor g769(n858 ,n692 ,n794);
    nor g770(n857 ,n774 ,n794);
    nor g771(n856 ,n719 ,n794);
    nor g772(n855 ,n766 ,n794);
    nor g773(n854 ,n690 ,n794);
    nor g774(n853 ,n748 ,n794);
    nor g775(n852 ,n776 ,n794);
    nor g776(n851 ,n737 ,n794);
    nor g777(n850 ,n733 ,n794);
    nor g778(n849 ,n700 ,n794);
    nor g779(n848 ,n708 ,n794);
    nor g780(n847 ,n745 ,n794);
    nor g781(n846 ,n752 ,n794);
    nor g782(n845 ,n753 ,n794);
    nor g783(n844 ,n749 ,n794);
    nor g784(n843 ,n754 ,n794);
    nor g785(n842 ,n764 ,n794);
    nor g786(n841 ,n740 ,n794);
    nor g787(n840 ,n735 ,n794);
    nor g788(n839 ,n759 ,n794);
    nor g789(n838 ,n742 ,n794);
    nor g790(n837 ,n762 ,n794);
    nor g791(n836 ,n679 ,n794);
    nor g792(n835 ,n763 ,n794);
    nor g793(n834 ,n710 ,n794);
    nor g794(n833 ,n714 ,n794);
    nor g795(n832 ,n709 ,n794);
    nor g796(n831 ,n769 ,n794);
    not g797(n828 ,n829);
    not g798(n491 ,n493);
    not g799(n492 ,n493);
    not g800(n493 ,n494);
    nor g801(n827 ,n724 ,n794);
    nor g802(n826 ,n704 ,n794);
    nor g803(n825 ,n680 ,n794);
    nor g804(n824 ,n779 ,n794);
    nor g805(n823 ,n777 ,n794);
    nor g806(n822 ,n683 ,n794);
    nor g807(n821 ,n734 ,n794);
    nor g808(n820 ,n677 ,n794);
    nor g809(n819 ,n676 ,n794);
    nor g810(n818 ,n512 ,n794);
    nor g811(n817 ,n685 ,n794);
    nor g812(n816 ,n746 ,n794);
    nor g813(n815 ,n785 ,n794);
    nor g814(n814 ,n696 ,n794);
    nor g815(n813 ,n722 ,n794);
    nor g816(n812 ,n689 ,n794);
    nor g817(n811 ,n751 ,n794);
    nor g818(n810 ,n747 ,n794);
    nor g819(n809 ,n687 ,n794);
    nor g820(n808 ,n789 ,n797);
    nor g821(n807 ,n643 ,n796);
    nor g822(n806 ,n641 ,n796);
    nor g823(n804 ,n797 ,n793);
    or g824(n830 ,n1 ,n799);
    nor g825(n829 ,n643 ,n801);
    or g826(n494 ,n1 ,n798);
    not g827(n801 ,n800);
    nor g828(n799 ,n641 ,n790);
    or g829(n798 ,n642 ,n788);
    nor g830(n800 ,n641 ,n791);
    not g831(n796 ,n797);
    or g832(n793 ,n792 ,n787);
    nor g833(n797 ,n642 ,n787);
    nor g834(n795 ,n788 ,n791);
    or g835(n794 ,n1 ,n787);
    nor g836(n792 ,n643 ,n641);
    or g837(n791 ,n6[2] ,n1);
    not g838(n790 ,n789);
    not g839(n788 ,n787);
    nor g840(n789 ,n6[0] ,n6[2]);
    nor g841(n787 ,n6[0] ,n6[1]);
    not g842(n786 ,n4[44]);
    not g843(n785 ,n3[56]);
    not g844(n784 ,n4[19]);
    not g845(n783 ,n4[17]);
    not g846(n782 ,n4[25]);
    not g847(n781 ,n5[4]);
    not g848(n780 ,n4[27]);
    not g849(n779 ,n3[47]);
    not g850(n778 ,n4[62]);
    not g851(n777 ,n3[48]);
    not g852(n776 ,n3[23]);
    not g853(n775 ,n4[57]);
    not g854(n774 ,n3[18]);
    not g855(n773 ,n5[11]);
    not g856(n772 ,n4[63]);
    not g857(n771 ,n4[39]);
    not g858(n770 ,n5[7]);
    not g859(n769 ,n3[43]);
    not g860(n768 ,n5[15]);
    not g861(n767 ,n5[12]);
    not g862(n766 ,n3[20]);
    not g863(n765 ,n4[37]);
    not g864(n764 ,n3[32]);
    not g865(n763 ,n3[39]);
    not g866(n762 ,n3[37]);
    not g867(n761 ,n4[22]);
    not g868(n760 ,n4[61]);
    not g869(n759 ,n3[35]);
    not g870(n758 ,n4[58]);
    not g871(n757 ,n3[29]);
    not g872(n756 ,n4[59]);
    not g873(n755 ,n4[49]);
    not g874(n754 ,n3[31]);
    not g875(n753 ,n3[16]);
    not g876(n752 ,n3[28]);
    not g877(n751 ,n3[63]);
    not g878(n750 ,n4[56]);
    not g879(n749 ,n3[30]);
    not g880(n748 ,n3[22]);
    not g881(n747 ,n3[62]);
    not g882(n746 ,n3[55]);
    not g883(n745 ,n3[27]);
    not g884(n744 ,n4[46]);
    not g885(n743 ,n4[43]);
    not g886(n742 ,n3[36]);
    not g887(n741 ,n4[36]);
    not g888(n740 ,n3[33]);
    not g889(n739 ,n4[26]);
    not g890(n738 ,n5[1]);
    not g891(n737 ,n3[24]);
    not g892(n736 ,n4[34]);
    not g893(n735 ,n3[34]);
    not g894(n734 ,n3[54]);
    not g895(n733 ,n3[25]);
    not g896(n732 ,n4[50]);
    not g897(n731 ,n4[21]);
    not g898(n730 ,n4[55]);
    not g899(n729 ,n4[20]);
    not g900(n728 ,n4[29]);
    not g901(n727 ,n5[9]);
    not g902(n726 ,n5[5]);
    not g903(n725 ,n4[18]);
    not g904(n724 ,n3[59]);
    not g905(n723 ,n4[53]);
    not g906(n722 ,n3[44]);
    not g907(n721 ,n4[47]);
    not g908(n720 ,n4[16]);
    not g909(n719 ,n3[19]);
    not g910(n718 ,n5[10]);
    not g911(n717 ,n4[35]);
    not g912(n716 ,n4[42]);
    not g913(n715 ,n4[40]);
    not g914(n714 ,n3[41]);
    not g915(n713 ,n5[13]);
    not g916(n712 ,n4[32]);
    not g917(n711 ,n4[51]);
    not g918(n710 ,n3[40]);
    not g919(n709 ,n3[42]);
    not g920(n708 ,n3[50]);
    not g921(n707 ,n4[28]);
    not g922(n706 ,n5[3]);
    not g923(n705 ,n5[14]);
    not g924(n704 ,n3[45]);
    not g925(n703 ,n4[24]);
    not g926(n702 ,n4[30]);
    not g927(n701 ,n4[23]);
    not g928(n700 ,n3[26]);
    not g929(n699 ,n4[52]);
    not g930(n698 ,n5[8]);
    not g931(n697 ,n5[6]);
    not g932(n696 ,n3[57]);
    not g933(n695 ,n5[2]);
    not g934(n694 ,n4[33]);
    not g935(n693 ,n4[48]);
    not g936(n692 ,n3[17]);
    not g937(n691 ,n4[31]);
    not g938(n690 ,n3[21]);
    not g939(n689 ,n3[60]);
    not g940(n688 ,n4[54]);
    not g941(n687 ,n3[58]);
    not g942(n686 ,n4[45]);
    not g943(n685 ,n3[61]);
    not g944(n684 ,n4[38]);
    not g945(n683 ,n3[49]);
    not g946(n682 ,n4[41]);
    not g947(n681 ,n5[0]);
    not g948(n680 ,n3[46]);
    not g949(n679 ,n3[38]);
    not g950(n678 ,n4[60]);
    not g951(n677 ,n3[51]);
    not g952(n676 ,n3[52]);
    not g953(n675 ,n4[12]);
    not g954(n674 ,n3[7]);
    not g955(n673 ,n4[13]);
    not g956(n672 ,n3[15]);
    not g957(n671 ,n4[4]);
    not g958(n670 ,n4[14]);
    not g959(n669 ,n4[6]);
    not g960(n668 ,n4[2]);
    not g961(n667 ,n3[12]);
    not g962(n666 ,n3[9]);
    not g963(n665 ,n3[0]);
    not g964(n664 ,n4[7]);
    not g965(n663 ,n4[15]);
    not g966(n662 ,n3[14]);
    not g967(n661 ,n3[10]);
    not g968(n660 ,n3[1]);
    not g969(n659 ,n4[10]);
    not g970(n658 ,n3[8]);
    not g971(n657 ,n4[9]);
    not g972(n656 ,n3[6]);
    not g973(n655 ,n3[13]);
    not g974(n654 ,n3[5]);
    not g975(n653 ,n3[11]);
    not g976(n652 ,n4[8]);
    not g977(n651 ,n4[11]);
    not g978(n650 ,n4[5]);
    not g979(n649 ,n3[4]);
    not g980(n648 ,n4[3]);
    not g981(n647 ,n4[1]);
    not g982(n646 ,n3[3]);
    not g983(n645 ,n3[2]);
    not g984(n644 ,n4[0]);
    not g985(n643 ,n6[0]);
    not g986(n642 ,n6[2]);
    not g987(n641 ,n6[1]);
    not g988(n640 ,n1556);
    not g989(n639 ,n1465);
    not g990(n638 ,n1505);
    not g991(n637 ,n1525);
    not g992(n636 ,n1456);
    not g993(n635 ,n1528);
    not g994(n634 ,n1441);
    not g995(n633 ,n1454);
    not g996(n632 ,n1522);
    not g997(n631 ,n1539);
    not g998(n630 ,n1455);
    not g999(n629 ,n1544);
    not g1000(n628 ,n1551);
    not g1001(n627 ,n1524);
    not g1002(n626 ,n1550);
    not g1003(n625 ,n1521);
    not g1004(n624 ,n1452);
    not g1005(n623 ,n1434);
    not g1006(n622 ,n1453);
    not g1007(n621 ,n1471);
    not g1008(n620 ,n1533);
    not g1009(n619 ,n1490);
    not g1010(n618 ,n1448);
    not g1011(n617 ,n1499);
    not g1012(n616 ,n1480);
    not g1013(n615 ,n1433);
    not g1014(n614 ,n1526);
    not g1015(n613 ,n1481);
    not g1016(n612 ,n1442);
    not g1017(n611 ,n1438);
    not g1018(n610 ,n1500);
    not g1019(n609 ,n1523);
    not g1020(n608 ,n1503);
    not g1021(n607 ,n1509);
    not g1022(n606 ,n1463);
    not g1023(n605 ,n1517);
    not g1024(n604 ,n1478);
    not g1025(n603 ,n1514);
    not g1026(n602 ,n1537);
    not g1027(n601 ,n1444);
    not g1028(n600 ,n1534);
    not g1029(n599 ,n1472);
    not g1030(n598 ,n1518);
    not g1031(n597 ,n1536);
    not g1032(n596 ,n1469);
    not g1033(n595 ,n1450);
    not g1034(n594 ,n1538);
    not g1035(n593 ,n1458);
    not g1036(n592 ,n1432);
    not g1037(n591 ,n1468);
    not g1038(n590 ,n1460);
    not g1039(n589 ,n1555);
    not g1040(n588 ,n1529);
    not g1041(n587 ,n1558);
    not g1042(n586 ,n1491);
    not g1043(n585 ,n1547);
    not g1044(n584 ,n1545);
    not g1045(n583 ,n1435);
    not g1046(n582 ,n1475);
    not g1047(n581 ,n1457);
    not g1048(n580 ,n1445);
    not g1049(n579 ,n1532);
    not g1050(n578 ,n1501);
    not g1051(n577 ,n1506);
    not g1052(n576 ,n1443);
    not g1053(n575 ,n1437);
    not g1054(n574 ,n1482);
    not g1055(n573 ,n1440);
    not g1056(n572 ,n1540);
    not g1057(n571 ,n1439);
    not g1058(n570 ,n1527);
    not g1059(n569 ,n1495);
    not g1060(n568 ,n1535);
    not g1061(n567 ,n1498);
    not g1062(n566 ,n1511);
    not g1063(n565 ,n1542);
    not g1064(n564 ,n1493);
    not g1065(n563 ,n1496);
    not g1066(n562 ,n1519);
    not g1067(n561 ,n1474);
    not g1068(n560 ,n1483);
    not g1069(n559 ,n1494);
    not g1070(n558 ,n1461);
    not g1071(n557 ,n1548);
    not g1072(n556 ,n1484);
    not g1073(n555 ,n1502);
    not g1074(n554 ,n1513);
    not g1075(n553 ,n1510);
    not g1076(n552 ,n1449);
    not g1077(n551 ,n1451);
    not g1078(n550 ,n1473);
    not g1079(n549 ,n1559);
    not g1080(n548 ,n1507);
    not g1081(n547 ,n1549);
    not g1082(n546 ,n1464);
    not g1083(n545 ,n1485);
    not g1084(n544 ,n1515);
    not g1085(n543 ,n1492);
    not g1086(n542 ,n1516);
    not g1087(n541 ,n1557);
    not g1088(n540 ,n1553);
    not g1089(n539 ,n1488);
    not g1090(n538 ,n1479);
    not g1091(n537 ,n1487);
    not g1092(n536 ,n1486);
    not g1093(n535 ,n1497);
    not g1094(n534 ,n1504);
    not g1095(n533 ,n1552);
    not g1096(n532 ,n1436);
    not g1097(n531 ,n1466);
    not g1098(n530 ,n1462);
    not g1099(n529 ,n1530);
    not g1100(n528 ,n1531);
    not g1101(n527 ,n1447);
    not g1102(n526 ,n1508);
    not g1103(n525 ,n1467);
    not g1104(n524 ,n1520);
    not g1105(n523 ,n1489);
    not g1106(n522 ,n1541);
    not g1107(n521 ,n1543);
    not g1108(n520 ,n1477);
    not g1109(n519 ,n1459);
    not g1110(n518 ,n1512);
    not g1111(n517 ,n1470);
    not g1112(n516 ,n1554);
    not g1113(n515 ,n1476);
    not g1114(n514 ,n1546);
    not g1115(n513 ,n1446);
    not g1116(n512 ,n3[53]);
    not g1117(n511 ,n7[6]);
    not g1118(n510 ,n7[3]);
    not g1119(n509 ,n7[4]);
    not g1120(n508 ,n7[2]);
    not g1121(n507 ,n7[7]);
    not g1122(n506 ,n7[13]);
    not g1123(n505 ,n7[0]);
    not g1124(n504 ,n7[14]);
    not g1125(n503 ,n7[9]);
    not g1126(n502 ,n7[15]);
    not g1127(n501 ,n7[8]);
    not g1128(n500 ,n7[11]);
    not g1129(n499 ,n7[12]);
    not g1130(n498 ,n7[1]);
    not g1131(n497 ,n7[5]);
    not g1132(n496 ,n7[10]);
    xor g1133(n1559 ,n3[63] ,n304);
    nor g1134(n1558 ,n303 ,n304);
    nor g1135(n304 ,n35 ,n302);
    nor g1136(n303 ,n3[62] ,n301);
    nor g1137(n1557 ,n300 ,n301);
    not g1138(n302 ,n301);
    nor g1139(n301 ,n69 ,n299);
    nor g1140(n300 ,n3[61] ,n298);
    nor g1141(n1556 ,n297 ,n298);
    not g1142(n299 ,n298);
    nor g1143(n298 ,n45 ,n296);
    nor g1144(n297 ,n3[60] ,n295);
    nor g1145(n1555 ,n294 ,n295);
    not g1146(n296 ,n295);
    nor g1147(n295 ,n36 ,n293);
    nor g1148(n294 ,n3[59] ,n292);
    nor g1149(n1554 ,n291 ,n292);
    not g1150(n293 ,n292);
    nor g1151(n292 ,n81 ,n290);
    nor g1152(n291 ,n3[58] ,n289);
    nor g1153(n1553 ,n288 ,n289);
    not g1154(n290 ,n289);
    nor g1155(n289 ,n76 ,n287);
    nor g1156(n288 ,n3[57] ,n286);
    nor g1157(n1552 ,n285 ,n286);
    not g1158(n287 ,n286);
    nor g1159(n286 ,n34 ,n284);
    nor g1160(n285 ,n3[56] ,n283);
    nor g1161(n1551 ,n282 ,n283);
    not g1162(n284 ,n283);
    nor g1163(n283 ,n75 ,n281);
    nor g1164(n282 ,n3[55] ,n280);
    nor g1165(n1550 ,n279 ,n280);
    not g1166(n281 ,n280);
    nor g1167(n280 ,n33 ,n278);
    nor g1168(n279 ,n3[54] ,n277);
    nor g1169(n1549 ,n276 ,n277);
    not g1170(n278 ,n277);
    nor g1171(n277 ,n32 ,n275);
    nor g1172(n276 ,n3[53] ,n274);
    nor g1173(n1548 ,n273 ,n274);
    not g1174(n275 ,n274);
    nor g1175(n274 ,n40 ,n272);
    nor g1176(n273 ,n3[52] ,n271);
    nor g1177(n1547 ,n270 ,n271);
    not g1178(n272 ,n271);
    nor g1179(n271 ,n31 ,n269);
    nor g1180(n270 ,n3[51] ,n268);
    nor g1181(n1546 ,n267 ,n268);
    not g1182(n269 ,n268);
    nor g1183(n268 ,n26 ,n266);
    nor g1184(n267 ,n3[50] ,n265);
    nor g1185(n1545 ,n264 ,n265);
    not g1186(n266 ,n265);
    nor g1187(n265 ,n68 ,n263);
    nor g1188(n264 ,n3[49] ,n262);
    nor g1189(n1544 ,n261 ,n262);
    not g1190(n263 ,n262);
    nor g1191(n262 ,n48 ,n260);
    nor g1192(n261 ,n3[48] ,n259);
    nor g1193(n1543 ,n258 ,n259);
    not g1194(n260 ,n259);
    nor g1195(n259 ,n78 ,n257);
    nor g1196(n258 ,n3[47] ,n256);
    nor g1197(n1542 ,n255 ,n256);
    not g1198(n257 ,n256);
    nor g1199(n256 ,n82 ,n254);
    nor g1200(n255 ,n3[46] ,n253);
    nor g1201(n1541 ,n252 ,n253);
    not g1202(n254 ,n253);
    nor g1203(n253 ,n74 ,n251);
    nor g1204(n252 ,n3[45] ,n250);
    nor g1205(n1540 ,n249 ,n250);
    not g1206(n251 ,n250);
    nor g1207(n250 ,n22 ,n248);
    nor g1208(n249 ,n3[44] ,n247);
    nor g1209(n1539 ,n246 ,n247);
    not g1210(n248 ,n247);
    nor g1211(n247 ,n85 ,n245);
    nor g1212(n246 ,n3[43] ,n244);
    nor g1213(n1538 ,n243 ,n244);
    not g1214(n245 ,n244);
    nor g1215(n244 ,n42 ,n242);
    nor g1216(n243 ,n3[42] ,n241);
    nor g1217(n1537 ,n240 ,n241);
    not g1218(n242 ,n241);
    nor g1219(n241 ,n72 ,n239);
    nor g1220(n240 ,n3[41] ,n238);
    nor g1221(n1536 ,n237 ,n238);
    not g1222(n239 ,n238);
    nor g1223(n238 ,n25 ,n236);
    nor g1224(n237 ,n3[40] ,n235);
    nor g1225(n1535 ,n234 ,n235);
    not g1226(n236 ,n235);
    nor g1227(n235 ,n27 ,n233);
    nor g1228(n234 ,n3[39] ,n232);
    nor g1229(n1534 ,n231 ,n232);
    not g1230(n233 ,n232);
    nor g1231(n232 ,n29 ,n230);
    nor g1232(n231 ,n3[38] ,n229);
    nor g1233(n1533 ,n228 ,n229);
    not g1234(n230 ,n229);
    nor g1235(n229 ,n84 ,n227);
    nor g1236(n228 ,n3[37] ,n226);
    nor g1237(n1532 ,n225 ,n226);
    not g1238(n227 ,n226);
    nor g1239(n226 ,n47 ,n224);
    nor g1240(n225 ,n3[36] ,n223);
    nor g1241(n1531 ,n222 ,n223);
    not g1242(n224 ,n223);
    nor g1243(n223 ,n86 ,n221);
    nor g1244(n222 ,n3[35] ,n220);
    nor g1245(n1530 ,n219 ,n220);
    not g1246(n221 ,n220);
    nor g1247(n220 ,n30 ,n218);
    nor g1248(n219 ,n3[34] ,n217);
    nor g1249(n1529 ,n216 ,n217);
    not g1250(n218 ,n217);
    nor g1251(n217 ,n41 ,n215);
    nor g1252(n216 ,n3[33] ,n214);
    nor g1253(n1528 ,n213 ,n214);
    not g1254(n215 ,n214);
    nor g1255(n214 ,n87 ,n212);
    nor g1256(n213 ,n3[32] ,n211);
    nor g1257(n1527 ,n210 ,n211);
    not g1258(n212 ,n211);
    nor g1259(n211 ,n71 ,n209);
    nor g1260(n210 ,n3[31] ,n208);
    nor g1261(n1526 ,n207 ,n208);
    not g1262(n209 ,n208);
    nor g1263(n208 ,n28 ,n206);
    nor g1264(n207 ,n3[30] ,n205);
    nor g1265(n1525 ,n204 ,n205);
    not g1266(n206 ,n205);
    nor g1267(n205 ,n23 ,n203);
    nor g1268(n204 ,n3[29] ,n202);
    nor g1269(n1524 ,n201 ,n202);
    not g1270(n203 ,n202);
    nor g1271(n202 ,n43 ,n200);
    nor g1272(n201 ,n3[28] ,n199);
    nor g1273(n1523 ,n198 ,n199);
    not g1274(n200 ,n199);
    nor g1275(n199 ,n80 ,n197);
    nor g1276(n198 ,n3[27] ,n196);
    nor g1277(n1522 ,n195 ,n196);
    not g1278(n197 ,n196);
    nor g1279(n196 ,n83 ,n194);
    nor g1280(n195 ,n3[26] ,n193);
    nor g1281(n1521 ,n192 ,n193);
    not g1282(n194 ,n193);
    nor g1283(n193 ,n24 ,n191);
    nor g1284(n192 ,n3[25] ,n190);
    nor g1285(n1520 ,n189 ,n190);
    not g1286(n191 ,n190);
    nor g1287(n190 ,n37 ,n188);
    nor g1288(n189 ,n3[24] ,n187);
    nor g1289(n1519 ,n186 ,n187);
    not g1290(n188 ,n187);
    nor g1291(n187 ,n46 ,n185);
    nor g1292(n186 ,n3[23] ,n184);
    nor g1293(n1518 ,n183 ,n184);
    not g1294(n185 ,n184);
    nor g1295(n184 ,n77 ,n182);
    nor g1296(n183 ,n3[22] ,n181);
    nor g1297(n1517 ,n180 ,n181);
    not g1298(n182 ,n181);
    nor g1299(n181 ,n73 ,n179);
    nor g1300(n180 ,n3[21] ,n178);
    nor g1301(n1516 ,n177 ,n178);
    not g1302(n179 ,n178);
    nor g1303(n178 ,n70 ,n176);
    nor g1304(n177 ,n3[20] ,n175);
    nor g1305(n1515 ,n174 ,n175);
    not g1306(n176 ,n175);
    nor g1307(n175 ,n21 ,n173);
    nor g1308(n174 ,n3[19] ,n172);
    nor g1309(n1514 ,n171 ,n172);
    not g1310(n173 ,n172);
    nor g1311(n172 ,n39 ,n170);
    nor g1312(n171 ,n3[18] ,n169);
    nor g1313(n1513 ,n168 ,n169);
    not g1314(n170 ,n169);
    nor g1315(n169 ,n38 ,n167);
    nor g1316(n168 ,n3[17] ,n166);
    xnor g1317(n1512 ,n3[16] ,n165);
    not g1318(n167 ,n166);
    nor g1319(n166 ,n67 ,n165);
    nor g1320(n165 ,n112 ,n164);
    xor g1321(n1511 ,n135 ,n163);
    nor g1322(n164 ,n92 ,n163);
    nor g1323(n163 ,n110 ,n162);
    xor g1324(n1510 ,n134 ,n161);
    nor g1325(n162 ,n97 ,n161);
    nor g1326(n161 ,n108 ,n160);
    xor g1327(n1509 ,n133 ,n159);
    nor g1328(n160 ,n89 ,n159);
    nor g1329(n159 ,n106 ,n158);
    xor g1330(n1508 ,n132 ,n157);
    nor g1331(n158 ,n101 ,n157);
    nor g1332(n157 ,n118 ,n156);
    xor g1333(n1507 ,n131 ,n155);
    nor g1334(n156 ,n88 ,n155);
    nor g1335(n155 ,n116 ,n154);
    xor g1336(n1506 ,n130 ,n153);
    nor g1337(n154 ,n100 ,n153);
    nor g1338(n153 ,n115 ,n152);
    xor g1339(n1505 ,n128 ,n151);
    nor g1340(n152 ,n102 ,n151);
    nor g1341(n151 ,n117 ,n150);
    xor g1342(n1504 ,n127 ,n149);
    nor g1343(n150 ,n96 ,n149);
    nor g1344(n149 ,n105 ,n148);
    xor g1345(n1503 ,n126 ,n147);
    nor g1346(n148 ,n103 ,n147);
    nor g1347(n147 ,n104 ,n146);
    xor g1348(n1502 ,n125 ,n145);
    nor g1349(n146 ,n95 ,n145);
    nor g1350(n145 ,n113 ,n144);
    xor g1351(n1501 ,n124 ,n143);
    nor g1352(n144 ,n90 ,n143);
    nor g1353(n143 ,n107 ,n142);
    xor g1354(n1500 ,n123 ,n141);
    nor g1355(n142 ,n98 ,n141);
    nor g1356(n141 ,n109 ,n140);
    xor g1357(n1499 ,n129 ,n139);
    nor g1358(n140 ,n91 ,n139);
    nor g1359(n139 ,n111 ,n138);
    xor g1360(n1498 ,n122 ,n137);
    nor g1361(n138 ,n99 ,n137);
    xnor g1362(n1497 ,n121 ,n119);
    nor g1363(n137 ,n114 ,n136);
    nor g1364(n1496 ,n119 ,n94);
    nor g1365(n136 ,n120 ,n93);
    xnor g1366(n135 ,n7[15] ,n3[15]);
    xnor g1367(n134 ,n7[14] ,n3[14]);
    xnor g1368(n133 ,n7[13] ,n3[13]);
    xnor g1369(n132 ,n7[12] ,n3[12]);
    xnor g1370(n131 ,n7[11] ,n3[11]);
    xnor g1371(n130 ,n7[10] ,n3[10]);
    xnor g1372(n129 ,n7[3] ,n3[3]);
    xnor g1373(n128 ,n7[9] ,n3[9]);
    xnor g1374(n127 ,n7[8] ,n3[8]);
    xnor g1375(n126 ,n7[7] ,n3[7]);
    xnor g1376(n125 ,n7[6] ,n3[6]);
    xnor g1377(n124 ,n7[5] ,n3[5]);
    xnor g1378(n123 ,n7[4] ,n3[4]);
    xnor g1379(n122 ,n7[2] ,n3[2]);
    xnor g1380(n121 ,n7[1] ,n3[1]);
    not g1381(n120 ,n119);
    nor g1382(n118 ,n20 ,n18);
    nor g1383(n117 ,n59 ,n19);
    nor g1384(n116 ,n13 ,n53);
    nor g1385(n115 ,n52 ,n58);
    nor g1386(n114 ,n54 ,n16);
    nor g1387(n113 ,n15 ,n62);
    nor g1388(n112 ,n10 ,n64);
    nor g1389(n111 ,n49 ,n12);
    nor g1390(n110 ,n57 ,n9);
    nor g1391(n109 ,n65 ,n66);
    nor g1392(n108 ,n63 ,n14);
    nor g1393(n107 ,n55 ,n56);
    nor g1394(n106 ,n11 ,n61);
    nor g1395(n105 ,n60 ,n17);
    nor g1396(n104 ,n50 ,n51);
    nor g1397(n119 ,n79 ,n44);
    nor g1398(n103 ,n3[7] ,n7[7]);
    nor g1399(n102 ,n3[9] ,n7[9]);
    nor g1400(n101 ,n3[12] ,n7[12]);
    nor g1401(n100 ,n3[10] ,n7[10]);
    nor g1402(n99 ,n3[2] ,n7[2]);
    nor g1403(n98 ,n3[4] ,n7[4]);
    nor g1404(n97 ,n3[14] ,n7[14]);
    nor g1405(n96 ,n3[8] ,n7[8]);
    nor g1406(n95 ,n3[6] ,n7[6]);
    nor g1407(n94 ,n3[0] ,n7[0]);
    nor g1408(n93 ,n3[1] ,n7[1]);
    nor g1409(n92 ,n3[15] ,n7[15]);
    nor g1410(n91 ,n3[3] ,n7[3]);
    nor g1411(n90 ,n3[5] ,n7[5]);
    nor g1412(n89 ,n3[13] ,n7[13]);
    nor g1413(n88 ,n3[11] ,n7[11]);
    not g1414(n87 ,n3[32]);
    not g1415(n86 ,n3[35]);
    not g1416(n85 ,n3[43]);
    not g1417(n84 ,n3[37]);
    not g1418(n83 ,n3[26]);
    not g1419(n82 ,n3[46]);
    not g1420(n81 ,n3[58]);
    not g1421(n80 ,n3[27]);
    not g1422(n79 ,n3[0]);
    not g1423(n78 ,n3[47]);
    not g1424(n77 ,n3[22]);
    not g1425(n76 ,n3[57]);
    not g1426(n75 ,n3[55]);
    not g1427(n74 ,n3[45]);
    not g1428(n73 ,n3[21]);
    not g1429(n72 ,n3[41]);
    not g1430(n71 ,n3[31]);
    not g1431(n70 ,n3[20]);
    not g1432(n69 ,n3[61]);
    not g1433(n68 ,n3[49]);
    not g1434(n67 ,n3[16]);
    not g1435(n66 ,n7[3]);
    not g1436(n65 ,n3[3]);
    not g1437(n64 ,n7[15]);
    not g1438(n63 ,n3[13]);
    not g1439(n62 ,n7[5]);
    not g1440(n61 ,n7[12]);
    not g1441(n60 ,n3[7]);
    not g1442(n59 ,n3[8]);
    not g1443(n58 ,n7[9]);
    not g1444(n57 ,n3[14]);
    not g1445(n56 ,n7[4]);
    not g1446(n55 ,n3[4]);
    not g1447(n54 ,n3[1]);
    not g1448(n53 ,n7[10]);
    not g1449(n52 ,n3[9]);
    not g1450(n51 ,n7[6]);
    not g1451(n50 ,n3[6]);
    not g1452(n49 ,n3[2]);
    not g1453(n48 ,n3[48]);
    not g1454(n47 ,n3[36]);
    not g1455(n46 ,n3[23]);
    not g1456(n45 ,n3[60]);
    not g1457(n44 ,n7[0]);
    not g1458(n43 ,n3[28]);
    not g1459(n42 ,n3[42]);
    not g1460(n41 ,n3[33]);
    not g1461(n40 ,n3[52]);
    not g1462(n39 ,n3[18]);
    not g1463(n38 ,n3[17]);
    not g1464(n37 ,n3[24]);
    not g1465(n36 ,n3[59]);
    not g1466(n35 ,n3[62]);
    not g1467(n34 ,n3[56]);
    not g1468(n33 ,n3[54]);
    not g1469(n32 ,n3[53]);
    not g1470(n31 ,n3[51]);
    not g1471(n30 ,n3[34]);
    not g1472(n29 ,n3[38]);
    not g1473(n28 ,n3[30]);
    not g1474(n27 ,n3[39]);
    not g1475(n26 ,n3[50]);
    not g1476(n25 ,n3[40]);
    not g1477(n24 ,n3[25]);
    not g1478(n23 ,n3[29]);
    not g1479(n22 ,n3[44]);
    not g1480(n21 ,n3[19]);
    not g1481(n20 ,n3[11]);
    not g1482(n19 ,n7[8]);
    not g1483(n18 ,n7[11]);
    not g1484(n17 ,n7[7]);
    not g1485(n16 ,n7[1]);
    not g1486(n15 ,n3[5]);
    not g1487(n14 ,n7[13]);
    not g1488(n13 ,n3[10]);
    not g1489(n12 ,n7[2]);
    not g1490(n11 ,n3[12]);
    not g1491(n10 ,n3[15]);
    not g1492(n9 ,n7[14]);
    xor g1493(n1495 ,n4[63] ,n490);
    xor g1494(n1494 ,n4[62] ,n488);
    nor g1495(n490 ,n4[62] ,n489);
    xor g1496(n1493 ,n4[61] ,n486);
    not g1497(n489 ,n488);
    nor g1498(n488 ,n4[61] ,n487);
    xor g1499(n1492 ,n4[60] ,n484);
    not g1500(n487 ,n486);
    nor g1501(n486 ,n4[60] ,n485);
    xor g1502(n1491 ,n4[59] ,n482);
    not g1503(n485 ,n484);
    nor g1504(n484 ,n4[59] ,n483);
    xor g1505(n1490 ,n4[58] ,n480);
    not g1506(n483 ,n482);
    nor g1507(n482 ,n4[58] ,n481);
    xor g1508(n1489 ,n4[57] ,n478);
    not g1509(n481 ,n480);
    nor g1510(n480 ,n4[57] ,n479);
    xor g1511(n1488 ,n4[56] ,n476);
    not g1512(n479 ,n478);
    nor g1513(n478 ,n4[56] ,n477);
    xor g1514(n1487 ,n4[55] ,n474);
    not g1515(n477 ,n476);
    nor g1516(n476 ,n4[55] ,n475);
    xor g1517(n1486 ,n4[54] ,n472);
    not g1518(n475 ,n474);
    nor g1519(n474 ,n4[54] ,n473);
    xor g1520(n1485 ,n4[53] ,n470);
    not g1521(n473 ,n472);
    nor g1522(n472 ,n4[53] ,n471);
    xor g1523(n1484 ,n4[52] ,n468);
    not g1524(n471 ,n470);
    nor g1525(n470 ,n4[52] ,n469);
    xor g1526(n1483 ,n4[51] ,n466);
    not g1527(n469 ,n468);
    nor g1528(n468 ,n4[51] ,n467);
    xor g1529(n1482 ,n4[50] ,n464);
    not g1530(n467 ,n466);
    nor g1531(n466 ,n4[50] ,n465);
    xor g1532(n1481 ,n4[49] ,n462);
    not g1533(n465 ,n464);
    nor g1534(n464 ,n4[49] ,n463);
    xor g1535(n1480 ,n4[48] ,n460);
    not g1536(n463 ,n462);
    nor g1537(n462 ,n4[48] ,n461);
    xor g1538(n1479 ,n4[47] ,n458);
    not g1539(n461 ,n460);
    nor g1540(n460 ,n4[47] ,n459);
    xor g1541(n1478 ,n4[46] ,n456);
    not g1542(n459 ,n458);
    nor g1543(n458 ,n4[46] ,n457);
    xor g1544(n1477 ,n4[45] ,n454);
    not g1545(n457 ,n456);
    nor g1546(n456 ,n4[45] ,n455);
    xor g1547(n1476 ,n4[44] ,n452);
    not g1548(n455 ,n454);
    nor g1549(n454 ,n4[44] ,n453);
    xor g1550(n1475 ,n4[43] ,n450);
    not g1551(n453 ,n452);
    nor g1552(n452 ,n4[43] ,n451);
    xor g1553(n1474 ,n4[42] ,n448);
    not g1554(n451 ,n450);
    nor g1555(n450 ,n4[42] ,n449);
    xor g1556(n1473 ,n4[41] ,n446);
    not g1557(n449 ,n448);
    nor g1558(n448 ,n4[41] ,n447);
    xor g1559(n1472 ,n4[40] ,n444);
    not g1560(n447 ,n446);
    nor g1561(n446 ,n4[40] ,n445);
    xor g1562(n1471 ,n4[39] ,n442);
    not g1563(n445 ,n444);
    nor g1564(n444 ,n4[39] ,n443);
    xor g1565(n1470 ,n4[38] ,n440);
    not g1566(n443 ,n442);
    nor g1567(n442 ,n4[38] ,n441);
    xor g1568(n1469 ,n4[37] ,n438);
    not g1569(n441 ,n440);
    nor g1570(n440 ,n4[37] ,n439);
    xor g1571(n1468 ,n4[36] ,n436);
    not g1572(n439 ,n438);
    nor g1573(n438 ,n4[36] ,n437);
    xor g1574(n1467 ,n4[35] ,n434);
    not g1575(n437 ,n436);
    nor g1576(n436 ,n4[35] ,n435);
    xor g1577(n1466 ,n4[34] ,n432);
    not g1578(n435 ,n434);
    nor g1579(n434 ,n4[34] ,n433);
    xor g1580(n1465 ,n4[33] ,n430);
    not g1581(n433 ,n432);
    nor g1582(n432 ,n4[33] ,n431);
    xor g1583(n1464 ,n4[32] ,n428);
    not g1584(n431 ,n430);
    nor g1585(n430 ,n4[32] ,n429);
    xor g1586(n1463 ,n4[31] ,n426);
    not g1587(n429 ,n428);
    nor g1588(n428 ,n4[31] ,n427);
    xor g1589(n1462 ,n4[30] ,n424);
    not g1590(n427 ,n426);
    nor g1591(n426 ,n4[30] ,n425);
    xor g1592(n1461 ,n4[29] ,n422);
    not g1593(n425 ,n424);
    nor g1594(n424 ,n4[29] ,n423);
    xor g1595(n1460 ,n4[28] ,n420);
    not g1596(n423 ,n422);
    nor g1597(n422 ,n4[28] ,n421);
    xor g1598(n1459 ,n4[27] ,n418);
    not g1599(n421 ,n420);
    nor g1600(n420 ,n4[27] ,n419);
    xor g1601(n1458 ,n4[26] ,n416);
    not g1602(n419 ,n418);
    nor g1603(n418 ,n4[26] ,n417);
    xor g1604(n1457 ,n4[25] ,n414);
    not g1605(n417 ,n416);
    nor g1606(n416 ,n4[25] ,n415);
    xor g1607(n1456 ,n4[24] ,n412);
    not g1608(n415 ,n414);
    nor g1609(n414 ,n4[24] ,n413);
    xor g1610(n1455 ,n4[23] ,n410);
    not g1611(n413 ,n412);
    nor g1612(n412 ,n4[23] ,n411);
    xor g1613(n1454 ,n4[22] ,n408);
    not g1614(n411 ,n410);
    nor g1615(n410 ,n4[22] ,n409);
    xor g1616(n1453 ,n4[21] ,n406);
    not g1617(n409 ,n408);
    nor g1618(n408 ,n4[21] ,n407);
    xor g1619(n1452 ,n4[20] ,n404);
    not g1620(n407 ,n406);
    nor g1621(n406 ,n4[20] ,n405);
    xor g1622(n1451 ,n4[19] ,n402);
    not g1623(n405 ,n404);
    nor g1624(n404 ,n4[19] ,n403);
    xor g1625(n1450 ,n4[18] ,n400);
    not g1626(n403 ,n402);
    nor g1627(n402 ,n4[18] ,n401);
    xor g1628(n1449 ,n4[17] ,n398);
    not g1629(n401 ,n400);
    nor g1630(n400 ,n4[17] ,n399);
    xnor g1631(n1448 ,n4[16] ,n397);
    not g1632(n399 ,n398);
    nor g1633(n398 ,n4[16] ,n397);
    nor g1634(n397 ,n323 ,n396);
    xor g1635(n1447 ,n395 ,n344);
    nor g1636(n396 ,n345 ,n395);
    nor g1637(n395 ,n324 ,n394);
    xor g1638(n1446 ,n393 ,n346);
    nor g1639(n394 ,n347 ,n393);
    nor g1640(n393 ,n336 ,n392);
    xor g1641(n1445 ,n391 ,n350);
    nor g1642(n392 ,n351 ,n391);
    nor g1643(n391 ,n321 ,n390);
    xor g1644(n1444 ,n389 ,n358);
    nor g1645(n390 ,n359 ,n389);
    nor g1646(n389 ,n322 ,n388);
    xor g1647(n1443 ,n387 ,n338);
    nor g1648(n388 ,n339 ,n387);
    nor g1649(n387 ,n332 ,n386);
    xor g1650(n1442 ,n385 ,n340);
    nor g1651(n386 ,n341 ,n385);
    nor g1652(n385 ,n326 ,n384);
    xor g1653(n1441 ,n383 ,n342);
    nor g1654(n384 ,n343 ,n383);
    nor g1655(n383 ,n333 ,n382);
    xor g1656(n1440 ,n381 ,n362);
    nor g1657(n382 ,n363 ,n381);
    nor g1658(n381 ,n325 ,n380);
    xor g1659(n1439 ,n379 ,n348);
    nor g1660(n380 ,n349 ,n379);
    nor g1661(n379 ,n335 ,n378);
    xor g1662(n1438 ,n377 ,n364);
    nor g1663(n378 ,n365 ,n377);
    nor g1664(n377 ,n334 ,n376);
    xor g1665(n1437 ,n375 ,n360);
    nor g1666(n376 ,n361 ,n375);
    nor g1667(n375 ,n337 ,n374);
    xor g1668(n1436 ,n373 ,n366);
    nor g1669(n374 ,n367 ,n373);
    nor g1670(n373 ,n327 ,n372);
    xor g1671(n1435 ,n371 ,n356);
    nor g1672(n372 ,n357 ,n371);
    nor g1673(n371 ,n331 ,n370);
    xor g1674(n1434 ,n369 ,n354);
    nor g1675(n370 ,n355 ,n369);
    nor g1676(n369 ,n330 ,n368);
    xnor g1677(n1433 ,n352 ,n328);
    nor g1678(n368 ,n329 ,n353);
    not g1679(n367 ,n366);
    not g1680(n365 ,n364);
    not g1681(n363 ,n362);
    not g1682(n361 ,n360);
    not g1683(n359 ,n358);
    not g1684(n357 ,n356);
    not g1685(n355 ,n354);
    not g1686(n353 ,n352);
    xnor g1687(n366 ,n4[4] ,n7[4]);
    xnor g1688(n364 ,n4[6] ,n7[6]);
    xnor g1689(n362 ,n4[8] ,n7[8]);
    xnor g1690(n360 ,n4[5] ,n7[5]);
    xnor g1691(n358 ,n4[12] ,n7[12]);
    xnor g1692(n356 ,n4[3] ,n7[3]);
    xnor g1693(n354 ,n4[2] ,n7[2]);
    xnor g1694(n352 ,n7[1] ,n4[1]);
    not g1695(n351 ,n350);
    not g1696(n349 ,n348);
    not g1697(n347 ,n346);
    not g1698(n345 ,n344);
    not g1699(n343 ,n342);
    not g1700(n341 ,n340);
    not g1701(n339 ,n338);
    xor g1702(n1432 ,n7[0] ,n4[0]);
    xnor g1703(n350 ,n4[13] ,n7[13]);
    xnor g1704(n348 ,n4[7] ,n7[7]);
    xnor g1705(n346 ,n4[14] ,n7[14]);
    xnor g1706(n344 ,n4[15] ,n7[15]);
    xnor g1707(n342 ,n4[9] ,n7[9]);
    xnor g1708(n340 ,n4[10] ,n7[10]);
    xnor g1709(n338 ,n4[11] ,n7[11]);
    nor g1710(n337 ,n314 ,n4[4]);
    nor g1711(n336 ,n313 ,n4[13]);
    nor g1712(n335 ,n319 ,n4[6]);
    nor g1713(n334 ,n317 ,n4[5]);
    nor g1714(n333 ,n316 ,n4[8]);
    nor g1715(n332 ,n312 ,n4[10]);
    nor g1716(n331 ,n315 ,n4[2]);
    nor g1717(n330 ,n310 ,n4[1]);
    not g1718(n329 ,n328);
    nor g1719(n327 ,n320 ,n4[3]);
    nor g1720(n326 ,n318 ,n4[9]);
    nor g1721(n325 ,n307 ,n4[7]);
    nor g1722(n324 ,n308 ,n4[14]);
    nor g1723(n323 ,n311 ,n4[15]);
    nor g1724(n322 ,n305 ,n4[11]);
    nor g1725(n321 ,n306 ,n4[12]);
    nor g1726(n328 ,n309 ,n4[0]);
    not g1727(n320 ,n7[3]);
    not g1728(n319 ,n7[6]);
    not g1729(n318 ,n7[9]);
    not g1730(n317 ,n7[5]);
    not g1731(n316 ,n7[8]);
    not g1732(n315 ,n7[2]);
    not g1733(n314 ,n7[4]);
    not g1734(n313 ,n7[13]);
    not g1735(n312 ,n7[10]);
    not g1736(n311 ,n7[15]);
    not g1737(n310 ,n7[1]);
    not g1738(n309 ,n7[0]);
    not g1739(n308 ,n7[14]);
    not g1740(n307 ,n7[7]);
    not g1741(n306 ,n7[12]);
    not g1742(n305 ,n7[11]);
    buf g1743(n803 ,n789);
    buf g1744(n805 ,n797);
    buf g1745(n802 ,n792);
    not g1746(n1702 ,n1);
    nor g1747(n1703 ,n1698 ,n1701);
    or g1748(n1701 ,n1690 ,n1700);
    or g1749(n1700 ,n1695 ,n1699);
    or g1750(n1699 ,n1697 ,n1696);
    or g1751(n1698 ,n1692 ,n1694);
    or g1752(n1697 ,n1691 ,n1688);
    or g1753(n1696 ,n1693 ,n1689);
    not g1754(n1695 ,n8[7]);
    not g1755(n1694 ,n8[5]);
    not g1756(n1693 ,n8[1]);
    not g1757(n1692 ,n8[6]);
    not g1758(n1691 ,n8[3]);
    not g1759(n1690 ,n8[4]);
    not g1760(n1689 ,n8[0]);
    not g1761(n1688 ,n8[2]);
    dff g1762(.RN(n1667), .SN(n1683), .CK(n0), .D(n1715), .Q(n7[4]));
    dff g1763(.RN(n1670), .SN(n1685), .CK(n0), .D(n1718), .Q(n7[1]));
    dff g1764(.RN(n1669), .SN(n1687), .CK(n0), .D(n1717), .Q(n7[2]));
    dff g1765(.RN(n1668), .SN(n1684), .CK(n0), .D(n1716), .Q(n7[3]));
    dff g1766(.RN(n1671), .SN(n1686), .CK(n0), .D(n2[0]), .Q(n7[0]));
    dff g1767(.RN(n1666), .SN(n1682), .CK(n0), .D(n1714), .Q(n7[5]));
    dff g1768(.RN(n1664), .SN(n1681), .CK(n0), .D(n1713), .Q(n7[6]));
    dff g1769(.RN(n1665), .SN(n1680), .CK(n0), .D(n1712), .Q(n7[7]));
    dff g1770(.RN(n1656), .SN(n1675), .CK(n0), .D(n1707), .Q(n7[12]));
    dff g1771(.RN(n1661), .SN(n1678), .CK(n0), .D(n1710), .Q(n7[9]));
    dff g1772(.RN(n1660), .SN(n1677), .CK(n0), .D(n1709), .Q(n7[10]));
    dff g1773(.RN(n1659), .SN(n1676), .CK(n0), .D(n1708), .Q(n7[11]));
    dff g1774(.RN(n1662), .SN(n1679), .CK(n0), .D(n1711), .Q(n7[8]));
    dff g1775(.RN(n1658), .SN(n1674), .CK(n0), .D(n1706), .Q(n7[13]));
    dff g1776(.RN(n1657), .SN(n1673), .CK(n0), .D(n1705), .Q(n7[14]));
    dff g1777(.RN(n1663), .SN(n1672), .CK(n0), .D(n1704), .Q(n7[15]));
    or g1778(n1687 ,n1702 ,n1654);
    dff g1779(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1722), .Q(n8[4]));
    dff g1780(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1721), .Q(n8[5]));
    dff g1781(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1725), .Q(n8[1]));
    dff g1782(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1719), .Q(n8[7]));
    dff g1783(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1724), .Q(n8[2]));
    dff g1784(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1720), .Q(n8[6]));
    or g1785(n1686 ,n1702 ,n1639);
    or g1786(n1685 ,n1702 ,n1648);
    dff g1787(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1723), .Q(n8[3]));
    or g1788(n1684 ,n1702 ,n1649);
    or g1789(n1683 ,n1702 ,n1643);
    or g1790(n1682 ,n1702 ,n1651);
    or g1791(n1681 ,n1702 ,n1647);
    or g1792(n1680 ,n1702 ,n1644);
    or g1793(n1679 ,n1702 ,n1650);
    or g1794(n1678 ,n1702 ,n1646);
    or g1795(n1677 ,n1702 ,n1652);
    or g1796(n1676 ,n1702 ,n1640);
    dff g1797(.RN(n1702), .SN(1'b1), .CK(n0), .D(n1653), .Q(n8[0]));
    or g1798(n1675 ,n1702 ,n1642);
    or g1799(n1674 ,n1702 ,n1645);
    or g1800(n1673 ,n1702 ,n1641);
    or g1801(n1672 ,n1702 ,n1655);
    or g1802(n1671 ,n1702 ,n2[0]);
    or g1803(n1670 ,n1702 ,n2[1]);
    or g1804(n1669 ,n1702 ,n2[2]);
    or g1805(n1668 ,n1702 ,n2[3]);
    or g1806(n1667 ,n1702 ,n2[4]);
    or g1807(n1666 ,n1702 ,n2[5]);
    or g1808(n1665 ,n1702 ,n2[7]);
    or g1809(n1664 ,n1702 ,n2[6]);
    or g1810(n1663 ,n1702 ,n2[15]);
    or g1811(n1662 ,n1702 ,n2[8]);
    or g1812(n1661 ,n1702 ,n2[9]);
    or g1813(n1660 ,n1702 ,n2[10]);
    or g1814(n1659 ,n1702 ,n2[11]);
    or g1815(n1658 ,n1702 ,n2[13]);
    or g1816(n1657 ,n1702 ,n2[14]);
    or g1817(n1656 ,n1702 ,n2[12]);
    not g1818(n1655 ,n2[15]);
    not g1819(n1654 ,n2[2]);
    not g1820(n1653 ,n8[0]);
    not g1821(n1652 ,n2[10]);
    not g1822(n1651 ,n2[5]);
    not g1823(n1650 ,n2[8]);
    not g1824(n1649 ,n2[3]);
    not g1825(n1648 ,n2[1]);
    not g1826(n1647 ,n2[6]);
    not g1827(n1646 ,n2[9]);
    not g1828(n1645 ,n2[13]);
    not g1829(n1644 ,n2[7]);
    not g1830(n1643 ,n2[4]);
    not g1831(n1642 ,n2[12]);
    not g1832(n1641 ,n2[14]);
    not g1833(n1640 ,n2[11]);
    not g1834(n1639 ,n2[0]);
    xor g1835(n1704 ,n2[15] ,n1614);
    nor g1836(n1705 ,n1613 ,n1614);
    nor g1837(n1614 ,n1567 ,n1612);
    nor g1838(n1613 ,n2[14] ,n1611);
    nor g1839(n1706 ,n1610 ,n1611);
    not g1840(n1612 ,n1611);
    nor g1841(n1611 ,n1563 ,n1609);
    nor g1842(n1610 ,n2[13] ,n1608);
    nor g1843(n1707 ,n1607 ,n1608);
    not g1844(n1609 ,n1608);
    nor g1845(n1608 ,n1573 ,n1606);
    nor g1846(n1607 ,n2[12] ,n1605);
    nor g1847(n1708 ,n1604 ,n1605);
    not g1848(n1606 ,n1605);
    nor g1849(n1605 ,n1564 ,n1603);
    nor g1850(n1604 ,n2[11] ,n1602);
    nor g1851(n1709 ,n1601 ,n1602);
    not g1852(n1603 ,n1602);
    nor g1853(n1602 ,n1571 ,n1600);
    nor g1854(n1601 ,n2[10] ,n1599);
    nor g1855(n1710 ,n1598 ,n1599);
    not g1856(n1600 ,n1599);
    nor g1857(n1599 ,n1566 ,n1597);
    nor g1858(n1598 ,n2[9] ,n1596);
    nor g1859(n1711 ,n1595 ,n1596);
    not g1860(n1597 ,n1596);
    nor g1861(n1596 ,n1570 ,n1594);
    nor g1862(n1595 ,n2[8] ,n1593);
    nor g1863(n1712 ,n1592 ,n1593);
    not g1864(n1594 ,n1593);
    nor g1865(n1593 ,n1572 ,n1591);
    nor g1866(n1592 ,n2[7] ,n1590);
    nor g1867(n1713 ,n1589 ,n1590);
    not g1868(n1591 ,n1590);
    nor g1869(n1590 ,n1562 ,n1588);
    nor g1870(n1589 ,n2[6] ,n1587);
    nor g1871(n1714 ,n1586 ,n1587);
    not g1872(n1588 ,n1587);
    nor g1873(n1587 ,n1565 ,n1585);
    nor g1874(n1586 ,n2[5] ,n1584);
    nor g1875(n1715 ,n1583 ,n1584);
    not g1876(n1585 ,n1584);
    nor g1877(n1584 ,n1561 ,n1582);
    nor g1878(n1583 ,n2[4] ,n1581);
    xor g1879(n1716 ,n2[3] ,n1579);
    not g1880(n1582 ,n1581);
    nor g1881(n1581 ,n1568 ,n1580);
    nor g1882(n1717 ,n1578 ,n1579);
    not g1883(n1580 ,n1579);
    nor g1884(n1579 ,n1560 ,n1577);
    nor g1885(n1578 ,n2[2] ,n1576);
    nor g1886(n1718 ,n1576 ,n1575);
    not g1887(n1577 ,n1576);
    nor g1888(n1576 ,n1574 ,n1569);
    nor g1889(n1575 ,n2[1] ,n1703);
    not g1890(n1574 ,n2[1]);
    not g1891(n1573 ,n2[12]);
    not g1892(n1572 ,n2[7]);
    not g1893(n1571 ,n2[10]);
    not g1894(n1570 ,n2[8]);
    not g1895(n1569 ,n1703);
    not g1896(n1568 ,n2[3]);
    not g1897(n1567 ,n2[14]);
    not g1898(n1566 ,n2[9]);
    not g1899(n1565 ,n2[5]);
    not g1900(n1564 ,n2[11]);
    not g1901(n1563 ,n2[13]);
    not g1902(n1562 ,n2[6]);
    not g1903(n1561 ,n2[4]);
    not g1904(n1560 ,n2[2]);
    xor g1905(n1719 ,n8[7] ,n1638);
    nor g1906(n1720 ,n1637 ,n1638);
    nor g1907(n1638 ,n1615 ,n1636);
    nor g1908(n1637 ,n8[6] ,n1635);
    nor g1909(n1721 ,n1634 ,n1635);
    not g1910(n1636 ,n1635);
    nor g1911(n1635 ,n1620 ,n1633);
    nor g1912(n1634 ,n8[5] ,n1632);
    nor g1913(n1722 ,n1631 ,n1632);
    not g1914(n1633 ,n1632);
    nor g1915(n1632 ,n1617 ,n1630);
    nor g1916(n1631 ,n8[4] ,n1629);
    nor g1917(n1723 ,n1628 ,n1629);
    not g1918(n1630 ,n1629);
    nor g1919(n1629 ,n1618 ,n1627);
    nor g1920(n1628 ,n8[3] ,n1626);
    nor g1921(n1724 ,n1625 ,n1626);
    not g1922(n1627 ,n1626);
    nor g1923(n1626 ,n1621 ,n1624);
    nor g1924(n1625 ,n8[2] ,n1623);
    nor g1925(n1725 ,n1623 ,n1622);
    not g1926(n1624 ,n1623);
    nor g1927(n1623 ,n1619 ,n1616);
    nor g1928(n1622 ,n8[1] ,n8[0]);
    not g1929(n1621 ,n8[2]);
    not g1930(n1620 ,n8[5]);
    not g1931(n1619 ,n8[1]);
    not g1932(n1618 ,n8[3]);
    not g1933(n1617 ,n8[4]);
    not g1934(n1616 ,n8[0]);
    not g1935(n1615 ,n8[6]);
endmodule
