module top (n0, n1, n2, n3, n4, n5, n6, n8, n9, n7, n10);
    input n0, n1, n2;
    input [13:0] n3;
    input [12:0] n4;
    input [7:0] n5, n6, n7;
    input [5:0] n8;
    input [9:0] n9;
    output [12:0] n10;
    wire n0, n1, n2;
    wire [13:0] n3;
    wire [12:0] n4;
    wire [7:0] n5, n6, n7;
    wire [5:0] n8;
    wire [9:0] n9;
    wire [12:0] n10;
    wire [13:0] n11;
    wire [9:0] n12;
    wire [12:0] n13;
    wire [13:0] n14;
    wire [7:0] n15;
    wire [7:0] n16;
    wire [12:0] n17;
    wire [5:0] n18;
    wire [7:0] n19;
    wire [7:0] n20;
    wire [7:0] n21;
    wire [7:0] n22;
    wire [7:0] n23;
    wire [7:0] n24;
    wire [12:0] n25;
    wire n26, n27, n28, n29, n30, n31, n32, n33;
    wire n34, n35, n36, n37, n38, n39, n40, n41;
    wire n42, n43, n44, n45, n46, n47, n48, n49;
    wire n50, n51, n52, n53, n54, n55, n56, n57;
    wire n58, n59, n60, n61, n62, n63, n64, n65;
    wire n66, n67, n68, n69, n70, n71, n72, n73;
    wire n74, n75, n76, n77, n78, n79, n80, n81;
    wire n82, n83, n84, n85, n86, n87, n88, n89;
    wire n90, n91, n92, n93, n94, n95, n96, n97;
    wire n98, n99, n100, n101, n102, n103, n104, n105;
    wire n106, n107, n108, n109, n110, n111, n112, n113;
    wire n114, n115, n116, n117, n118, n119, n120, n121;
    wire n122, n123, n124, n125, n126, n127, n128, n129;
    wire n130, n131, n132, n133, n134, n135, n136, n137;
    wire n138, n139, n140, n141, n142, n143, n144, n145;
    wire n146, n147, n148, n149, n150, n151, n152, n153;
    wire n154, n155, n156, n157, n158, n159, n160, n161;
    wire n162, n163, n164, n165, n166, n167, n168, n169;
    wire n170, n171, n172, n173, n174, n175, n176, n177;
    wire n178, n179, n180, n181, n182, n183, n184, n185;
    wire n186, n187, n188, n189, n190, n191, n192, n193;
    wire n194, n195, n196, n197, n198, n199, n200, n201;
    wire n202, n203, n204, n205, n206, n207, n208, n209;
    wire n210, n211, n212, n213, n214, n215, n216, n217;
    wire n218, n219, n220, n221, n222, n223, n224, n225;
    wire n226, n227, n228, n229, n230, n231, n232, n233;
    wire n234, n235, n236, n237, n238, n239, n240, n241;
    wire n242, n243, n244, n245, n246, n247, n248, n249;
    wire n250, n251, n252, n253, n254, n255, n256, n257;
    wire n258, n259, n260, n261, n262, n263, n264, n265;
    wire n266, n267, n268, n269, n270, n271, n272, n273;
    wire n274, n275, n276, n277, n278, n279, n280, n281;
    wire n282, n283, n284, n285, n286, n287, n288, n289;
    wire n290, n291, n292, n293, n294, n295, n296, n297;
    wire n298, n299, n300, n301, n302, n303, n304, n305;
    wire n306, n307, n308, n309, n310;
    dff g0(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[2]), .Q(n10[2]));
    not g1(n29 ,n12[2]);
    nor g2(n86 ,n11[10] ,n53);
    not g3(n269 ,n13[2]);
    nor g4(n165 ,n16[4] ,n137);
    xor g5(n13[2] ,n15[2] ,n239);
    or g6(n225 ,n185 ,n208);
    nor g7(n25[7] ,n288 ,n289);
    not g8(n259 ,n13[7]);
    not g9(n241 ,n240);
    not g10(n255 ,n12[8]);
    not g11(n63 ,n64);
    nor g12(n273 ,n13[2] ,n271);
    not g13(n254 ,n11[3]);
    buf g14(n10[9], 1'b0);
    nor g15(n279 ,n13[4] ,n277);
    xnor g16(n75 ,n20[0] ,n21[0]);
    dff g17(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[11]), .Q(n11[11]));
    nor g18(n229 ,n165 ,n219);
    not g19(n32 ,n12[4]);
    xnor g20(n100 ,n63 ,n11[6]);
    not g21(n135 ,n134);
    nor g22(n288 ,n13[7] ,n286);
    nor g23(n230 ,n188 ,n199);
    nor g24(n25[6] ,n285 ,n286);
    xnor g25(n70 ,n16[2] ,n29);
    not g26(n60 ,n59);
    nor g27(n276 ,n13[3] ,n274);
    not g28(n258 ,n13[1]);
    not g29(n272 ,n271);
    not g30(n33 ,n12[3]);
    xnor g31(n99 ,n66 ,n11[7]);
    nor g32(n85 ,n11[11] ,n59);
    xnor g33(n104 ,n66 ,n17[6]);
    or g34(n222 ,n213 ,n207);
    nor g35(n179 ,n102 ,n145);
    nor g36(n202 ,n134 ,n177);
    nor g37(n305 ,n14[13] ,n14[12]);
    dff g38(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[2]), .Q(n17[2]));
    xnor g39(n73 ,n19[2] ,n16[2]);
    xor g40(n13[1] ,n15[1] ,n238);
    nor g41(n80 ,n42 ,n64);
    buf g42(n10[11], 1'b0);
    not g43(n194 ,n193);
    nor g44(n220 ,n174 ,n217);
    xor g45(n124 ,n90 ,n58);
    or g46(n148 ,n36 ,n112);
    nor g47(n242 ,n196 ,n236);
    buf g48(n10[7], 1'b0);
    nor g49(n221 ,n167 ,n219);
    nor g50(n154 ,n56 ,n125);
    xnor g51(n52 ,n17[1] ,n17[11]);
    not g52(n128 ,n127);
    xnor g53(n78 ,n16[3] ,n18[3]);
    dff g54(.RN(n1), .SN(1'b1), .CK(n0), .D(n7[2]), .Q(n15[2]));
    nor g55(n297 ,n13[10] ,n295);
    xnor g56(n62 ,n20[0] ,n22[0]);
    nor g57(n177 ,n104 ,n149);
    not g58(n54 ,n53);
    nor g59(n118 ,n86 ,n109);
    or g60(n119 ,n61 ,n107);
    nor g61(n196 ,n132 ,n191);
    nor g62(n89 ,n40 ,n65);
    nor g63(n94 ,n256 ,n69);
    nor g64(n208 ,n12[7] ,n189);
    nor g65(n144 ,n55 ,n122);
    nor g66(n134 ,n77 ,n111);
    or g67(n14[12] ,n252 ,n251);
    not g68(n188 ,n187);
    or g69(n151 ,n47 ,n115);
    nor g70(n249 ,n203 ,n227);
    nor g71(n248 ,n168 ,n233);
    not g72(n299 ,n298);
    not g73(n123 ,n122);
    dff g74(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[7]), .Q(n12[7]));
    dff g75(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[12]), .Q(n10[12]));
    nor g76(n271 ,n258 ,n266);
    nor g77(n174 ,n39 ,n141);
    or g78(n234 ,n43 ,n215);
    not g79(n293 ,n292);
    nor g80(n240 ,n190 ,n197);
    xnor g81(n57 ,n18[4] ,n22[0]);
    or g82(n14[13] ,n253 ,n250);
    not g83(n130 ,n129);
    not g84(n41 ,n12[5]);
    buf g85(n10[10], 1'b0);
    not g86(n182 ,n181);
    or g87(n125 ,n87 ,n108);
    not g88(n45 ,n12[6]);
    nor g89(n167 ,n16[4] ,n140);
    not g90(n303 ,n14[12]);
    nor g91(n84 ,n44 ,n64);
    not g92(n156 ,n155);
    buf g93(n10[4], 1'b0);
    dff g94(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[1]), .Q(n10[1]));
    not g95(n268 ,n13[3]);
    nor g96(n169 ,n52 ,n152);
    buf g97(n10[12], 1'b0);
    not g98(n264 ,n13[6]);
    xnor g99(n58 ,n19[4] ,n21[0]);
    nor g100(n107 ,n73 ,n95);
    nor g101(n270 ,n13[1] ,n310);
    nor g102(n239 ,n29 ,n205);
    xnor g103(n101 ,n68 ,n17[8]);
    nor g104(n286 ,n264 ,n284);
    not g105(n184 ,n183);
    not g106(n28 ,n12[0]);
    nor g107(n90 ,n36 ,n54);
    or g108(n226 ,n193 ,n216);
    nor g109(n251 ,n226 ,n230);
    nor g110(n294 ,n13[9] ,n292);
    not g111(n27 ,n16[4]);
    not g112(n284 ,n283);
    dff g113(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[2]), .Q(n18[2]));
    nor g114(n283 ,n262 ,n281);
    or g115(n236 ,n255 ,n211);
    nor g116(n277 ,n268 ,n275);
    dff g117(.RN(n1), .SN(1'b1), .CK(n0), .D(n26), .Q(n10[0]));
    not g118(n275 ,n274);
    nor g119(n160 ,n154 ,n155);
    dff g120(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[4]), .Q(n10[4]));
    or g121(n110 ,n46 ,n93);
    or g122(n149 ,n40 ,n114);
    nor g123(n159 ,n70 ,n138);
    nor g124(n175 ,n69 ,n130);
    dff g125(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[11]), .Q(n10[11]));
    nor g126(n191 ,n101 ,n146);
    not g127(n140 ,n139);
    dff g128(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[4]), .Q(n11[4]));
    nor g129(n247 ,n202 ,n235);
    nor g130(n126 ,n56 ,n123);
    dff g131(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[8]), .Q(n12[8]));
    xor g132(n112 ,n82 ,n71);
    nor g133(n141 ,n56 ,n116);
    or g134(n145 ,n48 ,n111);
    not g135(n192 ,n191);
    nor g136(n93 ,n34 ,n60);
    nor g137(n244 ,n200 ,n222);
    not g138(n37 ,n11[10]);
    xnor g139(n102 ,n70 ,n17[7]);
    nor g140(n25[1] ,n271 ,n270);
    xnor g141(n64 ,n20[0] ,n12[0]);
    dff g142(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[5]), .Q(n12[5]));
    dff g143(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[0]), .Q(n22[0]));
    nor g144(n25[5] ,n282 ,n283);
    nor g145(n250 ,n225 ,n240);
    nor g146(n198 ,n169 ,n177);
    xnor g147(n51 ,n17[0] ,n17[10]);
    not g148(n190 ,n189);
    nor g149(n253 ,n186 ,n241);
    dff g150(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[3]), .Q(n18[3]));
    xor g151(n25[12] ,n13[12] ,n301);
    xor g152(n13[6] ,n247 ,n238);
    dff g153(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[6]), .Q(n10[6]));
    xor g154(n113 ,n79 ,n58);
    xor g155(n121 ,n81 ,n73);
    nor g156(n200 ,n136 ,n183);
    not g157(n69 ,n70);
    nor g158(n187 ,n100 ,n150);
    not g159(n309 ,n2);
    xnor g160(n66 ,n16[1] ,n30);
    dff g161(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[1]), .Q(n17[1]));
    dff g162(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[6]), .Q(n11[6]));
    buf g163(n10[2], 1'b0);
    or g164(n235 ,n45 ,n218);
    not g165(n42 ,n17[0]);
    or g166(n205 ,n159 ,n175);
    nor g167(n158 ,n63 ,n131);
    xor g168(n115 ,n88 ,n76);
    nor g169(n171 ,n66 ,n127);
    or g170(n146 ,n49 ,n121);
    dff g171(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[1]), .Q(n16[1]));
    nor g172(n301 ,n267 ,n299);
    nor g173(n228 ,n160 ,n212);
    dff g174(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[5]), .Q(n18[5]));
    nor g175(n214 ,n153 ,n182);
    not g176(n265 ,n13[8]);
    dff g177(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[4]), .Q(n18[4]));
    dff g178(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[1]), .Q(n19[1]));
    dff g179(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[3]), .Q(n17[3]));
    not g180(n142 ,n141);
    xor g181(n13[11] ,n245 ,n247);
    or g182(n108 ,n42 ,n84);
    dff g183(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[3]), .Q(n16[3]));
    dff g184(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[10]), .Q(n17[10]));
    or g185(n223 ,n210 ,n205);
    nor g186(n210 ,n170 ,n178);
    not g187(n30 ,n12[1]);
    xor g188(n116 ,n50 ,n91);
    nor g189(n298 ,n260 ,n296);
    not g190(n231 ,n230);
    nor g191(n274 ,n269 ,n272);
    nor g192(n138 ,n98 ,n119);
    dff g193(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[0]), .Q(n20[0]));
    nor g194(n96 ,n254 ,n67);
    dff g195(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[8]), .Q(n17[8]));
    nor g196(n127 ,n77 ,n115);
    buf g197(n10[0], 1'b0);
    nor g198(n282 ,n13[5] ,n280);
    nor g199(n307 ,n306 ,n304);
    dff g200(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[10]), .Q(n10[10]));
    not g201(n290 ,n289);
    nor g202(n237 ,n33 ,n206);
    nor g203(n216 ,n12[6] ,n187);
    xnor g204(n26 ,n257 ,n24[0]);
    not g205(n47 ,n11[1]);
    dff g206(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[5]), .Q(n11[5]));
    dff g207(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[2]), .Q(n19[2]));
    nor g208(n172 ,n153 ,n156);
    dff g209(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[0]), .Q(n17[0]));
    nor g210(n136 ,n57 ,n124);
    not g211(n267 ,n13[11]);
    nor g212(n91 ,n46 ,n60);
    nor g213(n105 ,n71 ,n97);
    dff g214(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[3]), .Q(n19[3]));
    nor g215(n79 ,n38 ,n54);
    dff g216(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[3]), .Q(n12[3]));
    dff g217(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[5]), .Q(n10[5]));
    nor g218(n218 ,n135 ,n178);
    not g219(n180 ,n179);
    not g220(n281 ,n280);
    dff g221(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[0]), .Q(n21[0]));
    not g222(n97 ,n96);
    xnor g223(n13[5] ,n257 ,n228);
    xor g224(n13[10] ,n249 ,n228);
    dff g225(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[5]), .Q(n19[5]));
    nor g226(n193 ,n45 ,n131);
    nor g227(n25[4] ,n279 ,n280);
    nor g228(n166 ,n65 ,n135);
    dff g229(.RN(n1), .SN(1'b1), .CK(n0), .D(n8[1]), .Q(n18[1]));
    or g230(n224 ,n171 ,n209);
    nor g231(n161 ,n65 ,n128);
    or g232(n120 ,n78 ,n105);
    dff g233(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[7]), .Q(n11[7]));
    not g234(n39 ,n16[5]);
    dff g235(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[5]), .Q(n16[5]));
    not g236(n266 ,n310);
    nor g237(n82 ,n49 ,n67);
    dff g238(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[2]), .Q(n11[2]));
    dff g239(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[3]), .Q(n10[3]));
    dff g240(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[8]), .Q(n10[8]));
    not g241(n74 ,n73);
    xor g242(n13[3] ,n15[3] ,n237);
    dff g243(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[6]), .Q(n17[6]));
    not g244(n35 ,n23[0]);
    xnor g245(n197 ,n67 ,n143);
    not g246(n95 ,n94);
    nor g247(n291 ,n13[8] ,n289);
    not g248(n133 ,n132);
    dff g249(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[0]), .Q(n12[0]));
    nor g250(n183 ,n103 ,n148);
    xor g251(n14[10] ,n248 ,n221);
    nor g252(n83 ,n35 ,n64);
    dff g253(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[7]), .Q(n17[7]));
    xnor g254(n50 ,n19[5] ,n19[1]);
    or g255(n209 ,n144 ,n162);
    nor g256(n139 ,n57 ,n113);
    not g257(n72 ,n71);
    not g258(n46 ,n11[5]);
    nor g259(n238 ,n30 ,n204);
    nor g260(n25[3] ,n276 ,n277);
    or g261(n257 ,n28 ,n207);
    nor g262(n289 ,n259 ,n287);
    not g263(n43 ,n12[7]);
    or g264(n206 ,n157 ,n164);
    nor g265(n164 ,n67 ,n133);
    buf g266(n10[3], 1'b0);
    xor g267(n114 ,n80 ,n75);
    xnor g268(n76 ,n16[1] ,n19[1]);
    dff g269(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[6]), .Q(n12[6]));
    xnor g270(n71 ,n19[3] ,n16[3]);
    not g271(n170 ,n169);
    or g272(n162 ,n126 ,n116);
    dff g273(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[4]), .Q(n16[4]));
    nor g274(n155 ,n62 ,n114);
    nor g275(n157 ,n68 ,n143);
    dff g276(.RN(n1), .SN(1'b1), .CK(n0), .D(n7[4]), .Q(n15[4]));
    xor g277(n168 ,n118 ,n57);
    dff g278(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[0]), .Q(n23[0]));
    xnor g279(n201 ,n63 ,n131);
    nor g280(n132 ,n78 ,n112);
    dff g281(.RN(n1), .SN(1'b1), .CK(n0), .D(n6[4]), .Q(n19[4]));
    not g282(n262 ,n13[5]);
    xnor g283(n61 ,n16[2] ,n18[2]);
    nor g284(n92 ,n37 ,n54);
    not g285(n49 ,n17[3]);
    xnor g286(n53 ,n27 ,n12[4]);
    nor g287(n185 ,n43 ,n127);
    not g288(n287 ,n286);
    dff g289(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[9]), .Q(n10[9]));
    nor g290(n106 ,n72 ,n96);
    nor g291(n243 ,n161 ,n224);
    nor g292(n88 ,n47 ,n65);
    nor g293(n310 ,n309 ,n308);
    or g294(n150 ,n35 ,n117);
    nor g295(n143 ,n106 ,n120);
    nor g296(n292 ,n265 ,n290);
    nor g297(n300 ,n13[11] ,n298);
    nor g298(n129 ,n61 ,n121);
    xor g299(n13[4] ,n15[4] ,n229);
    not g300(n178 ,n177);
    buf g301(n10[6], 1'b0);
    xor g302(n13[9] ,n244 ,n229);
    dff g303(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[2]), .Q(n12[2]));
    dff g304(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[10]), .Q(n11[10]));
    dff g305(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[4]), .Q(n12[4]));
    dff g306(.RN(n1), .SN(1'b1), .CK(n0), .D(n7[0]), .Q(n24[0]));
    or g307(n147 ,n44 ,n124);
    nor g308(n25[8] ,n291 ,n292);
    or g309(n109 ,n38 ,n92);
    xor g310(n111 ,n89 ,n76);
    nor g311(n211 ,n133 ,n192);
    nor g312(n280 ,n263 ,n278);
    not g313(n256 ,n11[2]);
    nor g314(n25[9] ,n294 ,n295);
    or g315(n306 ,n302 ,n303);
    or g316(n212 ,n41 ,n172);
    nor g317(n81 ,n48 ,n69);
    nor g318(n25[11] ,n300 ,n301);
    not g319(n153 ,n154);
    not g320(n40 ,n17[1]);
    not g321(n36 ,n17[4]);
    not g322(n65 ,n66);
    xnor g323(n103 ,n53 ,n17[9]);
    or g324(n227 ,n214 ,n204);
    not g325(n296 ,n295);
    buf g326(n10[8], 1'b0);
    nor g327(n203 ,n154 ,n181);
    dff g328(.RN(n1), .SN(1'b1), .CK(n0), .D(n7[3]), .Q(n15[3]));
    dff g329(.RN(n1), .SN(1'b1), .CK(n0), .D(n5[2]), .Q(n16[2]));
    dff g330(.RN(n1), .SN(1'b1), .CK(n0), .D(n9[1]), .Q(n12[1]));
    nor g331(n98 ,n74 ,n94);
    dff g332(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[5]), .Q(n17[5]));
    not g333(n186 ,n185);
    not g334(n137 ,n136);
    buf g335(n10[5], 1'b0);
    not g336(n48 ,n17[2]);
    not g337(n260 ,n13[10]);
    nor g338(n295 ,n261 ,n293);
    nor g339(n245 ,n198 ,n223);
    not g340(n263 ,n13[4]);
    xnor g341(n77 ,n16[1] ,n18[1]);
    nor g342(n215 ,n130 ,n180);
    not g343(n302 ,n14[13]);
    nor g344(n176 ,n16[5] ,n142);
    nor g345(n213 ,n137 ,n184);
    xnor g346(n68 ,n16[3] ,n33);
    dff g347(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[3]), .Q(n11[3]));
    not g348(n44 ,n17[5]);
    xnor g349(n59 ,n16[5] ,n41);
    or g350(n204 ,n171 ,n166);
    xor g351(n13[7] ,n246 ,n239);
    nor g352(n195 ,n129 ,n179);
    nor g353(n246 ,n195 ,n234);
    xnor g354(n199 ,n69 ,n138);
    xor g355(n14[11] ,n243 ,n220);
    nor g356(n304 ,n14[11] ,n14[10]);
    or g357(n217 ,n41 ,n176);
    dff g358(.RN(n1), .SN(1'b1), .CK(n0), .D(n3[1]), .Q(n11[1]));
    nor g359(n163 ,n64 ,n156);
    nor g360(n232 ,n180 ,n206);
    dff g361(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[9]), .Q(n17[9]));
    not g362(n67 ,n68);
    nor g363(n131 ,n62 ,n117);
    nor g364(n285 ,n13[6] ,n283);
    or g365(n308 ,n305 ,n307);
    nor g366(n25[10] ,n297 ,n298);
    not g367(n278 ,n277);
    not g368(n34 ,n11[11]);
    nor g369(n252 ,n194 ,n231);
    nor g370(n122 ,n85 ,n110);
    dff g371(.RN(n1), .SN(1'b1), .CK(n0), .D(n7[1]), .Q(n15[1]));
    not g372(n261 ,n13[9]);
    nor g373(n181 ,n51 ,n147);
    nor g374(n189 ,n99 ,n151);
    dff g375(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[11]), .Q(n17[11]));
    xnor g376(n56 ,n18[5] ,n18[1]);
    nor g377(n87 ,n17[5] ,n63);
    not g378(n31 ,n17[6]);
    xor g379(n13[8] ,n242 ,n237);
    dff g380(.RN(n1), .SN(1'b1), .CK(n0), .D(n4[4]), .Q(n17[4]));
    not g381(n38 ,n11[4]);
    or g382(n152 ,n31 ,n125);
    nor g383(n173 ,n27 ,n139);
    or g384(n207 ,n158 ,n163);
    xor g385(n117 ,n83 ,n75);
    dff g386(.RN(n1), .SN(1'b1), .CK(n0), .D(n25[7]), .Q(n10[7]));
    buf g387(n10[1], 1'b0);
    xor g388(n13[12] ,n232 ,n246);
    or g389(n233 ,n113 ,n201);
    nor g390(n25[2] ,n273 ,n274);
    or g391(n219 ,n32 ,n173);
    not g392(n55 ,n56);
endmodule
