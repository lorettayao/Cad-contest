module top(n0, n1, n2, n3, n4, n5, n13, n17, n18, n6, n7, n14, n19, n20, n8, n9, n15, n21, n22, n10, n11, n16, n23, n24, n12, n25, n26, n27, n28, n29, n30, n31, n32, n34, n33);
    input n0, n1;
    input [3:0] n2, n3;
    input [31:0] n4, n5, n6, n7, n8, n9, n10, n11, n12;
    input [15:0] n13, n14, n15, n16;
    input [1:0] n17, n18, n19, n20, n21, n22, n23, n24;
    output [31:0] n25, n26;
    output n27, n28;
    output [3:0] n29, n30;
    output [7:0] n31, n32, n33;
    output [15:0] n34;
    wire n0, n1;
    wire [3:0] n2, n3;
    wire [31:0] n4, n5, n6, n7, n8, n9, n10, n11, n12;
    wire [15:0] n13, n14, n15, n16;
    wire [1:0] n17, n18, n19, n20, n21, n22, n23, n24;
    wire [31:0] n25, n26;
    wire n27, n28;
    wire [3:0] n29, n30;
    wire [7:0] n31, n32, n33;
    wire [15:0] n34;
    wire [3:0] n35;
    wire [3:0] n36;
    wire [3:0] n37;
    wire [3:0] n38;
    wire [3:0] n39;
    wire [31:0] n40;
    wire [15:0] n41;
    wire [31:0] n42;
    wire [2:0] n43;
    wire [1:0] n44;
    wire [2:0] n45;
    wire [31:0] n46;
    wire [31:0] n47;
    wire [31:0] n48;
    wire [31:0] n49;
    wire [15:0] n50;
    wire [15:0] n51;
    wire [15:0] n52;
    wire [15:0] n53;
    wire n54, n55, n56, n57, n58, n59, n60, n61;
    wire n62, n63, n64, n65, n66, n67, n68, n69;
    wire n70, n71, n72, n73, n74, n75, n76, n77;
    wire n78, n79, n80, n81, n82, n83, n84, n85;
    wire n86, n87, n88, n89, n90, n91, n92, n93;
    wire n94, n95, n96, n97, n98, n99, n100, n101;
    wire n102, n103, n104, n105, n106, n107, n108, n109;
    wire n110, n111, n112, n113, n114, n115, n116, n117;
    wire n118, n119, n120, n121, n122, n123, n124, n125;
    wire n126, n127, n128, n129, n130, n131, n132, n133;
    wire n134, n135, n136, n137, n138, n139, n140, n141;
    wire n142, n143, n144, n145, n146, n147, n148, n149;
    wire n150, n151, n152, n153, n154, n155, n156, n157;
    wire n158, n159, n160, n161, n162, n163, n164, n165;
    wire n166, n167, n168, n169, n170, n171, n172, n173;
    wire n174, n175, n176, n177, n178, n179, n180, n181;
    wire n182, n183, n184, n185, n186, n187, n188, n189;
    wire n190, n191, n192, n193, n194, n195, n196, n197;
    wire n198, n199, n200, n201, n202, n203, n204, n205;
    wire n206, n207, n208, n209, n210, n211, n212, n213;
    wire n214, n215, n216, n217, n218, n219, n220, n221;
    wire n222, n223, n224, n225, n226, n227, n228, n229;
    wire n230, n231, n232, n233, n234, n235, n236, n237;
    wire n238, n239, n240, n241, n242, n243, n244, n245;
    wire n246, n247, n248, n249, n250, n251, n252, n253;
    wire n254, n255, n256, n257, n258, n259, n260, n261;
    wire n262, n263, n264, n265, n266, n267, n268, n269;
    wire n270, n271, n272, n273, n274, n275, n276, n277;
    wire n278, n279, n280, n281, n282, n283, n284, n285;
    wire n286, n287, n288, n289, n290, n291, n292, n293;
    wire n294, n295, n296, n297, n298, n299, n300, n301;
    wire n302, n303, n304, n305, n306, n307, n308, n309;
    wire n310, n311, n312, n313, n314, n315, n316, n317;
    wire n318, n319, n320, n321, n322, n323, n324, n325;
    wire n326, n327, n328, n329, n330, n331, n332, n333;
    wire n334, n335, n336, n337, n338, n339, n340, n341;
    wire n342, n343, n344, n345, n346, n347, n348, n349;
    wire n350, n351, n352, n353, n354, n355, n356, n357;
    wire n358, n359, n360, n361, n362, n363, n364, n365;
    wire n366, n367, n368, n369, n370, n371, n372, n373;
    wire n374, n375, n376, n377, n378, n379, n380, n381;
    wire n382, n383, n384, n385, n386, n387, n388, n389;
    wire n390, n391, n392, n393, n394, n395, n396, n397;
    wire n398, n399, n400, n401, n402, n403, n404, n405;
    wire n406, n407, n408, n409, n410, n411, n412, n413;
    wire n414, n415, n416, n417, n418, n419, n420, n421;
    wire n422, n423, n424, n425, n426, n427, n428, n429;
    wire n430, n431, n432, n433, n434, n435, n436, n437;
    wire n438, n439, n440, n441, n442, n443, n444, n445;
    wire n446, n447, n448, n449, n450, n451, n452, n453;
    wire n454, n455, n456, n457, n458, n459, n460, n461;
    wire n462, n463, n464, n465, n466, n467, n468, n469;
    wire n470, n471, n472, n473, n474, n475, n476, n477;
    wire n478, n479, n480, n481, n482, n483, n484, n485;
    wire n486, n487, n488, n489, n490, n491, n492, n493;
    wire n494, n495, n496, n497, n498, n499, n500, n501;
    wire n502, n503, n504, n505, n506, n507, n508, n509;
    wire n510, n511, n512, n513, n514, n515, n516, n517;
    wire n518, n519, n520, n521, n522, n523, n524, n525;
    wire n526, n527, n528, n529, n530, n531, n532, n533;
    wire n534, n535, n536, n537, n538, n539, n540, n541;
    wire n542, n543, n544, n545, n546, n547, n548, n549;
    wire n550, n551, n552, n553, n554, n555, n556, n557;
    wire n558, n559, n560, n561, n562, n563, n564, n565;
    wire n566, n567, n568, n569, n570, n571, n572, n573;
    wire n574, n575, n576, n577, n578, n579, n580, n581;
    wire n582, n583, n584, n585, n586, n587, n588, n589;
    wire n590, n591, n592, n593, n594, n595, n596, n597;
    wire n598, n599, n600, n601, n602, n603, n604, n605;
    wire n606, n607, n608, n609, n610, n611, n612, n613;
    wire n614, n615, n616, n617, n618, n619, n620, n621;
    wire n622, n623, n624, n625, n626, n627, n628, n629;
    wire n630, n631, n632, n633, n634, n635, n636, n637;
    wire n638, n639, n640, n641, n642, n643, n644, n645;
    wire n646, n647, n648, n649, n650, n651, n652, n653;
    wire n654, n655, n656, n657, n658, n659, n660, n661;
    wire n662, n663, n664, n665, n666, n667, n668, n669;
    wire n670, n671, n672, n673, n674, n675, n676, n677;
    wire n678, n679, n680, n681, n682, n683, n684, n685;
    wire n686, n687, n688, n689, n690, n691, n692, n693;
    wire n694, n695, n696, n697, n698, n699, n700, n701;
    wire n702, n703, n704, n705, n706, n707, n708, n709;
    wire n710, n711, n712, n713, n714, n715, n716, n717;
    wire n718, n719, n720, n721, n722, n723, n724, n725;
    wire n726, n727, n728, n729, n730, n731, n732, n733;
    wire n734, n735, n736, n737, n738, n739, n740, n741;
    wire n742, n743, n744, n745, n746, n747, n748, n749;
    wire n750, n751, n752, n753, n754, n755, n756, n757;
    wire n758, n759, n760, n761, n762, n763, n764, n765;
    wire n766, n767, n768, n769, n770, n771, n772, n773;
    wire n774, n775, n776, n777, n778, n779, n780, n781;
    wire n782, n783, n784, n785, n786, n787, n788, n789;
    wire n790, n791, n792, n793, n794, n795, n796, n797;
    wire n798, n799, n800, n801, n802, n803, n804, n805;
    wire n806, n807, n808, n809, n810, n811, n812, n813;
    wire n814, n815, n816, n817, n818, n819, n820, n821;
    wire n822, n823, n824, n825, n826, n827, n828, n829;
    wire n830, n831, n832, n833, n834, n835, n836, n837;
    wire n838, n839, n840, n841, n842, n843, n844, n845;
    wire n846, n847, n848, n849, n850, n851, n852, n853;
    wire n854, n855, n856, n857, n858, n859, n860, n861;
    wire n862, n863, n864, n865, n866, n867, n868, n869;
    wire n870, n871, n872, n873, n874, n875, n876, n877;
    wire n878, n879, n880, n881, n882, n883, n884, n885;
    wire n886, n887, n888, n889, n890, n891, n892, n893;
    wire n894, n895, n896, n897, n898, n899, n900, n901;
    wire n902, n903, n904, n905, n906, n907, n908, n909;
    wire n910, n911, n912, n913, n914, n915, n916, n917;
    wire n918, n919, n920, n921, n922, n923, n924, n925;
    wire n926, n927, n928, n929, n930, n931, n932, n933;
    wire n934, n935, n936, n937, n938, n939, n940, n941;
    wire n942, n943, n944, n945, n946, n947, n948, n949;
    wire n950, n951, n952, n953, n954, n955, n956, n957;
    wire n958, n959, n960, n961, n962, n963, n964, n965;
    wire n966, n967, n968, n969, n970, n971, n972, n973;
    wire n974, n975, n976, n977, n978, n979, n980, n981;
    wire n982, n983, n984, n985, n986, n987, n988, n989;
    wire n990, n991, n992, n993, n994, n995, n996, n997;
    wire n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
    wire n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013;
    wire n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
    wire n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
    wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
    wire n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;
    wire n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053;
    wire n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061;
    wire n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069;
    wire n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077;
    wire n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085;
    wire n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093;
    wire n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
    wire n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109;
    wire n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117;
    wire n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125;
    wire n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133;
    wire n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141;
    wire n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149;
    wire n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157;
    wire n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165;
    wire n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173;
    wire n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181;
    wire n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189;
    wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
    wire n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205;
    wire n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213;
    wire n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221;
    wire n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229;
    wire n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237;
    wire n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245;
    wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
    wire n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261;
    wire n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269;
    wire n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277;
    wire n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285;
    wire n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293;
    wire n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301;
    wire n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309;
    wire n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
    wire n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325;
    wire n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333;
    wire n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341;
    wire n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349;
    wire n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357;
    wire n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365;
    wire n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373;
    wire n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381;
    wire n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389;
    wire n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397;
    wire n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405;
    wire n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413;
    wire n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421;
    wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
    wire n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
    wire n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445;
    wire n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453;
    wire n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;
    wire n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469;
    wire n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477;
    wire n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485;
    wire n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493;
    wire n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501;
    wire n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509;
    wire n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517;
    wire n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525;
    wire n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533;
    wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
    wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
    wire n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
    wire n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565;
    wire n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573;
    wire n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581;
    wire n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589;
    wire n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597;
    wire n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605;
    wire n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613;
    wire n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621;
    wire n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629;
    wire n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
    wire n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645;
    wire n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653;
    wire n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661;
    wire n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;
    wire n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677;
    wire n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685;
    wire n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693;
    wire n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701;
    wire n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709;
    wire n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
    wire n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
    wire n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733;
    wire n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741;
    wire n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749;
    wire n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757;
    wire n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765;
    wire n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
    wire n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781;
    wire n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789;
    wire n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797;
    wire n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805;
    wire n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813;
    wire n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821;
    wire n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829;
    wire n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837;
    wire n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845;
    wire n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853;
    wire n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861;
    wire n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869;
    wire n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877;
    wire n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885;
    wire n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893;
    wire n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901;
    wire n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909;
    wire n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917;
    wire n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925;
    wire n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933;
    wire n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941;
    wire n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949;
    wire n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957;
    wire n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965;
    wire n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973;
    wire n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981;
    wire n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989;
    wire n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997;
    wire n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005;
    wire n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013;
    wire n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;
    wire n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029;
    wire n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037;
    wire n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045;
    wire n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053;
    wire n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061;
    wire n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069;
    wire n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077;
    wire n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085;
    wire n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093;
    wire n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101;
    wire n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109;
    wire n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117;
    wire n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125;
    wire n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133;
    wire n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141;
    wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
    wire n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157;
    wire n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165;
    wire n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
    wire n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181;
    wire n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189;
    wire n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197;
    wire n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205;
    wire n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213;
    wire n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;
    wire n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229;
    wire n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237;
    wire n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245;
    wire n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253;
    wire n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261;
    wire n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269;
    wire n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277;
    wire n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285;
    wire n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293;
    wire n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301;
    wire n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309;
    wire n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317;
    wire n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325;
    wire n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333;
    wire n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341;
    wire n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349;
    wire n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357;
    wire n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365;
    wire n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373;
    wire n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381;
    wire n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389;
    wire n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397;
    wire n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405;
    wire n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413;
    wire n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421;
    wire n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429;
    wire n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437;
    wire n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
    wire n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453;
    wire n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461;
    wire n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469;
    wire n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477;
    wire n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485;
    wire n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493;
    wire n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501;
    wire n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509;
    wire n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517;
    wire n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525;
    wire n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533;
    wire n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541;
    wire n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549;
    wire n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557;
    wire n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565;
    wire n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573;
    wire n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581;
    wire n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589;
    wire n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597;
    wire n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605;
    wire n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613;
    wire n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621;
    wire n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629;
    wire n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637;
    wire n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645;
    wire n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653;
    wire n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661;
    wire n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669;
    wire n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677;
    wire n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685;
    wire n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693;
    wire n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701;
    wire n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709;
    wire n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717;
    wire n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725;
    wire n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733;
    wire n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741;
    wire n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749;
    wire n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757;
    wire n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765;
    wire n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773;
    wire n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781;
    wire n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789;
    wire n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797;
    wire n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805;
    wire n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813;
    wire n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821;
    wire n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829;
    wire n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837;
    wire n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845;
    wire n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853;
    wire n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861;
    wire n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869;
    wire n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877;
    wire n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885;
    wire n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893;
    wire n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901;
    wire n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909;
    wire n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917;
    wire n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925;
    wire n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;
    wire n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941;
    wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
    wire n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957;
    wire n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965;
    wire n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973;
    wire n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981;
    wire n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989;
    wire n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997;
    wire n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005;
    wire n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013;
    wire n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021;
    wire n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029;
    wire n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037;
    wire n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045;
    wire n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053;
    wire n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061;
    wire n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069;
    wire n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077;
    wire n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085;
    wire n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093;
    wire n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101;
    wire n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109;
    wire n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117;
    wire n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125;
    wire n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133;
    wire n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141;
    wire n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149;
    wire n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157;
    wire n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165;
    wire n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173;
    wire n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181;
    wire n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189;
    wire n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197;
    wire n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205;
    wire n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213;
    wire n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221;
    wire n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229;
    wire n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237;
    wire n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245;
    wire n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253;
    wire n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261;
    wire n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269;
    wire n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277;
    wire n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285;
    wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
    wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
    wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
    wire n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317;
    wire n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325;
    wire n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333;
    wire n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341;
    wire n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349;
    wire n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357;
    wire n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365;
    wire n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373;
    wire n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381;
    wire n3382, n3383, n3384, n3385, n3386;
    buf g0(n33[0], 1'b0);
    buf g1(n33[1], 1'b0);
    buf g2(n33[2], 1'b0);
    buf g3(n32[4], 1'b0);
    buf g4(n32[5], 1'b0);
    buf g5(n32[6], 1'b0);
    buf g6(n32[7], 1'b0);
    not g7(n3258 ,n3262);
    not g8(n3257 ,n3265);
    not g9(n3256 ,n3268);
    not g10(n3255 ,n3367);
    or g11(n3267 ,n3252 ,n3254);
    or g12(n3266 ,n3251 ,n3253);
    nor g13(n3254 ,n3249 ,n3260);
    nor g14(n3253 ,n3248 ,n3260);
    nor g15(n3251 ,n3247 ,n3250);
    not g16(n3260 ,n3250);
    nor g17(n3250 ,n3246 ,n3256);
    not g18(n3249 ,n20[1]);
    not g19(n3248 ,n20[0]);
    not g20(n3247 ,n3269);
    not g21(n3246 ,n2[1]);
    nor g22(n3270 ,n3243 ,n3259);
    nor g23(n3269 ,n3244 ,n3259);
    or g24(n3259 ,n3245 ,n3255);
    not g25(n3245 ,n2[0]);
    not g26(n3244 ,n18[0]);
    not g27(n3243 ,n18[1]);
    or g28(n3264 ,n3240 ,n3242);
    or g29(n3263 ,n3239 ,n3241);
    nor g30(n3242 ,n3237 ,n3261);
    nor g31(n3241 ,n3235 ,n3261);
    nor g32(n3240 ,n3236 ,n3238);
    nor g33(n3239 ,n3234 ,n3238);
    not g34(n3261 ,n3238);
    nor g35(n3238 ,n3233 ,n3257);
    not g36(n3237 ,n22[1]);
    not g37(n3236 ,n3267);
    not g38(n3235 ,n22[0]);
    not g39(n3234 ,n3266);
    not g40(n3233 ,n2[2]);
    dff g41(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2661), .Q(n35[0]));
    dff g42(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2455), .Q(n35[1]));
    dff g43(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2454), .Q(n35[2]));
    dff g44(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2664), .Q(n35[3]));
    dff g45(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2663), .Q(n29[0]));
    dff g46(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2505), .Q(n29[1]));
    dff g47(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2450), .Q(n29[2]));
    dff g48(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2662), .Q(n29[3]));
    dff g49(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2660), .Q(n30[0]));
    dff g50(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2441), .Q(n30[1]));
    dff g51(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2445), .Q(n30[2]));
    dff g52(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2659), .Q(n30[3]));
    dff g53(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2439), .Q(n36[0]));
    dff g54(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2434), .Q(n36[1]));
    dff g55(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2429), .Q(n36[2]));
    dff g56(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2424), .Q(n36[3]));
    dff g57(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2658), .Q(n37[0]));
    dff g58(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2417), .Q(n37[1]));
    dff g59(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2414), .Q(n37[2]));
    dff g60(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2657), .Q(n37[3]));
    dff g61(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n38[0]));
    dff g62(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n38[1]));
    dff g63(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2026), .Q(n38[2]));
    dff g64(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n38[3]));
    dff g65(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1581), .Q(n39[0]));
    dff g66(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1580), .Q(n39[1]));
    dff g67(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1579), .Q(n39[2]));
    dff g68(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1578), .Q(n39[3]));
    dff g69(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2946), .Q(n40[0]));
    dff g70(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2948), .Q(n40[1]));
    dff g71(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2945), .Q(n40[2]));
    dff g72(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2944), .Q(n40[3]));
    dff g73(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2943), .Q(n40[4]));
    dff g74(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2942), .Q(n40[5]));
    dff g75(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2941), .Q(n40[6]));
    dff g76(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2940), .Q(n40[7]));
    dff g77(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2938), .Q(n40[8]));
    dff g78(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2939), .Q(n40[9]));
    dff g79(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2937), .Q(n40[10]));
    dff g80(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2936), .Q(n40[11]));
    dff g81(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2935), .Q(n40[12]));
    dff g82(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2934), .Q(n40[13]));
    dff g83(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3012), .Q(n40[14]));
    dff g84(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3011), .Q(n40[15]));
    dff g85(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3010), .Q(n40[16]));
    dff g86(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3009), .Q(n40[17]));
    dff g87(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3008), .Q(n40[18]));
    dff g88(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3006), .Q(n40[19]));
    dff g89(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3005), .Q(n40[20]));
    dff g90(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3004), .Q(n40[21]));
    dff g91(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3002), .Q(n40[22]));
    dff g92(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3001), .Q(n40[23]));
    dff g93(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2999), .Q(n40[24]));
    dff g94(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2998), .Q(n40[25]));
    dff g95(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2996), .Q(n40[26]));
    dff g96(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2995), .Q(n40[27]));
    dff g97(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2994), .Q(n40[28]));
    dff g98(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2993), .Q(n40[29]));
    dff g99(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2992), .Q(n40[30]));
    dff g100(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2991), .Q(n40[31]));
    dff g101(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2989), .Q(n41[0]));
    dff g102(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2990), .Q(n41[1]));
    dff g103(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2988), .Q(n41[2]));
    dff g104(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2987), .Q(n41[3]));
    dff g105(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2986), .Q(n41[4]));
    dff g106(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2985), .Q(n41[5]));
    dff g107(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2984), .Q(n41[6]));
    dff g108(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2983), .Q(n41[7]));
    dff g109(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2982), .Q(n41[8]));
    dff g110(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2981), .Q(n41[9]));
    dff g111(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2980), .Q(n41[10]));
    dff g112(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2979), .Q(n41[11]));
    dff g113(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2978), .Q(n41[12]));
    dff g114(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2977), .Q(n41[13]));
    dff g115(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3073), .Q(n41[14]));
    dff g116(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3074), .Q(n41[15]));
    dff g117(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3075), .Q(n42[0]));
    dff g118(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3076), .Q(n42[1]));
    dff g119(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3077), .Q(n42[2]));
    dff g120(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3079), .Q(n42[3]));
    dff g121(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3080), .Q(n42[4]));
    dff g122(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3081), .Q(n42[5]));
    dff g123(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2900), .Q(n42[6]));
    dff g124(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2973), .Q(n42[7]));
    dff g125(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3078), .Q(n42[8]));
    dff g126(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2972), .Q(n42[9]));
    dff g127(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2971), .Q(n42[10]));
    dff g128(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2970), .Q(n42[11]));
    dff g129(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2969), .Q(n42[12]));
    dff g130(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2967), .Q(n42[13]));
    dff g131(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2968), .Q(n42[14]));
    dff g132(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2966), .Q(n42[15]));
    dff g133(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2965), .Q(n42[16]));
    dff g134(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2964), .Q(n42[17]));
    dff g135(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2963), .Q(n42[18]));
    dff g136(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2961), .Q(n42[19]));
    dff g137(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2962), .Q(n42[20]));
    dff g138(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2960), .Q(n42[21]));
    dff g139(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2959), .Q(n42[22]));
    dff g140(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2958), .Q(n42[23]));
    dff g141(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2956), .Q(n42[24]));
    dff g142(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2957), .Q(n42[25]));
    dff g143(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2955), .Q(n42[26]));
    dff g144(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2954), .Q(n42[27]));
    dff g145(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2953), .Q(n42[28]));
    dff g146(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2952), .Q(n42[29]));
    dff g147(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2951), .Q(n42[30]));
    dff g148(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2950), .Q(n42[31]));
    dff g149(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1452), .Q(n43[0]));
    dff g150(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1453), .Q(n43[1]));
    dff g151(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1451), .Q(n43[2]));
    dff g152(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2949), .Q(n44[0]));
    dff g153(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2947), .Q(n44[1]));
    dff g154(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1577), .Q(n33[3]));
    dff g155(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1576), .Q(n33[4]));
    dff g156(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1582), .Q(n33[5]));
    dff g157(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1575), .Q(n33[6]));
    dff g158(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1397), .Q(n33[7]));
    dff g159(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n31[0]));
    dff g160(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1864), .Q(n31[1]));
    dff g161(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n31[2]));
    dff g162(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n31[3]));
    dff g163(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n31[4]));
    dff g164(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n31[5]));
    dff g165(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n31[6]));
    dff g166(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n31[7]));
    dff g167(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n32[0]));
    dff g168(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n32[1]));
    dff g169(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n32[2]));
    dff g170(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n32[3]));
    dff g171(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2928), .Q(n26[0]));
    dff g172(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2927), .Q(n26[1]));
    dff g173(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2926), .Q(n26[2]));
    dff g174(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2925), .Q(n26[3]));
    dff g175(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2924), .Q(n26[4]));
    dff g176(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2923), .Q(n26[5]));
    dff g177(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2922), .Q(n26[6]));
    dff g178(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2921), .Q(n26[7]));
    dff g179(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2920), .Q(n26[8]));
    dff g180(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2919), .Q(n26[9]));
    dff g181(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2918), .Q(n26[10]));
    dff g182(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2917), .Q(n26[11]));
    dff g183(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2916), .Q(n26[12]));
    dff g184(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2915), .Q(n26[13]));
    dff g185(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2914), .Q(n26[14]));
    dff g186(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2913), .Q(n26[15]));
    dff g187(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2912), .Q(n26[16]));
    dff g188(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2911), .Q(n26[17]));
    dff g189(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2910), .Q(n26[18]));
    dff g190(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2909), .Q(n26[19]));
    dff g191(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2908), .Q(n26[20]));
    dff g192(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2907), .Q(n26[21]));
    dff g193(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2906), .Q(n26[22]));
    dff g194(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2905), .Q(n26[23]));
    dff g195(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2904), .Q(n26[24]));
    dff g196(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2903), .Q(n26[25]));
    dff g197(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2902), .Q(n26[26]));
    dff g198(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2901), .Q(n26[27]));
    dff g199(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2932), .Q(n26[28]));
    dff g200(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2931), .Q(n26[29]));
    dff g201(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2930), .Q(n26[30]));
    dff g202(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2929), .Q(n26[31]));
    dff g203(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2665), .Q(n28));
    dff g204(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3118), .Q(n27));
    dff g205(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3232), .Q(n45[0]));
    dff g206(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3231), .Q(n45[1]));
    dff g207(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3230), .Q(n45[2]));
    dff g208(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n34[0]));
    dff g209(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n34[1]));
    dff g210(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n34[2]));
    dff g211(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n34[3]));
    dff g212(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n34[4]));
    dff g213(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n34[5]));
    dff g214(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n34[6]));
    dff g215(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n34[7]));
    dff g216(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n34[8]));
    dff g217(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n34[9]));
    dff g218(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n34[10]));
    dff g219(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n34[11]));
    dff g220(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n34[12]));
    dff g221(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n34[13]));
    dff g222(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n34[14]));
    dff g223(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n34[15]));
    dff g224(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2892), .Q(n25[0]));
    dff g225(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2891), .Q(n25[1]));
    dff g226(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2890), .Q(n25[2]));
    dff g227(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2889), .Q(n25[3]));
    dff g228(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2888), .Q(n25[4]));
    dff g229(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2887), .Q(n25[5]));
    dff g230(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2886), .Q(n25[6]));
    dff g231(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2885), .Q(n25[7]));
    dff g232(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2884), .Q(n25[8]));
    dff g233(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2883), .Q(n25[9]));
    dff g234(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2882), .Q(n25[10]));
    dff g235(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2881), .Q(n25[11]));
    dff g236(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2880), .Q(n25[12]));
    dff g237(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2879), .Q(n25[13]));
    dff g238(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2878), .Q(n25[14]));
    dff g239(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2877), .Q(n25[15]));
    dff g240(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2876), .Q(n25[16]));
    dff g241(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2875), .Q(n25[17]));
    dff g242(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2874), .Q(n25[18]));
    dff g243(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2873), .Q(n25[19]));
    dff g244(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2872), .Q(n25[20]));
    dff g245(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2871), .Q(n25[21]));
    dff g246(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2870), .Q(n25[22]));
    dff g247(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2869), .Q(n25[23]));
    dff g248(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2868), .Q(n25[24]));
    dff g249(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2867), .Q(n25[25]));
    dff g250(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2866), .Q(n25[26]));
    dff g251(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2865), .Q(n25[27]));
    dff g252(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2864), .Q(n25[28]));
    dff g253(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2863), .Q(n25[29]));
    dff g254(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2899), .Q(n25[30]));
    dff g255(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n2974), .Q(n25[31]));
    dff g256(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n46[0]));
    dff g257(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n46[1]));
    dff g258(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n46[2]));
    dff g259(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n46[3]));
    dff g260(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n46[4]));
    dff g261(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n46[5]));
    dff g262(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n46[6]));
    dff g263(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n46[7]));
    dff g264(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n46[8]));
    dff g265(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n46[9]));
    dff g266(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n47[0]));
    dff g267(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n47[1]));
    dff g268(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n47[2]));
    dff g269(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n47[3]));
    dff g270(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n47[4]));
    dff g271(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n47[5]));
    dff g272(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n47[6]));
    dff g273(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n47[7]));
    dff g274(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n47[8]));
    dff g275(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n47[9]));
    dff g276(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n48[0]));
    dff g277(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n48[1]));
    dff g278(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n48[2]));
    dff g279(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n48[3]));
    dff g280(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n48[4]));
    dff g281(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n48[5]));
    dff g282(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n48[6]));
    dff g283(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n48[7]));
    dff g284(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n48[8]));
    dff g285(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n48[9]));
    dff g286(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n49[0]));
    dff g287(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n49[1]));
    dff g288(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n49[2]));
    dff g289(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n49[3]));
    dff g290(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n49[4]));
    dff g291(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n49[5]));
    dff g292(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n49[6]));
    dff g293(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n49[7]));
    dff g294(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1767), .Q(n49[8]));
    dff g295(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n49[9]));
    dff g296(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3147), .Q(n50[0]));
    dff g297(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3152), .Q(n50[1]));
    dff g298(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3151), .Q(n50[2]));
    dff g299(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3150), .Q(n50[3]));
    dff g300(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3149), .Q(n50[4]));
    dff g301(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3148), .Q(n50[5]));
    dff g302(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3146), .Q(n50[6]));
    dff g303(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3145), .Q(n50[7]));
    dff g304(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3144), .Q(n50[8]));
    dff g305(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3143), .Q(n50[9]));
    dff g306(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3142), .Q(n50[10]));
    dff g307(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3141), .Q(n50[11]));
    dff g308(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3140), .Q(n50[12]));
    dff g309(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3139), .Q(n50[13]));
    dff g310(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3138), .Q(n50[14]));
    dff g311(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3137), .Q(n50[15]));
    dff g312(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3136), .Q(n51[0]));
    dff g313(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3135), .Q(n51[1]));
    dff g314(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3134), .Q(n51[2]));
    dff g315(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3133), .Q(n51[3]));
    dff g316(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3132), .Q(n51[4]));
    dff g317(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3131), .Q(n51[5]));
    dff g318(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3130), .Q(n51[6]));
    dff g319(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3129), .Q(n51[7]));
    dff g320(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3128), .Q(n51[8]));
    dff g321(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3127), .Q(n51[9]));
    dff g322(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3126), .Q(n51[10]));
    dff g323(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3123), .Q(n51[11]));
    dff g324(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3125), .Q(n51[12]));
    dff g325(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3124), .Q(n51[13]));
    dff g326(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3122), .Q(n51[14]));
    dff g327(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3121), .Q(n51[15]));
    dff g328(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3218), .Q(n52[0]));
    dff g329(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3217), .Q(n52[1]));
    dff g330(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3216), .Q(n52[2]));
    dff g331(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3215), .Q(n52[3]));
    dff g332(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3214), .Q(n52[4]));
    dff g333(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3213), .Q(n52[5]));
    dff g334(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3212), .Q(n52[6]));
    dff g335(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3211), .Q(n52[7]));
    dff g336(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3210), .Q(n52[8]));
    dff g337(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3209), .Q(n52[9]));
    dff g338(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3208), .Q(n52[10]));
    dff g339(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3206), .Q(n52[11]));
    dff g340(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3207), .Q(n52[12]));
    dff g341(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3205), .Q(n52[13]));
    dff g342(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3204), .Q(n52[14]));
    dff g343(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3219), .Q(n52[15]));
    dff g344(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3202), .Q(n53[0]));
    dff g345(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3201), .Q(n53[1]));
    dff g346(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3200), .Q(n53[2]));
    dff g347(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3199), .Q(n53[3]));
    dff g348(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3198), .Q(n53[4]));
    dff g349(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3197), .Q(n53[5]));
    dff g350(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3196), .Q(n53[6]));
    dff g351(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3195), .Q(n53[7]));
    dff g352(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3194), .Q(n53[8]));
    dff g353(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3191), .Q(n53[9]));
    dff g354(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3193), .Q(n53[10]));
    dff g355(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3192), .Q(n53[11]));
    dff g356(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3190), .Q(n53[12]));
    dff g357(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3189), .Q(n53[13]));
    dff g358(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3188), .Q(n53[14]));
    dff g359(.RN(1'b1), .SN(1'b1), .CK(n0), .D(n3187), .Q(n53[15]));
    or g360(n3232 ,n3229 ,n3226);
    or g361(n3231 ,n3227 ,n3225);
    or g362(n3230 ,n3228 ,n3224);
    nor g363(n3229 ,n1169 ,n3222);
    nor g364(n3228 ,n1171 ,n3222);
    nor g365(n3227 ,n1168 ,n3222);
    nor g366(n3226 ,n1854 ,n3223);
    nor g367(n3225 ,n2008 ,n3223);
    nor g368(n3224 ,n2006 ,n3223);
    not g369(n3222 ,n3223);
    nor g370(n3223 ,n2005 ,n3221);
    or g371(n3221 ,n1933 ,n3220);
    nor g372(n3220 ,n2197 ,n3203);
    or g373(n3219 ,n3023 ,n3171);
    or g374(n3218 ,n2894 ,n3155);
    or g375(n3217 ,n3039 ,n3184);
    or g376(n3216 ,n3038 ,n3185);
    or g377(n3215 ,n3037 ,n3183);
    or g378(n3214 ,n3036 ,n3182);
    or g379(n3213 ,n3035 ,n3181);
    or g380(n3212 ,n3034 ,n3180);
    or g381(n3211 ,n3033 ,n3179);
    or g382(n3210 ,n3031 ,n3178);
    or g383(n3209 ,n3030 ,n3177);
    or g384(n3208 ,n3029 ,n3176);
    or g385(n3207 ,n3027 ,n3174);
    or g386(n3206 ,n3028 ,n3175);
    or g387(n3205 ,n3026 ,n3173);
    or g388(n3204 ,n3025 ,n3172);
    nor g389(n3203 ,n3154 ,n3153);
    or g390(n3202 ,n2893 ,n3170);
    or g391(n3201 ,n3022 ,n3186);
    or g392(n3200 ,n3021 ,n3169);
    or g393(n3199 ,n3020 ,n3168);
    or g394(n3198 ,n3019 ,n3167);
    or g395(n3197 ,n3018 ,n3166);
    or g396(n3196 ,n3017 ,n3165);
    or g397(n3195 ,n3016 ,n3164);
    or g398(n3194 ,n3015 ,n3163);
    or g399(n3193 ,n3024 ,n3161);
    or g400(n3192 ,n3054 ,n3160);
    or g401(n3191 ,n3014 ,n3162);
    or g402(n3190 ,n3032 ,n3159);
    or g403(n3189 ,n3013 ,n3158);
    or g404(n3188 ,n3072 ,n3157);
    or g405(n3187 ,n3071 ,n3156);
    nor g406(n3186 ,n1026 ,n3120);
    nor g407(n3185 ,n1001 ,n3119);
    nor g408(n3184 ,n1002 ,n3119);
    nor g409(n3183 ,n1000 ,n3119);
    nor g410(n3182 ,n970 ,n3119);
    nor g411(n3181 ,n1029 ,n3119);
    nor g412(n3180 ,n992 ,n3119);
    nor g413(n3179 ,n1003 ,n3119);
    nor g414(n3178 ,n997 ,n3119);
    nor g415(n3177 ,n1004 ,n3119);
    nor g416(n3176 ,n995 ,n3119);
    nor g417(n3175 ,n989 ,n3119);
    nor g418(n3174 ,n985 ,n3119);
    nor g419(n3173 ,n990 ,n3119);
    nor g420(n3172 ,n993 ,n3119);
    nor g421(n3171 ,n973 ,n3119);
    nor g422(n3170 ,n966 ,n3120);
    nor g423(n3169 ,n1024 ,n3120);
    nor g424(n3168 ,n1023 ,n3120);
    nor g425(n3167 ,n1022 ,n3120);
    nor g426(n3166 ,n1021 ,n3120);
    nor g427(n3165 ,n1019 ,n3120);
    nor g428(n3164 ,n1017 ,n3120);
    nor g429(n3163 ,n1031 ,n3120);
    nor g430(n3162 ,n1006 ,n3120);
    nor g431(n3161 ,n1011 ,n3120);
    nor g432(n3160 ,n1020 ,n3120);
    nor g433(n3159 ,n1010 ,n3120);
    nor g434(n3158 ,n1008 ,n3120);
    nor g435(n3157 ,n1007 ,n3120);
    nor g436(n3156 ,n1005 ,n3120);
    nor g437(n3155 ,n963 ,n3119);
    or g438(n3154 ,n3114 ,n3115);
    or g439(n3153 ,n3116 ,n3117);
    or g440(n3152 ,n3070 ,n3082);
    or g441(n3151 ,n3069 ,n3083);
    or g442(n3150 ,n3068 ,n3084);
    or g443(n3149 ,n3067 ,n3085);
    or g444(n3148 ,n3066 ,n3086);
    or g445(n3147 ,n2896 ,n3112);
    or g446(n3146 ,n3065 ,n3087);
    or g447(n3145 ,n3064 ,n3088);
    or g448(n3144 ,n3063 ,n3089);
    or g449(n3143 ,n3062 ,n3090);
    or g450(n3142 ,n3061 ,n3091);
    or g451(n3141 ,n3060 ,n3092);
    or g452(n3140 ,n3059 ,n3093);
    or g453(n3139 ,n3058 ,n3094);
    or g454(n3138 ,n3057 ,n3095);
    or g455(n3137 ,n3056 ,n3096);
    or g456(n3136 ,n2895 ,n3113);
    or g457(n3135 ,n3055 ,n3097);
    or g458(n3134 ,n3053 ,n3099);
    or g459(n3133 ,n3052 ,n3098);
    or g460(n3132 ,n3051 ,n3100);
    or g461(n3131 ,n3050 ,n3101);
    or g462(n3130 ,n3049 ,n3102);
    or g463(n3129 ,n3048 ,n3103);
    or g464(n3128 ,n3047 ,n3104);
    or g465(n3127 ,n3046 ,n3105);
    or g466(n3126 ,n3045 ,n3106);
    or g467(n3125 ,n3043 ,n3108);
    or g468(n3124 ,n3042 ,n3109);
    or g469(n3123 ,n3044 ,n3107);
    or g470(n3122 ,n3041 ,n3110);
    or g471(n3121 ,n3040 ,n3111);
    or g472(n3118 ,n2933 ,n2670);
    nor g473(n3117 ,n2850 ,n2997);
    nor g474(n3116 ,n2544 ,n3000);
    nor g475(n3115 ,n2546 ,n3003);
    nor g476(n3114 ,n2548 ,n3007);
    nor g477(n3113 ,n965 ,n2975);
    nor g478(n3112 ,n968 ,n2976);
    nor g479(n3111 ,n987 ,n2975);
    nor g480(n3110 ,n982 ,n2975);
    nor g481(n3109 ,n1014 ,n2975);
    nor g482(n3108 ,n976 ,n2975);
    nor g483(n3107 ,n984 ,n2975);
    nor g484(n3106 ,n1009 ,n2975);
    nor g485(n3105 ,n1013 ,n2975);
    nor g486(n3104 ,n1033 ,n2975);
    nor g487(n3103 ,n1015 ,n2975);
    nor g488(n3102 ,n988 ,n2975);
    nor g489(n3101 ,n979 ,n2975);
    nor g490(n3100 ,n1030 ,n2975);
    nor g491(n3099 ,n981 ,n2975);
    nor g492(n3098 ,n998 ,n2975);
    nor g493(n3097 ,n986 ,n2975);
    nor g494(n3096 ,n1012 ,n2976);
    nor g495(n3095 ,n974 ,n2976);
    nor g496(n3094 ,n991 ,n2976);
    nor g497(n3093 ,n1025 ,n2976);
    nor g498(n3092 ,n1016 ,n2976);
    nor g499(n3091 ,n971 ,n2976);
    nor g500(n3090 ,n978 ,n2976);
    nor g501(n3089 ,n972 ,n2976);
    nor g502(n3088 ,n1034 ,n2976);
    nor g503(n3087 ,n1028 ,n2976);
    nor g504(n3086 ,n1035 ,n2976);
    nor g505(n3085 ,n1018 ,n2976);
    nor g506(n3084 ,n999 ,n2976);
    nor g507(n3083 ,n969 ,n2976);
    nor g508(n3082 ,n975 ,n2976);
    or g509(n3120 ,n1599 ,n2897);
    or g510(n3119 ,n1598 ,n2898);
    or g511(n3081 ,n2462 ,n2713);
    or g512(n3080 ,n2492 ,n2710);
    or g513(n3079 ,n2464 ,n2714);
    or g514(n3078 ,n2456 ,n2716);
    or g515(n3077 ,n2517 ,n2715);
    or g516(n3076 ,n2468 ,n2717);
    or g517(n3075 ,n2470 ,n2718);
    or g518(n3074 ,n2472 ,n2719);
    or g519(n3073 ,n2474 ,n2720);
    nor g520(n3072 ,n855 ,n2858);
    nor g521(n3071 ,n561 ,n2858);
    nor g522(n3070 ,n796 ,n2862);
    nor g523(n3069 ,n564 ,n2862);
    nor g524(n3068 ,n851 ,n2862);
    nor g525(n3067 ,n613 ,n2862);
    nor g526(n3066 ,n1302 ,n2862);
    nor g527(n3065 ,n1303 ,n2862);
    nor g528(n3064 ,n1272 ,n2862);
    nor g529(n3063 ,n856 ,n2862);
    nor g530(n3062 ,n793 ,n2862);
    nor g531(n3061 ,n1307 ,n2862);
    nor g532(n3060 ,n1309 ,n2862);
    nor g533(n3059 ,n864 ,n2862);
    nor g534(n3058 ,n714 ,n2862);
    nor g535(n3057 ,n894 ,n2862);
    nor g536(n3056 ,n827 ,n2862);
    nor g537(n3055 ,n683 ,n2856);
    nor g538(n3054 ,n938 ,n2858);
    nor g539(n3053 ,n742 ,n2856);
    nor g540(n3052 ,n1333 ,n2856);
    nor g541(n3051 ,n597 ,n2856);
    nor g542(n3050 ,n805 ,n2856);
    nor g543(n3049 ,n584 ,n2856);
    nor g544(n3048 ,n721 ,n2856);
    nor g545(n3047 ,n792 ,n2856);
    nor g546(n3046 ,n808 ,n2856);
    nor g547(n3045 ,n1288 ,n2856);
    nor g548(n3044 ,n889 ,n2856);
    nor g549(n3043 ,n1258 ,n2856);
    nor g550(n3042 ,n634 ,n2856);
    nor g551(n3041 ,n725 ,n2856);
    nor g552(n3040 ,n704 ,n2856);
    nor g553(n3039 ,n563 ,n2860);
    nor g554(n3038 ,n846 ,n2860);
    nor g555(n3037 ,n556 ,n2860);
    nor g556(n3036 ,n774 ,n2860);
    nor g557(n3035 ,n839 ,n2860);
    nor g558(n3034 ,n1259 ,n2860);
    nor g559(n3033 ,n812 ,n2860);
    nor g560(n3032 ,n892 ,n2858);
    nor g561(n3031 ,n862 ,n2860);
    nor g562(n3030 ,n929 ,n2860);
    nor g563(n3029 ,n931 ,n2860);
    nor g564(n3028 ,n879 ,n2860);
    nor g565(n3027 ,n588 ,n2860);
    nor g566(n3026 ,n798 ,n2860);
    nor g567(n3025 ,n645 ,n2860);
    nor g568(n3024 ,n587 ,n2858);
    nor g569(n3023 ,n691 ,n2860);
    nor g570(n3022 ,n1267 ,n2858);
    nor g571(n3021 ,n871 ,n2858);
    nor g572(n3020 ,n887 ,n2858);
    nor g573(n3019 ,n859 ,n2858);
    nor g574(n3018 ,n868 ,n2858);
    nor g575(n3017 ,n567 ,n2858);
    nor g576(n3016 ,n717 ,n2858);
    nor g577(n3015 ,n866 ,n2858);
    nor g578(n3014 ,n723 ,n2858);
    nor g579(n3013 ,n939 ,n2858);
    or g580(n3012 ,n2538 ,n2852);
    or g581(n3011 ,n2535 ,n2853);
    or g582(n3010 ,n2532 ,n2629);
    or g583(n3009 ,n2530 ,n2748);
    or g584(n3008 ,n2528 ,n2747);
    or g585(n3007 ,n1838 ,n2847);
    or g586(n3006 ,n2526 ,n2746);
    or g587(n3005 ,n2525 ,n2745);
    or g588(n3004 ,n2522 ,n2744);
    or g589(n3003 ,n1488 ,n2848);
    or g590(n3002 ,n2520 ,n2743);
    or g591(n3001 ,n2518 ,n2742);
    or g592(n3000 ,n1484 ,n2849);
    or g593(n2999 ,n2515 ,n2741);
    or g594(n2998 ,n2513 ,n2739);
    or g595(n2997 ,n1479 ,n2851);
    or g596(n2996 ,n2512 ,n2740);
    or g597(n2995 ,n2509 ,n2738);
    or g598(n2994 ,n2507 ,n2737);
    or g599(n2993 ,n2503 ,n2736);
    or g600(n2992 ,n2501 ,n2735);
    or g601(n2991 ,n2499 ,n2734);
    or g602(n2990 ,n2558 ,n2732);
    or g603(n2989 ,n2498 ,n2733);
    or g604(n2988 ,n2368 ,n2673);
    or g605(n2987 ,n2496 ,n2731);
    or g606(n2986 ,n2494 ,n2730);
    or g607(n2985 ,n2537 ,n2728);
    or g608(n2984 ,n2491 ,n2729);
    or g609(n2983 ,n2488 ,n2727);
    or g610(n2982 ,n2486 ,n2726);
    or g611(n2981 ,n2484 ,n2725);
    or g612(n2980 ,n2482 ,n2724);
    or g613(n2979 ,n2480 ,n2723);
    or g614(n2978 ,n2478 ,n2722);
    or g615(n2977 ,n2476 ,n2721);
    or g616(n2974 ,n2843 ,n2778);
    or g617(n2973 ,n2458 ,n2711);
    or g618(n2972 ,n2451 ,n2709);
    or g619(n2971 ,n2460 ,n2854);
    or g620(n2970 ,n2449 ,n2708);
    or g621(n2969 ,n2447 ,n2707);
    or g622(n2968 ,n2442 ,n2705);
    or g623(n2967 ,n2444 ,n2706);
    or g624(n2966 ,n2438 ,n2704);
    or g625(n2965 ,n2436 ,n2703);
    or g626(n2964 ,n2433 ,n2702);
    or g627(n2963 ,n2431 ,n2701);
    or g628(n2962 ,n2426 ,n2699);
    or g629(n2961 ,n2428 ,n2700);
    or g630(n2960 ,n2423 ,n2698);
    or g631(n2959 ,n2421 ,n2697);
    or g632(n2958 ,n2419 ,n2696);
    or g633(n2957 ,n2413 ,n2694);
    or g634(n2956 ,n2416 ,n2695);
    or g635(n2955 ,n2411 ,n2693);
    or g636(n2954 ,n2409 ,n2692);
    or g637(n2953 ,n2407 ,n2691);
    or g638(n2952 ,n2405 ,n2690);
    or g639(n2951 ,n2403 ,n2688);
    or g640(n2950 ,n2401 ,n2687);
    or g641(n2949 ,n2397 ,n2686);
    or g642(n2948 ,n2394 ,n2684);
    or g643(n2947 ,n2393 ,n2685);
    or g644(n2946 ,n2400 ,n2689);
    or g645(n2945 ,n2390 ,n2682);
    or g646(n2944 ,n2388 ,n2683);
    or g647(n2943 ,n2386 ,n2681);
    or g648(n2942 ,n2382 ,n2680);
    or g649(n2941 ,n2381 ,n2679);
    or g650(n2940 ,n2379 ,n2678);
    or g651(n2939 ,n2375 ,n2676);
    or g652(n2938 ,n2376 ,n2677);
    or g653(n2937 ,n2373 ,n2675);
    or g654(n2936 ,n2371 ,n2674);
    or g655(n2935 ,n2369 ,n2672);
    or g656(n2934 ,n2366 ,n2671);
    nor g657(n2933 ,n539 ,n2842);
    or g658(n2932 ,n2841 ,n2669);
    or g659(n2931 ,n2840 ,n2668);
    or g660(n2930 ,n2839 ,n2667);
    or g661(n2929 ,n2838 ,n2666);
    or g662(n2928 ,n2837 ,n2656);
    or g663(n2927 ,n2836 ,n2655);
    or g664(n2926 ,n2835 ,n2654);
    or g665(n2925 ,n2834 ,n2653);
    or g666(n2924 ,n2833 ,n2652);
    or g667(n2923 ,n2832 ,n2651);
    or g668(n2922 ,n2831 ,n2650);
    or g669(n2921 ,n2830 ,n2649);
    or g670(n2920 ,n2829 ,n2648);
    or g671(n2919 ,n2828 ,n2647);
    or g672(n2918 ,n2827 ,n2646);
    or g673(n2917 ,n2826 ,n2645);
    or g674(n2916 ,n2825 ,n2644);
    or g675(n2915 ,n2824 ,n2643);
    or g676(n2914 ,n2823 ,n2642);
    or g677(n2913 ,n2822 ,n2641);
    or g678(n2912 ,n2821 ,n2640);
    or g679(n2911 ,n2820 ,n2639);
    or g680(n2910 ,n2819 ,n2638);
    or g681(n2909 ,n2818 ,n2637);
    or g682(n2908 ,n2817 ,n2636);
    or g683(n2907 ,n2816 ,n2635);
    or g684(n2906 ,n2815 ,n2634);
    or g685(n2905 ,n2814 ,n2633);
    or g686(n2904 ,n2813 ,n2632);
    or g687(n2903 ,n2812 ,n2631);
    or g688(n2902 ,n2811 ,n2630);
    or g689(n2901 ,n2810 ,n2749);
    or g690(n2900 ,n2452 ,n2712);
    or g691(n2899 ,n2777 ,n2779);
    or g692(n2898 ,n544 ,n2859);
    or g693(n2897 ,n537 ,n2857);
    nor g694(n2896 ,n50[0] ,n2862);
    nor g695(n2895 ,n51[0] ,n2856);
    nor g696(n2894 ,n52[0] ,n2860);
    nor g697(n2893 ,n53[0] ,n2858);
    or g698(n2892 ,n2776 ,n2809);
    or g699(n2891 ,n2775 ,n2808);
    or g700(n2890 ,n2774 ,n2807);
    or g701(n2889 ,n2773 ,n2806);
    or g702(n2888 ,n2772 ,n2805);
    or g703(n2887 ,n2771 ,n2804);
    or g704(n2886 ,n2770 ,n2803);
    or g705(n2885 ,n2769 ,n2802);
    or g706(n2884 ,n2768 ,n2801);
    or g707(n2883 ,n2767 ,n2800);
    or g708(n2882 ,n2766 ,n2799);
    or g709(n2881 ,n2765 ,n2798);
    or g710(n2880 ,n2764 ,n2797);
    or g711(n2879 ,n2763 ,n2796);
    or g712(n2878 ,n2846 ,n2795);
    or g713(n2877 ,n2762 ,n2794);
    or g714(n2876 ,n2761 ,n2793);
    or g715(n2875 ,n2760 ,n2792);
    or g716(n2874 ,n2845 ,n2791);
    or g717(n2873 ,n2759 ,n2790);
    or g718(n2872 ,n2758 ,n2789);
    or g719(n2871 ,n2757 ,n2788);
    or g720(n2870 ,n2844 ,n2787);
    or g721(n2869 ,n2756 ,n2786);
    or g722(n2868 ,n2755 ,n2785);
    or g723(n2867 ,n2754 ,n2784);
    or g724(n2866 ,n2753 ,n2783);
    or g725(n2865 ,n2752 ,n2782);
    or g726(n2864 ,n2751 ,n2781);
    or g727(n2863 ,n2750 ,n2780);
    or g728(n2976 ,n1935 ,n2861);
    or g729(n2975 ,n1934 ,n2855);
    not g730(n2862 ,n2861);
    not g731(n2860 ,n2859);
    not g732(n2858 ,n2857);
    not g733(n2856 ,n2855);
    or g734(n2854 ,n2258 ,n2504);
    or g735(n2853 ,n2318 ,n2533);
    or g736(n2852 ,n2322 ,n2536);
    or g737(n2851 ,n1814 ,n2541);
    or g738(n2850 ,n1480 ,n2542);
    or g739(n2849 ,n1817 ,n2543);
    or g740(n2848 ,n1819 ,n2545);
    or g741(n2847 ,n1548 ,n2547);
    nor g742(n2846 ,n1215 ,n2625);
    nor g743(n2845 ,n1149 ,n2625);
    nor g744(n2844 ,n1178 ,n2625);
    nor g745(n2843 ,n1249 ,n2625);
    or g746(n2842 ,n1197 ,n2628);
    nor g747(n2841 ,n1163 ,n2497);
    nor g748(n2840 ,n1232 ,n2497);
    nor g749(n2839 ,n1057 ,n2497);
    nor g750(n2838 ,n1111 ,n2497);
    nor g751(n2837 ,n1239 ,n2497);
    nor g752(n2836 ,n1113 ,n2497);
    nor g753(n2835 ,n1245 ,n2497);
    nor g754(n2834 ,n1066 ,n2497);
    nor g755(n2833 ,n1069 ,n2497);
    nor g756(n2832 ,n1065 ,n2497);
    nor g757(n2831 ,n1058 ,n2497);
    nor g758(n2830 ,n1150 ,n2497);
    nor g759(n2829 ,n1214 ,n2497);
    nor g760(n2828 ,n1096 ,n2497);
    nor g761(n2827 ,n1103 ,n2497);
    nor g762(n2826 ,n1094 ,n2497);
    nor g763(n2825 ,n1132 ,n2497);
    nor g764(n2824 ,n1107 ,n2497);
    nor g765(n2823 ,n1138 ,n2497);
    nor g766(n2822 ,n1185 ,n2497);
    nor g767(n2821 ,n1182 ,n2497);
    nor g768(n2820 ,n1237 ,n2497);
    nor g769(n2819 ,n1221 ,n2497);
    nor g770(n2818 ,n1133 ,n2497);
    nor g771(n2817 ,n1165 ,n2497);
    nor g772(n2816 ,n1052 ,n2497);
    nor g773(n2815 ,n1090 ,n2497);
    nor g774(n2814 ,n1211 ,n2497);
    nor g775(n2813 ,n1143 ,n2497);
    nor g776(n2812 ,n1189 ,n2497);
    nor g777(n2811 ,n1190 ,n2497);
    nor g778(n2810 ,n1072 ,n2497);
    nor g779(n2809 ,n901 ,n2624);
    nor g780(n2808 ,n708 ,n2624);
    nor g781(n2807 ,n697 ,n2624);
    nor g782(n2806 ,n877 ,n2624);
    nor g783(n2805 ,n787 ,n2624);
    nor g784(n2804 ,n895 ,n2624);
    nor g785(n2803 ,n825 ,n2624);
    nor g786(n2802 ,n716 ,n2624);
    nor g787(n2801 ,n574 ,n2624);
    nor g788(n2800 ,n620 ,n2624);
    nor g789(n2799 ,n705 ,n2624);
    nor g790(n2798 ,n1300 ,n2624);
    nor g791(n2797 ,n596 ,n2624);
    nor g792(n2796 ,n850 ,n2624);
    nor g793(n2795 ,n809 ,n2624);
    nor g794(n2794 ,n678 ,n2624);
    nor g795(n2793 ,n664 ,n2624);
    nor g796(n2792 ,n577 ,n2624);
    nor g797(n2791 ,n600 ,n2624);
    nor g798(n2790 ,n874 ,n2624);
    nor g799(n2789 ,n633 ,n2624);
    nor g800(n2788 ,n566 ,n2624);
    nor g801(n2787 ,n730 ,n2624);
    nor g802(n2786 ,n803 ,n2624);
    nor g803(n2785 ,n914 ,n2624);
    nor g804(n2784 ,n845 ,n2624);
    nor g805(n2783 ,n776 ,n2624);
    nor g806(n2782 ,n608 ,n2624);
    nor g807(n2781 ,n737 ,n2624);
    nor g808(n2780 ,n817 ,n2624);
    nor g809(n2779 ,n1275 ,n2624);
    nor g810(n2778 ,n1338 ,n2624);
    nor g811(n2777 ,n1251 ,n2625);
    nor g812(n2776 ,n1079 ,n2625);
    nor g813(n2775 ,n1095 ,n2625);
    nor g814(n2774 ,n1120 ,n2625);
    nor g815(n2773 ,n1076 ,n2625);
    nor g816(n2772 ,n1088 ,n2625);
    nor g817(n2771 ,n1105 ,n2625);
    nor g818(n2770 ,n1135 ,n2625);
    nor g819(n2769 ,n1157 ,n2625);
    nor g820(n2768 ,n1184 ,n2625);
    nor g821(n2767 ,n1201 ,n2625);
    nor g822(n2766 ,n1100 ,n2625);
    nor g823(n2765 ,n1235 ,n2625);
    nor g824(n2764 ,n1241 ,n2625);
    nor g825(n2763 ,n1073 ,n2625);
    nor g826(n2762 ,n1082 ,n2625);
    nor g827(n2761 ,n1220 ,n2625);
    nor g828(n2760 ,n1060 ,n2625);
    nor g829(n2759 ,n1128 ,n2625);
    nor g830(n2758 ,n1187 ,n2625);
    nor g831(n2757 ,n1114 ,n2625);
    nor g832(n2756 ,n1175 ,n2625);
    nor g833(n2755 ,n1246 ,n2625);
    nor g834(n2754 ,n1248 ,n2625);
    nor g835(n2753 ,n1181 ,n2625);
    nor g836(n2752 ,n1074 ,n2625);
    nor g837(n2751 ,n1110 ,n2625);
    nor g838(n2750 ,n1126 ,n2625);
    nor g839(n2861 ,n1562 ,n2626);
    nor g840(n2859 ,n1563 ,n2626);
    nor g841(n2857 ,n1564 ,n2626);
    nor g842(n2855 ,n1565 ,n2626);
    or g843(n2749 ,n2550 ,n2582);
    or g844(n2748 ,n2312 ,n2529);
    or g845(n2747 ,n2309 ,n2527);
    or g846(n2746 ,n1955 ,n2523);
    or g847(n2745 ,n2303 ,n2524);
    or g848(n2744 ,n1953 ,n2521);
    or g849(n2743 ,n1952 ,n2519);
    or g850(n2742 ,n2295 ,n2516);
    or g851(n2741 ,n2291 ,n2514);
    or g852(n2740 ,n2284 ,n2511);
    or g853(n2739 ,n2288 ,n2510);
    or g854(n2738 ,n2281 ,n2508);
    or g855(n2737 ,n1967 ,n2506);
    or g856(n2736 ,n2274 ,n2502);
    or g857(n2735 ,n2270 ,n2500);
    or g858(n2734 ,n2365 ,n2534);
    or g859(n2733 ,n2254 ,n2549);
    or g860(n2732 ,n2263 ,n2622);
    or g861(n2731 ,n2119 ,n2495);
    or g862(n2730 ,n2255 ,n2493);
    or g863(n2729 ,n2249 ,n2489);
    or g864(n2728 ,n1982 ,n2490);
    or g865(n2727 ,n2247 ,n2487);
    or g866(n2726 ,n2244 ,n2485);
    or g867(n2725 ,n2241 ,n2483);
    or g868(n2724 ,n2238 ,n2481);
    or g869(n2723 ,n2236 ,n2479);
    or g870(n2722 ,n2232 ,n2477);
    or g871(n2721 ,n2228 ,n2475);
    or g872(n2720 ,n2225 ,n2473);
    or g873(n2719 ,n2233 ,n2471);
    or g874(n2718 ,n2219 ,n2395);
    or g875(n2717 ,n2216 ,n2467);
    or g876(n2716 ,n2224 ,n2469);
    or g877(n2715 ,n1956 ,n2466);
    or g878(n2714 ,n2218 ,n2465);
    or g879(n2713 ,n2204 ,n2461);
    or g880(n2712 ,n2201 ,n2459);
    or g881(n2711 ,n1986 ,n2457);
    or g882(n2710 ,n2208 ,n2463);
    or g883(n2709 ,n2220 ,n2453);
    or g884(n2708 ,n2340 ,n2448);
    or g885(n2707 ,n1993 ,n2446);
    or g886(n2706 ,n2345 ,n2443);
    or g887(n2705 ,n2349 ,n2440);
    or g888(n2704 ,n2352 ,n2437);
    or g889(n2703 ,n2354 ,n2435);
    or g890(n2702 ,n2358 ,n2432);
    or g891(n2701 ,n1887 ,n2430);
    or g892(n2700 ,n1855 ,n2427);
    or g893(n2699 ,n1930 ,n2425);
    or g894(n2698 ,n1929 ,n2422);
    or g895(n2697 ,n1928 ,n2420);
    or g896(n2696 ,n1927 ,n2418);
    or g897(n2695 ,n2177 ,n2415);
    or g898(n2694 ,n2174 ,n2412);
    or g899(n2693 ,n1924 ,n2410);
    or g900(n2692 ,n2168 ,n2408);
    or g901(n2691 ,n2165 ,n2406);
    or g902(n2690 ,n2162 ,n2404);
    or g903(n2689 ,n2153 ,n2398);
    or g904(n2688 ,n2159 ,n2402);
    or g905(n2687 ,n2156 ,n2399);
    or g906(n2686 ,n2149 ,n2396);
    or g907(n2685 ,n1916 ,n2392);
    or g908(n2684 ,n2144 ,n2391);
    or g909(n2683 ,n2137 ,n2387);
    or g910(n2682 ,n1914 ,n2389);
    or g911(n2681 ,n2134 ,n2385);
    or g912(n2680 ,n2131 ,n2384);
    or g913(n2679 ,n2125 ,n2380);
    or g914(n2678 ,n2123 ,n2378);
    or g915(n2677 ,n2118 ,n2377);
    or g916(n2676 ,n2114 ,n2374);
    or g917(n2675 ,n2111 ,n2372);
    or g918(n2674 ,n1903 ,n2370);
    or g919(n2673 ,n2259 ,n2539);
    or g920(n2672 ,n1902 ,n2367);
    or g921(n2671 ,n1901 ,n2383);
    nor g922(n2670 ,n1549 ,n2627);
    or g923(n2669 ,n2581 ,n2613);
    or g924(n2668 ,n2580 ,n2612);
    or g925(n2667 ,n2579 ,n2611);
    or g926(n2666 ,n2578 ,n2610);
    or g927(n2665 ,n2540 ,n2004);
    or g928(n2664 ,n525 ,n2620);
    or g929(n2663 ,n534 ,n2619);
    or g930(n2662 ,n525 ,n2618);
    or g931(n2661 ,n534 ,n2621);
    or g932(n2660 ,n1936 ,n2617);
    or g933(n2659 ,n1937 ,n2616);
    or g934(n2658 ,n1936 ,n2615);
    or g935(n2657 ,n1937 ,n2614);
    or g936(n2656 ,n2577 ,n2609);
    or g937(n2655 ,n2576 ,n2608);
    or g938(n2654 ,n2575 ,n2607);
    or g939(n2653 ,n2574 ,n2606);
    or g940(n2652 ,n2573 ,n2605);
    or g941(n2651 ,n2572 ,n2604);
    or g942(n2650 ,n2571 ,n2603);
    or g943(n2649 ,n2570 ,n2602);
    or g944(n2648 ,n2569 ,n2601);
    or g945(n2647 ,n2568 ,n2600);
    or g946(n2646 ,n2567 ,n2599);
    or g947(n2645 ,n2566 ,n2598);
    or g948(n2644 ,n2565 ,n2597);
    or g949(n2643 ,n2564 ,n2596);
    or g950(n2642 ,n2563 ,n2595);
    or g951(n2641 ,n2562 ,n2594);
    or g952(n2640 ,n2561 ,n2593);
    or g953(n2639 ,n2560 ,n2592);
    or g954(n2638 ,n2559 ,n2591);
    or g955(n2637 ,n2623 ,n2590);
    or g956(n2636 ,n2557 ,n2589);
    or g957(n2635 ,n2556 ,n2588);
    or g958(n2634 ,n2555 ,n2587);
    or g959(n2633 ,n2554 ,n2586);
    or g960(n2632 ,n2553 ,n2585);
    or g961(n2631 ,n2552 ,n2584);
    or g962(n2630 ,n2551 ,n2583);
    or g963(n2629 ,n1959 ,n2531);
    not g964(n2628 ,n2627);
    not g965(n2624 ,n2625);
    nor g966(n2623 ,n1091 ,n2192);
    or g967(n2622 ,n2262 ,n2013);
    nor g968(n2621 ,n1032 ,n2195);
    nor g969(n2620 ,n977 ,n2196);
    nor g970(n2619 ,n1240 ,n2195);
    nor g971(n2618 ,n1064 ,n2196);
    nor g972(n2617 ,n1210 ,n2195);
    nor g973(n2616 ,n1205 ,n2196);
    nor g974(n2615 ,n1044 ,n2195);
    nor g975(n2614 ,n1039 ,n2196);
    nor g976(n2613 ,n1101 ,n2194);
    nor g977(n2612 ,n1109 ,n2194);
    nor g978(n2611 ,n1118 ,n2194);
    nor g979(n2610 ,n1152 ,n2194);
    nor g980(n2609 ,n1250 ,n2194);
    nor g981(n2608 ,n1253 ,n2194);
    nor g982(n2607 ,n1180 ,n2194);
    nor g983(n2606 ,n1116 ,n2194);
    nor g984(n2605 ,n1238 ,n2194);
    nor g985(n2604 ,n1130 ,n2194);
    nor g986(n2603 ,n1097 ,n2194);
    nor g987(n2602 ,n1200 ,n2194);
    nor g988(n2601 ,n1242 ,n2194);
    nor g989(n2600 ,n1055 ,n2194);
    nor g990(n2599 ,n1193 ,n2194);
    nor g991(n2598 ,n1188 ,n2194);
    nor g992(n2597 ,n1183 ,n2194);
    nor g993(n2596 ,n1172 ,n2194);
    nor g994(n2595 ,n1177 ,n2194);
    nor g995(n2594 ,n1125 ,n2194);
    nor g996(n2593 ,n1252 ,n2194);
    nor g997(n2592 ,n1199 ,n2194);
    nor g998(n2591 ,n1159 ,n2194);
    nor g999(n2590 ,n1154 ,n2194);
    nor g1000(n2589 ,n1206 ,n2194);
    nor g1001(n2588 ,n1085 ,n2194);
    nor g1002(n2587 ,n1099 ,n2194);
    nor g1003(n2586 ,n1137 ,n2194);
    nor g1004(n2585 ,n1131 ,n2194);
    nor g1005(n2584 ,n1117 ,n2194);
    nor g1006(n2583 ,n1122 ,n2194);
    nor g1007(n2582 ,n1089 ,n2194);
    nor g1008(n2581 ,n1166 ,n2192);
    nor g1009(n2580 ,n1084 ,n2192);
    nor g1010(n2579 ,n1162 ,n2192);
    nor g1011(n2578 ,n1213 ,n2192);
    nor g1012(n2577 ,n1158 ,n2192);
    nor g1013(n2576 ,n1191 ,n2192);
    nor g1014(n2575 ,n1233 ,n2192);
    nor g1015(n2574 ,n1086 ,n2192);
    nor g1016(n2573 ,n1080 ,n2192);
    nor g1017(n2572 ,n1081 ,n2192);
    nor g1018(n2571 ,n1164 ,n2192);
    nor g1019(n2570 ,n1225 ,n2192);
    nor g1020(n2569 ,n1056 ,n2192);
    nor g1021(n2568 ,n1108 ,n2192);
    nor g1022(n2567 ,n1229 ,n2192);
    nor g1023(n2566 ,n1104 ,n2192);
    nor g1024(n2565 ,n1167 ,n2192);
    nor g1025(n2564 ,n1209 ,n2192);
    nor g1026(n2563 ,n1144 ,n2192);
    nor g1027(n2562 ,n1234 ,n2192);
    nor g1028(n2561 ,n1141 ,n2192);
    nor g1029(n2560 ,n1151 ,n2192);
    nor g1030(n2559 ,n1106 ,n2192);
    or g1031(n2558 ,n1969 ,n2261);
    nor g1032(n2557 ,n1236 ,n2192);
    nor g1033(n2556 ,n1136 ,n2192);
    nor g1034(n2555 ,n1145 ,n2192);
    nor g1035(n2554 ,n1228 ,n2192);
    nor g1036(n2553 ,n1148 ,n2192);
    nor g1037(n2552 ,n1247 ,n2192);
    nor g1038(n2551 ,n1075 ,n2192);
    nor g1039(n2550 ,n1134 ,n2192);
    or g1040(n2549 ,n1971 ,n2264);
    or g1041(n2548 ,n1899 ,n2034);
    or g1042(n2547 ,n1477 ,n2033);
    or g1043(n2546 ,n1543 ,n2032);
    or g1044(n2545 ,n1895 ,n2031);
    or g1045(n2544 ,n1486 ,n2030);
    or g1046(n2543 ,n1892 ,n2029);
    or g1047(n2542 ,n1511 ,n2028);
    or g1048(n2541 ,n1888 ,n2027);
    nor g1049(n2540 ,n537 ,n2336);
    or g1050(n2539 ,n2010 ,n2115);
    or g1051(n2538 ,n2323 ,n2100);
    or g1052(n2537 ,n2252 ,n2022);
    or g1053(n2536 ,n1962 ,n2321);
    or g1054(n2535 ,n2319 ,n2098);
    or g1055(n2534 ,n1991 ,n2266);
    or g1056(n2533 ,n1960 ,n2317);
    or g1057(n2532 ,n2315 ,n2316);
    or g1058(n2531 ,n2096 ,n2314);
    or g1059(n2530 ,n2313 ,n2095);
    or g1060(n2529 ,n1958 ,n2311);
    or g1061(n2528 ,n2310 ,n2094);
    or g1062(n2527 ,n1957 ,n2308);
    or g1063(n2526 ,n2307 ,n2191);
    or g1064(n2525 ,n2304 ,n2092);
    or g1065(n2524 ,n1954 ,n2302);
    or g1066(n2523 ,n2306 ,n2305);
    or g1067(n2522 ,n2301 ,n2091);
    or g1068(n2521 ,n2300 ,n2299);
    or g1069(n2520 ,n2297 ,n2298);
    or g1070(n2519 ,n2090 ,n2296);
    or g1071(n2518 ,n1951 ,n2089);
    or g1072(n2517 ,n2214 ,n2215);
    or g1073(n2516 ,n2294 ,n2293);
    or g1074(n2515 ,n2292 ,n2088);
    or g1075(n2514 ,n1950 ,n2290);
    or g1076(n2513 ,n2289 ,n2087);
    or g1077(n2512 ,n2286 ,n2086);
    or g1078(n2511 ,n1965 ,n2283);
    or g1079(n2510 ,n1964 ,n2287);
    or g1080(n2509 ,n2282 ,n2085);
    or g1081(n2508 ,n1966 ,n2280);
    or g1082(n2507 ,n2279 ,n2084);
    or g1083(n2506 ,n2277 ,n2276);
    or g1084(n2505 ,n531 ,n2329);
    or g1085(n2504 ,n2278 ,n2082);
    or g1086(n2503 ,n2275 ,n2081);
    or g1087(n2502 ,n1968 ,n2273);
    or g1088(n2501 ,n2271 ,n2080);
    or g1089(n2500 ,n1908 ,n2269);
    or g1090(n2499 ,n2268 ,n2079);
    or g1091(n2498 ,n2265 ,n2025);
    nor g1092(n2627 ,n1573 ,n2193);
    or g1093(n2626 ,n945 ,n2197);
    nor g1094(n2625 ,n44[1] ,n2192);
    or g1095(n2496 ,n1963 ,n2126);
    or g1096(n2495 ,n2023 ,n2142);
    or g1097(n2494 ,n2256 ,n2011);
    or g1098(n2493 ,n1997 ,n2202);
    or g1099(n2492 ,n2211 ,n2210);
    or g1100(n2491 ,n2251 ,n2024);
    or g1101(n2490 ,n2209 ,n2129);
    or g1102(n2489 ,n1973 ,n2250);
    or g1103(n2488 ,n2248 ,n2021);
    or g1104(n2487 ,n1974 ,n2246);
    or g1105(n2486 ,n2245 ,n2020);
    or g1106(n2485 ,n1975 ,n2243);
    or g1107(n2484 ,n2242 ,n2019);
    or g1108(n2483 ,n1976 ,n2240);
    or g1109(n2482 ,n2239 ,n2018);
    or g1110(n2481 ,n1977 ,n2237);
    or g1111(n2480 ,n1978 ,n2017);
    or g1112(n2479 ,n2235 ,n2234);
    or g1113(n2478 ,n1979 ,n2016);
    or g1114(n2477 ,n2230 ,n2231);
    or g1115(n2476 ,n1980 ,n2229);
    or g1116(n2475 ,n2227 ,n2015);
    or g1117(n2474 ,n1981 ,n2226);
    or g1118(n2473 ,n2348 ,n2012);
    or g1119(n2472 ,n2223 ,n2014);
    or g1120(n2471 ,n1984 ,n2222);
    or g1121(n2470 ,n2221 ,n2083);
    or g1122(n2469 ,n1972 ,n2072);
    or g1123(n2468 ,n1904 ,n2257);
    or g1124(n2467 ,n2078 ,n2272);
    or g1125(n2466 ,n2097 ,n2253);
    or g1126(n2465 ,n1985 ,n2099);
    or g1127(n2464 ,n2213 ,n2212);
    or g1128(n2463 ,n1990 ,n2076);
    or g1129(n2462 ,n2207 ,n2206);
    or g1130(n2461 ,n1987 ,n2075);
    or g1131(n2460 ,n1961 ,n2285);
    or g1132(n2459 ,n2199 ,n2200);
    or g1133(n2458 ,n2267 ,n2205);
    or g1134(n2457 ,n2077 ,n2217);
    or g1135(n2456 ,n2198 ,n2105);
    or g1136(n2455 ,n531 ,n2330);
    or g1137(n2454 ,n528 ,n2331);
    or g1138(n2453 ,n1988 ,n2203);
    or g1139(n2452 ,n1989 ,n2073);
    or g1140(n2451 ,n2337 ,n2074);
    or g1141(n2450 ,n528 ,n2328);
    or g1142(n2449 ,n2338 ,n2339);
    or g1143(n2448 ,n1992 ,n2071);
    or g1144(n2447 ,n2341 ,n2342);
    or g1145(n2446 ,n2070 ,n2343);
    or g1146(n2445 ,n1849 ,n2326);
    or g1147(n2444 ,n1994 ,n2344);
    or g1148(n2443 ,n2069 ,n2346);
    or g1149(n2442 ,n2347 ,n2068);
    or g1150(n2441 ,n1850 ,n2327);
    or g1151(n2440 ,n1995 ,n2350);
    or g1152(n2439 ,n2003 ,n2335);
    or g1153(n2438 ,n1996 ,n2351);
    or g1154(n2437 ,n2067 ,n2353);
    or g1155(n2436 ,n1998 ,n2066);
    or g1156(n2435 ,n2355 ,n2356);
    or g1157(n2434 ,n2002 ,n2334);
    or g1158(n2433 ,n1999 ,n2357);
    or g1159(n2432 ,n2359 ,n2065);
    or g1160(n2431 ,n2360 ,n2064);
    or g1161(n2430 ,n2361 ,n2362);
    or g1162(n2429 ,n2001 ,n2333);
    or g1163(n2428 ,n2363 ,n2063);
    or g1164(n2427 ,n2364 ,n2093);
    or g1165(n2426 ,n2190 ,n2062);
    or g1166(n2425 ,n2188 ,n2189);
    or g1167(n2424 ,n2000 ,n2332);
    or g1168(n2423 ,n2187 ,n2061);
    or g1169(n2422 ,n2186 ,n2185);
    or g1170(n2421 ,n2184 ,n2060);
    or g1171(n2420 ,n2183 ,n2182);
    or g1172(n2419 ,n2181 ,n2059);
    or g1173(n2418 ,n2180 ,n2179);
    or g1174(n2417 ,n1850 ,n2325);
    or g1175(n2416 ,n2178 ,n2058);
    or g1176(n2415 ,n1926 ,n2176);
    or g1177(n2414 ,n1849 ,n2324);
    or g1178(n2413 ,n2175 ,n2057);
    or g1179(n2412 ,n1925 ,n2173);
    or g1180(n2411 ,n2172 ,n2056);
    or g1181(n2410 ,n2171 ,n2170);
    or g1182(n2409 ,n2169 ,n2055);
    or g1183(n2408 ,n1923 ,n2167);
    or g1184(n2407 ,n2166 ,n2054);
    or g1185(n2406 ,n1922 ,n2164);
    or g1186(n2405 ,n2163 ,n2053);
    or g1187(n2404 ,n1921 ,n2161);
    or g1188(n2403 ,n2160 ,n2052);
    or g1189(n2402 ,n1920 ,n2158);
    or g1190(n2401 ,n2157 ,n2050);
    or g1191(n2400 ,n2154 ,n2051);
    or g1192(n2399 ,n1919 ,n2155);
    or g1193(n2398 ,n1918 ,n2152);
    or g1194(n2397 ,n2151 ,n2150);
    or g1195(n2396 ,n1917 ,n2049);
    or g1196(n2395 ,n1983 ,n2121);
    or g1197(n2394 ,n2148 ,n2048);
    or g1198(n2393 ,n2147 ,n2146);
    or g1199(n2392 ,n2145 ,n2035);
    or g1200(n2391 ,n1915 ,n2143);
    or g1201(n2390 ,n2140 ,n2047);
    or g1202(n2389 ,n2139 ,n2141);
    or g1203(n2388 ,n2138 ,n2046);
    or g1204(n2387 ,n1913 ,n2136);
    or g1205(n2386 ,n2135 ,n2045);
    or g1206(n2385 ,n1912 ,n2133);
    or g1207(n2384 ,n1911 ,n2130);
    or g1208(n2383 ,n2101 ,n2320);
    or g1209(n2382 ,n2132 ,n2044);
    or g1210(n2381 ,n2128 ,n2043);
    or g1211(n2380 ,n1910 ,n2127);
    or g1212(n2379 ,n2124 ,n2042);
    or g1213(n2378 ,n1909 ,n2122);
    or g1214(n2377 ,n1907 ,n2117);
    or g1215(n2376 ,n2120 ,n2041);
    or g1216(n2375 ,n2116 ,n2040);
    or g1217(n2374 ,n1906 ,n2113);
    or g1218(n2373 ,n1905 ,n2112);
    or g1219(n2372 ,n2110 ,n2039);
    or g1220(n2371 ,n2109 ,n2038);
    or g1221(n2370 ,n2108 ,n2107);
    or g1222(n2369 ,n2106 ,n2037);
    or g1223(n2368 ,n1970 ,n2260);
    or g1224(n2367 ,n2103 ,n2104);
    or g1225(n2366 ,n2102 ,n2036);
    or g1226(n2497 ,n1847 ,n2193);
    nor g1227(n2365 ,n671 ,n529);
    nor g1228(n2364 ,n844 ,n526);
    nor g1229(n2363 ,n674 ,n530);
    nor g1230(n2362 ,n1306 ,n532);
    nor g1231(n2361 ,n595 ,n527);
    nor g1232(n2360 ,n647 ,n529);
    nor g1233(n2359 ,n858 ,n526);
    nor g1234(n2358 ,n1304 ,n533);
    nor g1235(n2357 ,n882 ,n530);
    nor g1236(n2356 ,n558 ,n532);
    nor g1237(n2355 ,n773 ,n527);
    nor g1238(n2354 ,n1261 ,n529);
    nor g1239(n2353 ,n729 ,n533);
    nor g1240(n2352 ,n1313 ,n526);
    nor g1241(n2351 ,n778 ,n530);
    nor g1242(n2350 ,n1269 ,n527);
    nor g1243(n2349 ,n667 ,n532);
    nor g1244(n2348 ,n586 ,n527);
    nor g1245(n2347 ,n701 ,n530);
    nor g1246(n2346 ,n665 ,n533);
    nor g1247(n2345 ,n685 ,n527);
    nor g1248(n2344 ,n744 ,n530);
    nor g1249(n2343 ,n893 ,n533);
    nor g1250(n2342 ,n731 ,n530);
    nor g1251(n2341 ,n676 ,n527);
    nor g1252(n2340 ,n888 ,n533);
    nor g1253(n2339 ,n712 ,n529);
    nor g1254(n2338 ,n1334 ,n526);
    nor g1255(n2337 ,n652 ,n530);
    or g1256(n2336 ,n1068 ,n1943);
    nor g1257(n2335 ,n1049 ,n1939);
    nor g1258(n2334 ,n1041 ,n1949);
    nor g1259(n2333 ,n1046 ,n1947);
    nor g1260(n2332 ,n1047 ,n1945);
    nor g1261(n2331 ,n980 ,n1934);
    nor g1262(n2330 ,n994 ,n1935);
    nor g1263(n2329 ,n1219 ,n1935);
    nor g1264(n2328 ,n1061 ,n1934);
    nor g1265(n2327 ,n1222 ,n1935);
    nor g1266(n2326 ,n1155 ,n1934);
    nor g1267(n2325 ,n1048 ,n1935);
    nor g1268(n2324 ,n1051 ,n1934);
    nor g1269(n2323 ,n881 ,n529);
    nor g1270(n2322 ,n624 ,n533);
    nor g1271(n2321 ,n797 ,n527);
    nor g1272(n2320 ,n649 ,n532);
    nor g1273(n2319 ,n763 ,n526);
    nor g1274(n2318 ,n896 ,n530);
    nor g1275(n2317 ,n784 ,n533);
    nor g1276(n2316 ,n861 ,n530);
    nor g1277(n2315 ,n732 ,n527);
    nor g1278(n2314 ,n1310 ,n532);
    nor g1279(n2313 ,n695 ,n529);
    nor g1280(n2312 ,n765 ,n527);
    nor g1281(n2311 ,n758 ,n533);
    nor g1282(n2310 ,n636 ,n530);
    nor g1283(n2309 ,n1335 ,n533);
    nor g1284(n2308 ,n842 ,n526);
    nor g1285(n2307 ,n786 ,n530);
    nor g1286(n2306 ,n909 ,n527);
    nor g1287(n2305 ,n576 ,n532);
    nor g1288(n2304 ,n852 ,n527);
    nor g1289(n2303 ,n603 ,n529);
    nor g1290(n2302 ,n1277 ,n533);
    nor g1291(n2301 ,n818 ,n529);
    nor g1292(n2300 ,n835 ,n526);
    nor g1293(n2299 ,n766 ,n533);
    nor g1294(n2298 ,n694 ,n530);
    nor g1295(n2297 ,n598 ,n526);
    nor g1296(n2296 ,n637 ,n532);
    nor g1297(n2295 ,n823 ,n530);
    nor g1298(n2294 ,n824 ,n527);
    nor g1299(n2293 ,n746 ,n532);
    nor g1300(n2292 ,n924 ,n530);
    nor g1301(n2291 ,n770 ,n527);
    nor g1302(n2290 ,n693 ,n533);
    nor g1303(n2289 ,n781 ,n527);
    nor g1304(n2288 ,n814 ,n530);
    nor g1305(n2287 ,n684 ,n533);
    nor g1306(n2286 ,n897 ,n530);
    nor g1307(n2285 ,n575 ,n530);
    nor g1308(n2284 ,n822 ,n533);
    nor g1309(n2283 ,n891 ,n527);
    nor g1310(n2282 ,n795 ,n530);
    nor g1311(n2281 ,n745 ,n533);
    nor g1312(n2280 ,n790 ,n527);
    nor g1313(n2279 ,n606 ,n529);
    nor g1314(n2278 ,n560 ,n527);
    nor g1315(n2277 ,n826 ,n527);
    nor g1316(n2276 ,n1295 ,n533);
    nor g1317(n2275 ,n1256 ,n530);
    nor g1318(n2274 ,n660 ,n526);
    nor g1319(n2273 ,n661 ,n533);
    nor g1320(n2272 ,n869 ,n533);
    nor g1321(n2271 ,n666 ,n529);
    nor g1322(n2270 ,n689 ,n532);
    nor g1323(n2269 ,n1298 ,n527);
    nor g1324(n2268 ,n1299 ,n526);
    nor g1325(n2267 ,n935 ,n526);
    nor g1326(n2266 ,n794 ,n533);
    nor g1327(n2265 ,n1337 ,n529);
    nor g1328(n2264 ,n752 ,n532);
    nor g1329(n2263 ,n585 ,n532);
    nor g1330(n2262 ,n646 ,n527);
    nor g1331(n2261 ,n1329 ,n530);
    nor g1332(n2260 ,n905 ,n529);
    nor g1333(n2259 ,n583 ,n526);
    nor g1334(n2258 ,n769 ,n533);
    nor g1335(n2257 ,n1274 ,n530);
    nor g1336(n2256 ,n865 ,n529);
    nor g1337(n2255 ,n722 ,n532);
    nor g1338(n2254 ,n1318 ,n527);
    nor g1339(n2253 ,n750 ,n533);
    nor g1340(n2252 ,n1262 ,n529);
    nor g1341(n2251 ,n747 ,n530);
    nor g1342(n2250 ,n937 ,n532);
    nor g1343(n2249 ,n1293 ,n526);
    nor g1344(n2248 ,n1278 ,n529);
    nor g1345(n2247 ,n880 ,n526);
    nor g1346(n2246 ,n1315 ,n532);
    nor g1347(n2245 ,n911 ,n530);
    nor g1348(n2244 ,n838 ,n527);
    nor g1349(n2243 ,n565 ,n533);
    nor g1350(n2242 ,n642 ,n530);
    nor g1351(n2241 ,n799 ,n532);
    nor g1352(n2240 ,n771 ,n526);
    nor g1353(n2239 ,n807 ,n530);
    nor g1354(n2238 ,n913 ,n533);
    nor g1355(n2237 ,n1280 ,n527);
    nor g1356(n2236 ,n625 ,n530);
    nor g1357(n2235 ,n662 ,n527);
    nor g1358(n2234 ,n885 ,n533);
    nor g1359(n2233 ,n1292 ,n530);
    nor g1360(n2232 ,n1294 ,n529);
    nor g1361(n2231 ,n1287 ,n533);
    nor g1362(n2230 ,n1325 ,n527);
    nor g1363(n2229 ,n622 ,n529);
    nor g1364(n2228 ,n559 ,n533);
    nor g1365(n2227 ,n1336 ,n527);
    nor g1366(n2226 ,n1290 ,n529);
    nor g1367(n2225 ,n830 ,n533);
    nor g1368(n2224 ,n821 ,n532);
    nor g1369(n2223 ,n902 ,n527);
    nor g1370(n2222 ,n1264 ,n532);
    nor g1371(n2221 ,n578 ,n530);
    nor g1372(n2220 ,n922 ,n532);
    nor g1373(n2219 ,n579 ,n533);
    nor g1374(n2218 ,n1296 ,n533);
    nor g1375(n2217 ,n857 ,n533);
    nor g1376(n2216 ,n658 ,n526);
    nor g1377(n2215 ,n677 ,n530);
    nor g1378(n2214 ,n1323 ,n526);
    nor g1379(n2213 ,n648 ,n526);
    nor g1380(n2212 ,n933 ,n530);
    nor g1381(n2211 ,n672 ,n527);
    nor g1382(n2210 ,n568 ,n530);
    nor g1383(n2209 ,n900 ,n527);
    nor g1384(n2208 ,n687 ,n533);
    nor g1385(n2207 ,n680 ,n527);
    nor g1386(n2206 ,n738 ,n529);
    nor g1387(n2205 ,n640 ,n530);
    nor g1388(n2204 ,n1270 ,n532);
    nor g1389(n2203 ,n557 ,n527);
    nor g1390(n2202 ,n916 ,n526);
    nor g1391(n2201 ,n686 ,n529);
    nor g1392(n2200 ,n607 ,n533);
    nor g1393(n2199 ,n690 ,n527);
    nor g1394(n2198 ,n847 ,n526);
    not g1395(n2192 ,n2193);
    nor g1396(n2191 ,n1091 ,n536);
    nor g1397(n2190 ,n884 ,n529);
    nor g1398(n2189 ,n829 ,n532);
    nor g1399(n2188 ,n679 ,n526);
    nor g1400(n2187 ,n706 ,n529);
    nor g1401(n2186 ,n760 ,n526);
    nor g1402(n2185 ,n644 ,n532);
    nor g1403(n2184 ,n1268 ,n530);
    nor g1404(n2183 ,n656 ,n527);
    nor g1405(n2182 ,n734 ,n532);
    nor g1406(n2181 ,n1308 ,n530);
    nor g1407(n2180 ,n655 ,n527);
    nor g1408(n2179 ,n643 ,n533);
    nor g1409(n2178 ,n1279 ,n526);
    nor g1410(n2177 ,n610 ,n529);
    nor g1411(n2176 ,n753 ,n533);
    nor g1412(n2175 ,n912 ,n530);
    nor g1413(n2174 ,n833 ,n527);
    nor g1414(n2173 ,n925 ,n532);
    nor g1415(n2172 ,n800 ,n529);
    nor g1416(n2171 ,n837 ,n526);
    nor g1417(n2170 ,n571 ,n533);
    nor g1418(n2169 ,n785 ,n527);
    nor g1419(n2168 ,n1285 ,n530);
    nor g1420(n2167 ,n1322 ,n532);
    nor g1421(n2166 ,n1301 ,n527);
    nor g1422(n2165 ,n872 ,n530);
    nor g1423(n2164 ,n668 ,n533);
    nor g1424(n2163 ,n1273 ,n527);
    nor g1425(n2162 ,n727 ,n530);
    nor g1426(n2161 ,n1260 ,n533);
    nor g1427(n2160 ,n612 ,n526);
    nor g1428(n2159 ,n860 ,n529);
    nor g1429(n2158 ,n867 ,n533);
    nor g1430(n2157 ,n711 ,n527);
    nor g1431(n2156 ,n601 ,n530);
    nor g1432(n2155 ,n779 ,n532);
    nor g1433(n2154 ,n589 ,n527);
    nor g1434(n2153 ,n718 ,n530);
    nor g1435(n2152 ,n802 ,n533);
    nor g1436(n2151 ,n638 ,n527);
    nor g1437(n2150 ,n599 ,n533);
    nor g1438(n2149 ,n593 ,n530);
    nor g1439(n2148 ,n650 ,n526);
    nor g1440(n2147 ,n1312 ,n529);
    nor g1441(n2146 ,n927 ,n533);
    nor g1442(n2145 ,n1324 ,n526);
    nor g1443(n2144 ,n926 ,n529);
    nor g1444(n2143 ,n1289 ,n532);
    nor g1445(n2142 ,n700 ,n532);
    nor g1446(n2141 ,n663 ,n533);
    nor g1447(n2140 ,n703 ,n530);
    nor g1448(n2139 ,n934 ,n527);
    nor g1449(n2138 ,n724 ,n529);
    nor g1450(n2137 ,n582 ,n526);
    nor g1451(n2136 ,n569 ,n532);
    nor g1452(n2135 ,n675 ,n527);
    nor g1453(n2134 ,n920 ,n530);
    nor g1454(n2133 ,n555 ,n533);
    nor g1455(n2132 ,n873 ,n527);
    nor g1456(n2131 ,n626 ,n530);
    nor g1457(n2130 ,n878 ,n533);
    nor g1458(n2129 ,n918 ,n533);
    nor g1459(n2128 ,n617 ,n527);
    nor g1460(n2127 ,n688 ,n532);
    nor g1461(n2126 ,n903 ,n530);
    nor g1462(n2125 ,n651 ,n529);
    nor g1463(n2124 ,n849 ,n526);
    nor g1464(n2123 ,n843 ,n529);
    nor g1465(n2122 ,n623 ,n532);
    nor g1466(n2121 ,n759 ,n526);
    nor g1467(n2120 ,n940 ,n527);
    nor g1468(n2119 ,n1326 ,n526);
    nor g1469(n2118 ,n1271 ,n530);
    nor g1470(n2117 ,n681 ,n533);
    nor g1471(n2116 ,n836 ,n529);
    nor g1472(n2115 ,n910 ,n532);
    nor g1473(n2114 ,n1266 ,n527);
    nor g1474(n2113 ,n631 ,n533);
    nor g1475(n2112 ,n692 ,n530);
    nor g1476(n2111 ,n936 ,n533);
    nor g1477(n2110 ,n923 ,n527);
    nor g1478(n2109 ,n580 ,n530);
    nor g1479(n2108 ,n554 ,n526);
    nor g1480(n2107 ,n1319 ,n532);
    nor g1481(n2106 ,n720 ,n529);
    nor g1482(n2105 ,n741 ,n530);
    nor g1483(n2104 ,n813 ,n533);
    nor g1484(n2103 ,n669 ,n527);
    nor g1485(n2102 ,n682 ,n530);
    nor g1486(n2101 ,n615 ,n527);
    nor g1487(n2100 ,n1144 ,n1933);
    nor g1488(n2099 ,n1116 ,n535);
    nor g1489(n2098 ,n1234 ,n536);
    nor g1490(n2097 ,n1180 ,n1933);
    nor g1491(n2096 ,n1141 ,n1933);
    nor g1492(n2095 ,n1151 ,n536);
    nor g1493(n2094 ,n1106 ,n1933);
    nor g1494(n2093 ,n930 ,n533);
    nor g1495(n2092 ,n1236 ,n1933);
    nor g1496(n2091 ,n1136 ,n1933);
    nor g1497(n2090 ,n1145 ,n535);
    nor g1498(n2089 ,n1228 ,n536);
    nor g1499(n2088 ,n1148 ,n1933);
    nor g1500(n2087 ,n1247 ,n1933);
    nor g1501(n2086 ,n1075 ,n1933);
    nor g1502(n2085 ,n1134 ,n1933);
    nor g1503(n2084 ,n1166 ,n1933);
    nor g1504(n2083 ,n1250 ,n536);
    nor g1505(n2082 ,n1193 ,n1933);
    nor g1506(n2081 ,n1084 ,n536);
    nor g1507(n2080 ,n1162 ,n535);
    nor g1508(n2079 ,n1213 ,n536);
    nor g1509(n2078 ,n1253 ,n1933);
    nor g1510(n2077 ,n1200 ,n535);
    nor g1511(n2076 ,n1238 ,n536);
    nor g1512(n2075 ,n1130 ,n1933);
    nor g1513(n2074 ,n1055 ,n1933);
    nor g1514(n2073 ,n1097 ,n1933);
    nor g1515(n2072 ,n1242 ,n535);
    nor g1516(n2071 ,n1188 ,n536);
    nor g1517(n2070 ,n1183 ,n536);
    nor g1518(n2069 ,n1172 ,n536);
    nor g1519(n2068 ,n1177 ,n536);
    nor g1520(n2067 ,n1125 ,n1933);
    nor g1521(n2066 ,n1252 ,n1933);
    nor g1522(n2065 ,n1199 ,n536);
    nor g1523(n2064 ,n1159 ,n536);
    nor g1524(n2063 ,n1154 ,n1933);
    nor g1525(n2062 ,n1206 ,n1933);
    nor g1526(n2061 ,n1085 ,n535);
    nor g1527(n2060 ,n1099 ,n1933);
    nor g1528(n2059 ,n1137 ,n1933);
    nor g1529(n2058 ,n1131 ,n536);
    nor g1530(n2057 ,n1117 ,n536);
    nor g1531(n2056 ,n1122 ,n536);
    nor g1532(n2055 ,n1089 ,n1933);
    nor g1533(n2054 ,n1101 ,n1933);
    nor g1534(n2053 ,n1109 ,n1933);
    nor g1535(n2052 ,n1118 ,n536);
    nor g1536(n2051 ,n1158 ,n1933);
    nor g1537(n2050 ,n1152 ,n1933);
    nor g1538(n2049 ,n1027 ,n535);
    nor g1539(n2048 ,n1191 ,n535);
    nor g1540(n2047 ,n1233 ,n1933);
    nor g1541(n2046 ,n1086 ,n1933);
    nor g1542(n2045 ,n1080 ,n535);
    nor g1543(n2044 ,n1081 ,n535);
    nor g1544(n2043 ,n1164 ,n535);
    nor g1545(n2042 ,n1225 ,n536);
    nor g1546(n2041 ,n1056 ,n535);
    nor g1547(n2040 ,n1108 ,n1933);
    nor g1548(n2039 ,n1229 ,n536);
    nor g1549(n2038 ,n1104 ,n536);
    nor g1550(n2037 ,n1167 ,n536);
    nor g1551(n2036 ,n1209 ,n536);
    nor g1552(n2035 ,n964 ,n535);
    or g1553(n2034 ,n1541 ,n1898);
    or g1554(n2033 ,n1542 ,n1897);
    or g1555(n2032 ,n1499 ,n1896);
    or g1556(n2031 ,n1476 ,n1894);
    or g1557(n2030 ,n1485 ,n1893);
    or g1558(n2029 ,n1500 ,n1891);
    or g1559(n2028 ,n1510 ,n1890);
    or g1560(n2027 ,n1501 ,n1889);
    or g1561(n2026 ,n1841 ,n528);
    nor g1562(n2025 ,n951 ,n536);
    nor g1563(n2024 ,n950 ,n535);
    nor g1564(n2023 ,n947 ,n536);
    nor g1565(n2022 ,n952 ,n535);
    nor g1566(n2021 ,n958 ,n536);
    nor g1567(n2020 ,n957 ,n536);
    nor g1568(n2019 ,n959 ,n535);
    nor g1569(n2018 ,n954 ,n536);
    nor g1570(n2017 ,n960 ,n535);
    nor g1571(n2016 ,n955 ,n536);
    nor g1572(n2015 ,n956 ,n536);
    nor g1573(n2014 ,n948 ,n535);
    nor g1574(n2013 ,n944 ,n1933);
    nor g1575(n2012 ,n946 ,n536);
    nor g1576(n2011 ,n949 ,n535);
    nor g1577(n2010 ,n953 ,n536);
    or g1578(n2009 ,n1840 ,n531);
    nor g1579(n2008 ,n1545 ,n1883);
    or g1580(n2007 ,n1824 ,n534);
    nor g1581(n2006 ,n1550 ,n1885);
    nor g1582(n2005 ,n538 ,n1900);
    nor g1583(n2004 ,n1549 ,n1942);
    nor g1584(n2003 ,n542 ,n1938);
    nor g1585(n2002 ,n542 ,n1948);
    nor g1586(n2001 ,n540 ,n1946);
    nor g1587(n2000 ,n538 ,n1944);
    or g1588(n2197 ,n544 ,n1884);
    or g1589(n2196 ,n537 ,n1937);
    or g1590(n2195 ,n544 ,n1936);
    or g1591(n2194 ,n1848 ,n1940);
    nor g1592(n2193 ,n1661 ,n1941);
    nor g1593(n1999 ,n715 ,n523);
    nor g1594(n1998 ,n904 ,n524);
    nor g1595(n1997 ,n748 ,n523);
    nor g1596(n1996 ,n801 ,n524);
    nor g1597(n1995 ,n780 ,n523);
    nor g1598(n1994 ,n764 ,n524);
    nor g1599(n1993 ,n831 ,n524);
    nor g1600(n1992 ,n832 ,n524);
    nor g1601(n1991 ,n653 ,n524);
    nor g1602(n1990 ,n1282 ,n523);
    nor g1603(n1989 ,n673 ,n524);
    nor g1604(n1988 ,n1297 ,n523);
    nor g1605(n1987 ,n616 ,n524);
    nor g1606(n1986 ,n782 ,n524);
    nor g1607(n1985 ,n768 ,n523);
    nor g1608(n1984 ,n942 ,n524);
    nor g1609(n1983 ,n1328 ,n524);
    nor g1610(n1982 ,n1265 ,n523);
    nor g1611(n1981 ,n719 ,n523);
    nor g1612(n1980 ,n762 ,n524);
    nor g1613(n1979 ,n819 ,n524);
    nor g1614(n1978 ,n761 ,n524);
    nor g1615(n1977 ,n917 ,n524);
    nor g1616(n1976 ,n811 ,n524);
    nor g1617(n1975 ,n1283 ,n524);
    nor g1618(n1974 ,n757 ,n524);
    nor g1619(n1973 ,n899 ,n523);
    nor g1620(n1972 ,n941 ,n524);
    nor g1621(n1971 ,n572 ,n523);
    nor g1622(n1970 ,n562 ,n523);
    nor g1623(n1969 ,n594 ,n524);
    nor g1624(n1968 ,n654 ,n523);
    nor g1625(n1967 ,n573 ,n524);
    nor g1626(n1966 ,n928 ,n523);
    nor g1627(n1965 ,n696 ,n523);
    nor g1628(n1964 ,n848 ,n524);
    nor g1629(n1963 ,n635 ,n523);
    nor g1630(n1962 ,n919 ,n524);
    nor g1631(n1961 ,n870 ,n524);
    nor g1632(n1960 ,n755 ,n524);
    nor g1633(n1959 ,n590 ,n524);
    nor g1634(n1958 ,n641 ,n524);
    nor g1635(n1957 ,n707 ,n523);
    nor g1636(n1956 ,n1330 ,n523);
    nor g1637(n1955 ,n1257 ,n523);
    nor g1638(n1954 ,n609 ,n524);
    nor g1639(n1953 ,n709 ,n524);
    nor g1640(n1952 ,n627 ,n524);
    nor g1641(n1951 ,n728 ,n524);
    nor g1642(n1950 ,n621 ,n523);
    not g1643(n1949 ,n1948);
    not g1644(n1947 ,n1946);
    not g1645(n1945 ,n1944);
    not g1646(n1943 ,n1942);
    not g1647(n1941 ,n1940);
    not g1648(n1939 ,n1938);
    not g1649(n1933 ,n1932);
    not g1650(n536 ,n1932);
    not g1651(n535 ,n1932);
    not g1652(n533 ,n534);
    not g1653(n532 ,n534);
    not g1654(n530 ,n531);
    not g1655(n529 ,n531);
    not g1656(n527 ,n528);
    not g1657(n526 ,n528);
    nor g1658(n1931 ,n538 ,n1757);
    nor g1659(n1930 ,n1320 ,n524);
    nor g1660(n1929 ,n614 ,n523);
    nor g1661(n1928 ,n1281 ,n523);
    nor g1662(n1927 ,n553 ,n523);
    nor g1663(n1926 ,n886 ,n524);
    nor g1664(n1925 ,n772 ,n524);
    nor g1665(n1924 ,n1317 ,n523);
    nor g1666(n1923 ,n1276 ,n524);
    nor g1667(n1922 ,n751 ,n523);
    nor g1668(n1921 ,n670 ,n524);
    nor g1669(n1920 ,n570 ,n524);
    nor g1670(n1919 ,n739 ,n524);
    nor g1671(n1918 ,n840 ,n523);
    nor g1672(n1917 ,n789 ,n524);
    nor g1673(n1916 ,n775 ,n524);
    nor g1674(n1915 ,n733 ,n524);
    nor g1675(n1914 ,n906 ,n523);
    nor g1676(n1913 ,n1316 ,n523);
    nor g1677(n1912 ,n804 ,n524);
    nor g1678(n1911 ,n875 ,n523);
    nor g1679(n1910 ,n591 ,n524);
    nor g1680(n1909 ,n736 ,n524);
    nor g1681(n1908 ,n639 ,n524);
    nor g1682(n1907 ,n841 ,n523);
    nor g1683(n1906 ,n908 ,n523);
    nor g1684(n1905 ,n619 ,n524);
    nor g1685(n1904 ,n816 ,n523);
    nor g1686(n1903 ,n915 ,n524);
    nor g1687(n1902 ,n1291 ,n524);
    nor g1688(n1901 ,n629 ,n523);
    nor g1689(n1900 ,n1807 ,n1852);
    or g1690(n1899 ,n1535 ,n1839);
    or g1691(n1898 ,n1544 ,n1821);
    or g1692(n1897 ,n1489 ,n1820);
    or g1693(n1896 ,n1523 ,n1837);
    or g1694(n1895 ,n1520 ,n1836);
    or g1695(n1894 ,n1565 ,n1818);
    or g1696(n1893 ,n1492 ,n1835);
    or g1697(n1892 ,n1498 ,n1834);
    or g1698(n1891 ,n1481 ,n1816);
    or g1699(n1890 ,n1509 ,n1815);
    or g1700(n1889 ,n1504 ,n1813);
    or g1701(n1888 ,n1507 ,n1833);
    nor g1702(n1887 ,n1263 ,n524);
    or g1703(n1886 ,n1842 ,n525);
    nor g1704(n1885 ,n1851 ,n1853);
    or g1705(n1884 ,n1571 ,n1803);
    or g1706(n1883 ,n1566 ,n1852);
    nor g1707(n1882 ,n538 ,n1812);
    nor g1708(n1881 ,n540 ,n1755);
    nor g1709(n1880 ,n537 ,n1811);
    nor g1710(n1879 ,n539 ,n1747);
    nor g1711(n1878 ,n538 ,n1750);
    nor g1712(n1877 ,n542 ,n1752);
    nor g1713(n1876 ,n539 ,n1830);
    nor g1714(n1875 ,n539 ,n1769);
    nor g1715(n1874 ,n541 ,n1832);
    nor g1716(n1873 ,n538 ,n1844);
    nor g1717(n1872 ,n539 ,n1846);
    nor g1718(n1871 ,n543 ,n1774);
    nor g1719(n1870 ,n541 ,n1804);
    nor g1720(n1869 ,n541 ,n1845);
    nor g1721(n1868 ,n541 ,n1801);
    nor g1722(n1867 ,n543 ,n1823);
    nor g1723(n1866 ,n539 ,n1756);
    nor g1724(n1865 ,n537 ,n1766);
    nor g1725(n1864 ,n539 ,n1765);
    nor g1726(n1863 ,n540 ,n1764);
    nor g1727(n1862 ,n543 ,n1763);
    nor g1728(n1861 ,n540 ,n1762);
    nor g1729(n1860 ,n540 ,n1761);
    nor g1730(n1859 ,n542 ,n1760);
    nor g1731(n1858 ,n542 ,n1759);
    nor g1732(n1857 ,n540 ,n1758);
    nor g1733(n1856 ,n542 ,n1822);
    nor g1734(n1855 ,n834 ,n524);
    nor g1735(n1948 ,n1526 ,n1827);
    nor g1736(n1946 ,n1527 ,n1826);
    nor g1737(n1944 ,n1529 ,n1825);
    nor g1738(n1942 ,n1573 ,n1847);
    nor g1739(n1940 ,n44[0] ,n1803);
    nor g1740(n1938 ,n1525 ,n1828);
    nor g1741(n1937 ,n1406 ,n1831);
    nor g1742(n1936 ,n1400 ,n1829);
    or g1743(n1935 ,n544 ,n1850);
    or g1744(n1934 ,n544 ,n1849);
    or g1745(n1932 ,n1655 ,n1843);
    nor g1746(n534 ,n1746 ,n1810);
    nor g1747(n531 ,n1572 ,n1809);
    nor g1748(n528 ,n3261 ,n1808);
    not g1749(n1854 ,n1853);
    not g1750(n1852 ,n1851);
    not g1751(n1848 ,n1847);
    not g1752(n524 ,n525);
    not g1753(n523 ,n525);
    nor g1754(n1846 ,n1624 ,n1640);
    nor g1755(n1845 ,n1629 ,n1638);
    nor g1756(n1844 ,n1622 ,n1642);
    nor g1757(n1843 ,n551 ,n1746);
    nor g1758(n1842 ,n996 ,n1656);
    nor g1759(n1841 ,n967 ,n1656);
    nor g1760(n1840 ,n962 ,n1656);
    or g1761(n1839 ,n1537 ,n1606);
    or g1762(n1838 ,n1547 ,n1605);
    or g1763(n1837 ,n1503 ,n1604);
    or g1764(n1836 ,n1519 ,n1603);
    or g1765(n1835 ,n1475 ,n1602);
    or g1766(n1834 ,n1512 ,n1601);
    or g1767(n1833 ,n1478 ,n1600);
    nor g1768(n1832 ,n1618 ,n1637);
    or g1769(n1831 ,n1402 ,n1657);
    nor g1770(n1830 ,n1613 ,n1643);
    or g1771(n1829 ,n1401 ,n1657);
    nor g1772(n1828 ,n1568 ,n1659);
    nor g1773(n1827 ,n1574 ,n1659);
    nor g1774(n1826 ,n1568 ,n1658);
    nor g1775(n1825 ,n1574 ,n1658);
    nor g1776(n1824 ,n943 ,n1656);
    nor g1777(n1823 ,n1614 ,n1645);
    nor g1778(n1822 ,n1631 ,n1653);
    or g1779(n1821 ,n1393 ,n1593);
    or g1780(n1820 ,n1368 ,n1592);
    or g1781(n1819 ,n1357 ,n1591);
    or g1782(n1818 ,n1408 ,n1590);
    or g1783(n1817 ,n1362 ,n1589);
    or g1784(n1816 ,n1373 ,n1588);
    or g1785(n1815 ,n1448 ,n1587);
    or g1786(n1814 ,n1384 ,n1586);
    or g1787(n1813 ,n1377 ,n1585);
    nor g1788(n1812 ,n1610 ,n1647);
    nor g1789(n1811 ,n1611 ,n1636);
    or g1790(n1810 ,n3259 ,n1655);
    or g1791(n1809 ,n3260 ,n1655);
    or g1792(n1808 ,n1465 ,n1655);
    or g1793(n1807 ,n43[2] ,n1597);
    or g1794(n1806 ,n1726 ,n1744);
    or g1795(n1805 ,n1743 ,n1728);
    nor g1796(n1804 ,n1625 ,n1639);
    nor g1797(n1853 ,n1654 ,n1660);
    nor g1798(n1851 ,n1528 ,n1660);
    nor g1799(n1850 ,n1657 ,n1562);
    nor g1800(n1849 ,n1657 ,n1565);
    nor g1801(n1847 ,n44[1] ,n1661);
    nor g1802(n525 ,n1464 ,n1655);
    or g1803(n1802 ,n1708 ,n1732);
    nor g1804(n1801 ,n1621 ,n1641);
    or g1805(n1800 ,n1740 ,n1583);
    or g1806(n1799 ,n1669 ,n1672);
    or g1807(n1798 ,n1739 ,n1688);
    or g1808(n1797 ,n1691 ,n1689);
    or g1809(n1796 ,n1690 ,n1692);
    or g1810(n1795 ,n1694 ,n1693);
    or g1811(n1794 ,n1738 ,n1698);
    or g1812(n1793 ,n1737 ,n1695);
    or g1813(n1792 ,n1736 ,n1696);
    or g1814(n1791 ,n1697 ,n1699);
    or g1815(n1790 ,n1735 ,n1594);
    or g1816(n1789 ,n1731 ,n1741);
    or g1817(n1788 ,n1727 ,n1710);
    or g1818(n1787 ,n1724 ,n1723);
    or g1819(n1786 ,n1745 ,n1722);
    or g1820(n1785 ,n1700 ,n1702);
    or g1821(n1784 ,n1712 ,n1711);
    or g1822(n1783 ,n1680 ,n1671);
    or g1823(n1782 ,n1670 ,n1719);
    or g1824(n1781 ,n1687 ,n1595);
    or g1825(n1780 ,n1717 ,n1674);
    or g1826(n1779 ,n1715 ,n1682);
    or g1827(n1778 ,n1714 ,n1681);
    or g1828(n1777 ,n1730 ,n1742);
    or g1829(n1776 ,n1707 ,n1709);
    or g1830(n1775 ,n1733 ,n1704);
    nor g1831(n1774 ,n1632 ,n1649);
    or g1832(n1773 ,n1705 ,n1721);
    or g1833(n1772 ,n1734 ,n1701);
    or g1834(n1771 ,n1725 ,n1596);
    or g1835(n1770 ,n1729 ,n1683);
    nor g1836(n1769 ,n1630 ,n1650);
    or g1837(n1768 ,n1686 ,n1685);
    or g1838(n1767 ,n1713 ,n1684);
    nor g1839(n1766 ,n1617 ,n1667);
    nor g1840(n1765 ,n1619 ,n1666);
    nor g1841(n1764 ,n1616 ,n1665);
    nor g1842(n1763 ,n1628 ,n1664);
    nor g1843(n1762 ,n1620 ,n1663);
    nor g1844(n1761 ,n1623 ,n1662);
    nor g1845(n1760 ,n1615 ,n1703);
    nor g1846(n1759 ,n1627 ,n1607);
    nor g1847(n1758 ,n1633 ,n1668);
    nor g1848(n1757 ,n1634 ,n1652);
    nor g1849(n1756 ,n1635 ,n1651);
    xnor g1850(n1755 ,n1550 ,n34[0]);
    or g1851(n1754 ,n1676 ,n1677);
    or g1852(n1753 ,n1716 ,n1675);
    nor g1853(n1752 ,n1626 ,n1644);
    or g1854(n1751 ,n1679 ,n1678);
    nor g1855(n1750 ,n1612 ,n1646);
    or g1856(n1749 ,n1718 ,n1673);
    or g1857(n1748 ,n1706 ,n1720);
    nor g1858(n1747 ,n1609 ,n1648);
    nor g1859(n1803 ,n1608 ,n1584);
    nor g1860(n1745 ,n1243 ,n1559);
    nor g1861(n1744 ,n791 ,n1555);
    nor g1862(n1743 ,n1077 ,n1558);
    nor g1863(n1742 ,n754 ,n1555);
    nor g1864(n1741 ,n749 ,n1555);
    nor g1865(n1740 ,n1042 ,n1553);
    nor g1866(n1739 ,n1170 ,n1553);
    nor g1867(n1738 ,n1083 ,n1553);
    nor g1868(n1737 ,n1244 ,n1553);
    nor g1869(n1736 ,n1224 ,n1553);
    nor g1870(n1735 ,n1045 ,n1558);
    nor g1871(n1734 ,n1063 ,n1558);
    nor g1872(n1733 ,n1067 ,n1558);
    nor g1873(n1732 ,n699 ,n1555);
    nor g1874(n1731 ,n1216 ,n1558);
    nor g1875(n1730 ,n1140 ,n1558);
    nor g1876(n1729 ,n1093 ,n1558);
    nor g1877(n1728 ,n1284 ,n1555);
    nor g1878(n1727 ,n1053 ,n1558);
    nor g1879(n1726 ,n1054 ,n1558);
    nor g1880(n1725 ,n1050 ,n1559);
    nor g1881(n1724 ,n1198 ,n1559);
    nor g1882(n1723 ,n932 ,n1554);
    nor g1883(n1722 ,n898 ,n1554);
    nor g1884(n1721 ,n1286 ,n1554);
    nor g1885(n1720 ,n1327 ,n1554);
    nor g1886(n1719 ,n713 ,n1554);
    nor g1887(n1718 ,n1059 ,n1557);
    nor g1888(n1717 ,n1112 ,n1557);
    nor g1889(n1716 ,n1147 ,n1557);
    nor g1890(n1715 ,n1255 ,n1557);
    nor g1891(n1714 ,n1254 ,n1557);
    nor g1892(n1713 ,n1087 ,n1557);
    nor g1893(n1712 ,n1098 ,n1559);
    nor g1894(n1711 ,n777 ,n1554);
    nor g1895(n1710 ,n806 ,n1555);
    nor g1896(n1709 ,n632 ,n1554);
    nor g1897(n1708 ,n1119 ,n1558);
    nor g1898(n1707 ,n1062 ,n1559);
    nor g1899(n1706 ,n1161 ,n1559);
    nor g1900(n1705 ,n1218 ,n1559);
    nor g1901(n1704 ,n743 ,n1555);
    nor g1902(n1703 ,n1046 ,n1551);
    nor g1903(n1702 ,n1311 ,n1554);
    nor g1904(n1701 ,n611 ,n1555);
    nor g1905(n1700 ,n1196 ,n1559);
    nor g1906(n1699 ,n1305 ,n1556);
    nor g1907(n1698 ,n921 ,n1556);
    nor g1908(n1697 ,n1202 ,n1553);
    nor g1909(n1696 ,n783 ,n1556);
    nor g1910(n1695 ,n820 ,n1556);
    nor g1911(n1694 ,n1115 ,n1553);
    nor g1912(n1693 ,n810 ,n1556);
    nor g1913(n1692 ,n698 ,n1556);
    nor g1914(n1691 ,n1070 ,n1553);
    nor g1915(n1690 ,n1208 ,n1553);
    nor g1916(n1689 ,n726 ,n1556);
    nor g1917(n1688 ,n756 ,n1556);
    nor g1918(n1687 ,n1043 ,n1557);
    nor g1919(n1686 ,n1124 ,n1557);
    nor g1920(n1685 ,n710 ,n1560);
    nor g1921(n1684 ,n605 ,n1560);
    nor g1922(n1683 ,n890 ,n1555);
    nor g1923(n1682 ,n883 ,n1560);
    nor g1924(n1681 ,n853 ,n1560);
    nor g1925(n1680 ,n1078 ,n1559);
    nor g1926(n1679 ,n1156 ,n1557);
    nor g1927(n1678 ,n628 ,n1560);
    nor g1928(n1677 ,n592 ,n1560);
    nor g1929(n1676 ,n1223 ,n1557);
    nor g1930(n1675 ,n815 ,n1560);
    nor g1931(n1674 ,n740 ,n1560);
    nor g1932(n1673 ,n702 ,n1560);
    nor g1933(n1672 ,n1332 ,n1556);
    nor g1934(n1671 ,n907 ,n1554);
    nor g1935(n1670 ,n1146 ,n1559);
    nor g1936(n1669 ,n1102 ,n1553);
    nor g1937(n1668 ,n1044 ,n1551);
    nor g1938(n1667 ,n1037 ,n1551);
    nor g1939(n1666 ,n1036 ,n1551);
    nor g1940(n1665 ,n1038 ,n1551);
    nor g1941(n1664 ,n1040 ,n1551);
    nor g1942(n1663 ,n1049 ,n1551);
    nor g1943(n1662 ,n1041 ,n1551);
    or g1944(n1746 ,n550 ,n1572);
    not g1945(n1655 ,n1656);
    nor g1946(n1654 ,n1403 ,n1570);
    nor g1947(n1653 ,n1048 ,n1551);
    nor g1948(n1652 ,n1051 ,n1551);
    nor g1949(n1651 ,n1039 ,n1551);
    nor g1950(n1650 ,n657 ,n1549);
    nor g1951(n1649 ,n618 ,n1549);
    nor g1952(n1648 ,n1331 ,n1549);
    nor g1953(n1647 ,n602 ,n1549);
    nor g1954(n1646 ,n1321 ,n1549);
    nor g1955(n1645 ,n1314 ,n1549);
    nor g1956(n1644 ,n604 ,n1549);
    nor g1957(n1643 ,n854 ,n1549);
    nor g1958(n1642 ,n767 ,n1549);
    nor g1959(n1641 ,n876 ,n1549);
    nor g1960(n1640 ,n735 ,n1549);
    nor g1961(n1639 ,n863 ,n1549);
    nor g1962(n1638 ,n581 ,n1549);
    nor g1963(n1637 ,n659 ,n1549);
    nor g1964(n1636 ,n788 ,n1549);
    nor g1965(n1635 ,n1231 ,n1552);
    nor g1966(n1634 ,n1195 ,n1552);
    nor g1967(n1633 ,n1092 ,n1552);
    nor g1968(n1632 ,n1160 ,n1550);
    nor g1969(n1631 ,n1071 ,n1552);
    nor g1970(n1630 ,n1203 ,n1550);
    nor g1971(n1629 ,n1127 ,n1550);
    nor g1972(n1628 ,n1230 ,n1552);
    nor g1973(n1627 ,n1227 ,n1552);
    nor g1974(n1626 ,n1194 ,n1550);
    nor g1975(n1625 ,n1153 ,n1550);
    nor g1976(n1624 ,n1139 ,n1550);
    nor g1977(n1623 ,n1176 ,n1552);
    nor g1978(n1622 ,n1121 ,n1550);
    nor g1979(n1621 ,n1129 ,n1550);
    nor g1980(n1620 ,n1217 ,n1552);
    nor g1981(n1619 ,n1174 ,n1552);
    nor g1982(n1618 ,n1204 ,n1550);
    nor g1983(n1617 ,n1142 ,n1552);
    nor g1984(n1616 ,n1226 ,n1552);
    nor g1985(n1615 ,n1123 ,n1552);
    nor g1986(n1614 ,n1192 ,n1550);
    nor g1987(n1613 ,n1207 ,n1550);
    nor g1988(n1612 ,n1186 ,n1550);
    nor g1989(n1611 ,n1212 ,n1550);
    nor g1990(n1610 ,n1179 ,n1550);
    nor g1991(n1609 ,n1173 ,n1550);
    nor g1992(n1608 ,n962 ,n1513);
    nor g1993(n1607 ,n1047 ,n1551);
    or g1994(n1606 ,n1538 ,n1539);
    or g1995(n1605 ,n1490 ,n1563);
    or g1996(n1604 ,n1522 ,n1521);
    or g1997(n1603 ,n1518 ,n1517);
    or g1998(n1602 ,n1515 ,n1514);
    or g1999(n1601 ,n1524 ,n1482);
    or g2000(n1600 ,n1506 ,n1505);
    nor g2001(n1599 ,n1561 ,n1564);
    nor g2002(n1598 ,n1561 ,n1563);
    nor g2003(n1597 ,n43[0] ,n1540);
    nor g2004(n1596 ,n48[0] ,n1554);
    nor g2005(n1595 ,n49[0] ,n1560);
    nor g2006(n1594 ,n47[0] ,n1555);
    or g2007(n1593 ,n1414 ,n1546);
    or g2008(n1592 ,n1429 ,n1491);
    or g2009(n1591 ,n1432 ,n1487);
    or g2010(n1590 ,n1370 ,n1516);
    or g2011(n1589 ,n1425 ,n1483);
    or g2012(n1588 ,n1462 ,n1564);
    or g2013(n1587 ,n1440 ,n1508);
    or g2014(n1586 ,n1417 ,n1562);
    or g2015(n1585 ,n1379 ,n1502);
    nor g2016(n1584 ,n1348 ,n1493);
    nor g2017(n1583 ,n46[0] ,n1556);
    nor g2018(n1582 ,n537 ,n1532);
    nor g2019(n1581 ,n543 ,n1495);
    nor g2020(n1580 ,n541 ,n1494);
    nor g2021(n1579 ,n541 ,n1496);
    nor g2022(n1578 ,n541 ,n1497);
    nor g2023(n1577 ,n538 ,n1533);
    nor g2024(n1576 ,n538 ,n1536);
    nor g2025(n1575 ,n542 ,n1531);
    or g2026(n1661 ,n544 ,n1549);
    or g2027(n1660 ,n1530 ,n1534);
    or g2028(n1659 ,n1400 ,n1569);
    or g2029(n1658 ,n1402 ,n1569);
    or g2030(n1657 ,n537 ,n1561);
    nor g2031(n1656 ,n542 ,n1567);
    not g2032(n1571 ,n1570);
    not g2033(n1567 ,n1566);
    not g2034(n1551 ,n1552);
    not g2035(n1549 ,n1550);
    or g2036(n1548 ,n1439 ,n1391);
    or g2037(n1547 ,n1392 ,n1351);
    or g2038(n1546 ,n1441 ,n1365);
    nor g2039(n1545 ,n961 ,n1404);
    or g2040(n1544 ,n1454 ,n1455);
    or g2041(n1543 ,n1438 ,n1361);
    or g2042(n1542 ,n1356 ,n1350);
    or g2043(n1541 ,n1442 ,n1416);
    nor g2044(n1540 ,n1342 ,n1345);
    or g2045(n1539 ,n1446 ,n1388);
    or g2046(n1538 ,n1443 ,n1380);
    or g2047(n1537 ,n1444 ,n1383);
    nor g2048(n1536 ,n1347 ,n1343);
    or g2049(n1535 ,n1445 ,n1395);
    or g2050(n1534 ,n1469 ,n1467);
    nor g2051(n1533 ,n1339 ,n1346);
    nor g2052(n1532 ,n1367 ,n1340);
    nor g2053(n1531 ,n1398 ,n1341);
    or g2054(n1530 ,n1466 ,n1468);
    or g2055(n1529 ,n544 ,n1467);
    nor g2056(n1528 ,n43[0] ,n1463);
    or g2057(n1527 ,n544 ,n1468);
    or g2058(n1526 ,n537 ,n1469);
    or g2059(n1525 ,n537 ,n1466);
    or g2060(n1574 ,n943 ,n1473);
    nor g2061(n1573 ,n43[2] ,n1404);
    or g2062(n1572 ,n552 ,n1465);
    nor g2063(n1570 ,n1457 ,n1463);
    or g2064(n1569 ,n1460 ,n1463);
    or g2065(n1568 ,n38[0] ,n1473);
    nor g2066(n1566 ,n43[2] ,n1405);
    or g2067(n1565 ,n1402 ,n1401);
    or g2068(n1564 ,n1419 ,n1401);
    or g2069(n1563 ,n1366 ,n1400);
    or g2070(n1562 ,n1406 ,n1400);
    or g2071(n1561 ,n961 ,n1405);
    or g2072(n1560 ,n3386 ,n1471);
    or g2073(n1559 ,n545 ,n1474);
    or g2074(n1558 ,n546 ,n1472);
    or g2075(n1557 ,n547 ,n1471);
    or g2076(n1556 ,n3383 ,n1470);
    or g2077(n1555 ,n3384 ,n1472);
    or g2078(n1554 ,n3385 ,n1474);
    or g2079(n1553 ,n548 ,n1470);
    nor g2080(n1552 ,n961 ,n1415);
    nor g2081(n1550 ,n945 ,n1463);
    or g2082(n1524 ,n1427 ,n1378);
    or g2083(n1523 ,n1461 ,n1355);
    or g2084(n1522 ,n1412 ,n1413);
    or g2085(n1521 ,n1435 ,n1375);
    or g2086(n1520 ,n1449 ,n1450);
    or g2087(n1519 ,n1411 ,n1410);
    or g2088(n1518 ,n1352 ,n1389);
    or g2089(n1517 ,n1385 ,n1354);
    or g2090(n1516 ,n1369 ,n1371);
    or g2091(n1515 ,n1387 ,n1399);
    or g2092(n1514 ,n1407 ,n1372);
    nor g2093(n1513 ,n1456 ,n1434);
    or g2094(n1512 ,n1430 ,n1364);
    or g2095(n1511 ,n1420 ,n1381);
    or g2096(n1510 ,n1421 ,n1396);
    or g2097(n1509 ,n1426 ,n1436);
    or g2098(n1508 ,n1394 ,n1360);
    or g2099(n1507 ,n1363 ,n1359);
    or g2100(n1506 ,n1428 ,n1424);
    or g2101(n1505 ,n1423 ,n1376);
    or g2102(n1504 ,n1458 ,n1422);
    or g2103(n1503 ,n1447 ,n1390);
    or g2104(n1502 ,n1382 ,n1374);
    or g2105(n1501 ,n1418 ,n1358);
    or g2106(n1500 ,n1459 ,n1386);
    or g2107(n1499 ,n1437 ,n1353);
    or g2108(n1498 ,n1409 ,n1431);
    nor g2109(n1497 ,n39[3] ,n1467);
    nor g2110(n1496 ,n39[2] ,n1468);
    nor g2111(n1495 ,n39[0] ,n1466);
    nor g2112(n1494 ,n39[1] ,n1469);
    or g2113(n1493 ,n38[1] ,n1344);
    or g2114(n1492 ,n1433 ,n1349);
    xnor g2115(n1491 ,n963 ,n41[0]);
    xnor g2116(n1490 ,n953 ,n52[2]);
    xnor g2117(n1489 ,n949 ,n52[4]);
    xnor g2118(n1488 ,n953 ,n51[2]);
    xnor g2119(n1487 ,n954 ,n51[10]);
    xnor g2120(n1486 ,n948 ,n53[15]);
    xnor g2121(n1485 ,n946 ,n53[14]);
    xnor g2122(n1484 ,n947 ,n53[3]);
    xnor g2123(n1483 ,n958 ,n53[7]);
    xnor g2124(n1482 ,n952 ,n53[5]);
    xnor g2125(n1481 ,n957 ,n53[8]);
    xnor g2126(n1480 ,n950 ,n50[6]);
    xnor g2127(n1479 ,n947 ,n50[3]);
    xnor g2128(n1478 ,n953 ,n50[2]);
    xnor g2129(n1477 ,n960 ,n52[11]);
    xnor g2130(n1476 ,n957 ,n51[8]);
    xnor g2131(n1475 ,n959 ,n53[9]);
    not g2132(n1464 ,n1465);
    nor g2133(n1462 ,n1020 ,n41[11]);
    nor g2134(n1461 ,n965 ,n41[0]);
    or g2135(n1460 ,n964 ,n38[2]);
    nor g2136(n1459 ,n966 ,n41[0]);
    nor g2137(n1458 ,n968 ,n41[0]);
    nor g2138(n1457 ,n1027 ,n964);
    nor g2139(n1456 ,n943 ,n630);
    nor g2140(n1455 ,n1029 ,n41[5]);
    nor g2141(n1454 ,n1002 ,n41[1]);
    nor g2142(n1453 ,n1168 ,n539);
    nor g2143(n1452 ,n1169 ,n540);
    nor g2144(n1451 ,n1171 ,n540);
    nor g2145(n1450 ,n987 ,n41[15]);
    nor g2146(n1449 ,n1015 ,n41[7]);
    nor g2147(n1448 ,n991 ,n41[13]);
    nor g2148(n1447 ,n998 ,n41[3]);
    nor g2149(n1446 ,n997 ,n41[8]);
    nor g2150(n1445 ,n993 ,n41[14]);
    nor g2151(n1444 ,n985 ,n41[12]);
    nor g2152(n1443 ,n1004 ,n41[9]);
    nor g2153(n1442 ,n992 ,n41[6]);
    nor g2154(n1441 ,n990 ,n41[13]);
    nor g2155(n1440 ,n975 ,n41[1]);
    nor g2156(n1439 ,n1003 ,n41[7]);
    nor g2157(n1438 ,n1013 ,n41[9]);
    nor g2158(n1437 ,n976 ,n41[12]);
    nor g2159(n1436 ,n971 ,n41[10]);
    nor g2160(n1435 ,n986 ,n41[1]);
    nor g2161(n1434 ,n828 ,n38[0]);
    nor g2162(n1433 ,n1011 ,n41[10]);
    nor g2163(n1432 ,n988 ,n41[6]);
    nor g2164(n1431 ,n1008 ,n41[13]);
    nor g2165(n1430 ,n1010 ,n41[12]);
    nor g2166(n1429 ,n995 ,n41[10]);
    nor g2167(n1428 ,n1035 ,n41[5]);
    nor g2168(n1427 ,n1019 ,n41[6]);
    nor g2169(n1426 ,n972 ,n41[8]);
    nor g2170(n1425 ,n1022 ,n41[4]);
    nor g2171(n1424 ,n974 ,n41[14]);
    nor g2172(n1423 ,n1012 ,n41[15]);
    nor g2173(n1422 ,n1034 ,n41[7]);
    nor g2174(n1421 ,n978 ,n41[9]);
    nor g2175(n1420 ,n1016 ,n41[11]);
    or g2176(n1419 ,n996 ,n38[1]);
    nor g2177(n1418 ,n1018 ,n41[4]);
    nor g2178(n1417 ,n1025 ,n41[12]);
    nor g2179(n1416 ,n973 ,n41[15]);
    or g2180(n1415 ,n983 ,n43[0]);
    nor g2181(n1414 ,n1000 ,n41[3]);
    nor g2182(n1413 ,n984 ,n41[11]);
    nor g2183(n1412 ,n979 ,n41[5]);
    nor g2184(n1411 ,n1014 ,n41[13]);
    nor g2185(n1410 ,n982 ,n41[14]);
    nor g2186(n1409 ,n1024 ,n41[2]);
    nor g2187(n1408 ,n1030 ,n41[4]);
    nor g2188(n1407 ,n1026 ,n41[1]);
    or g2189(n1474 ,n980 ,n543);
    or g2190(n1473 ,n1027 ,n43[0]);
    or g2191(n1472 ,n994 ,n543);
    or g2192(n1471 ,n977 ,n543);
    or g2193(n1470 ,n1032 ,n537);
    nor g2194(n1469 ,n994 ,n546);
    nor g2195(n1468 ,n980 ,n545);
    nor g2196(n1467 ,n977 ,n547);
    nor g2197(n1466 ,n1032 ,n548);
    nor g2198(n1465 ,n549 ,n3258);
    or g2199(n1463 ,n983 ,n43[2]);
    not g2200(n1404 ,n1403);
    nor g2201(n1399 ,n954 ,n53[10]);
    or g2202(n1398 ,n35[1] ,n35[2]);
    nor g2203(n1397 ,n945 ,n541);
    nor g2204(n1396 ,n957 ,n50[8]);
    nor g2205(n1395 ,n956 ,n52[13]);
    nor g2206(n1394 ,n959 ,n50[9]);
    nor g2207(n1393 ,n946 ,n52[14]);
    nor g2208(n1392 ,n947 ,n52[3]);
    nor g2209(n1391 ,n957 ,n52[8]);
    nor g2210(n1390 ,n951 ,n51[0]);
    nor g2211(n1389 ,n959 ,n51[9]);
    nor g2212(n1388 ,n950 ,n52[6]);
    nor g2213(n1387 ,n950 ,n53[6]);
    nor g2214(n1386 ,n944 ,n53[1]);
    nor g2215(n1385 ,n949 ,n51[4]);
    nor g2216(n1384 ,n955 ,n50[12]);
    nor g2217(n1383 ,n952 ,n52[5]);
    nor g2218(n1382 ,n952 ,n50[5]);
    nor g2219(n1381 ,n954 ,n50[10]);
    nor g2220(n1380 ,n944 ,n52[1]);
    nor g2221(n1379 ,n944 ,n50[1]);
    nor g2222(n1378 ,n953 ,n53[2]);
    nor g2223(n1377 ,n960 ,n50[11]);
    nor g2224(n1376 ,n949 ,n50[4]);
    nor g2225(n1375 ,n960 ,n51[11]);
    nor g2226(n1374 ,n946 ,n50[14]);
    nor g2227(n1373 ,n960 ,n53[11]);
    nor g2228(n1372 ,n955 ,n53[12]);
    nor g2229(n1371 ,n946 ,n51[14]);
    nor g2230(n1370 ,n958 ,n51[7]);
    nor g2231(n1369 ,n956 ,n51[13]);
    nor g2232(n1368 ,n954 ,n52[10]);
    or g2233(n1367 ,n36[0] ,n36[1]);
    or g2234(n1366 ,n967 ,n38[0]);
    nor g2235(n1365 ,n959 ,n52[9]);
    nor g2236(n1364 ,n951 ,n53[0]);
    nor g2237(n1363 ,n951 ,n50[0]);
    nor g2238(n1362 ,n949 ,n53[4]);
    nor g2239(n1361 ,n944 ,n51[1]);
    nor g2240(n1360 ,n948 ,n50[15]);
    nor g2241(n1359 ,n956 ,n50[13]);
    nor g2242(n1358 ,n958 ,n50[7]);
    nor g2243(n1357 ,n950 ,n51[6]);
    nor g2244(n1356 ,n955 ,n52[12]);
    nor g2245(n1355 ,n952 ,n51[5]);
    nor g2246(n1354 ,n955 ,n51[12]);
    nor g2247(n1353 ,n948 ,n51[15]);
    nor g2248(n1352 ,n947 ,n51[3]);
    nor g2249(n1351 ,n958 ,n52[7]);
    nor g2250(n1350 ,n948 ,n52[15]);
    nor g2251(n1349 ,n956 ,n53[13]);
    nor g2252(n1348 ,n943 ,n3[1]);
    or g2253(n1347 ,n39[0] ,n39[1]);
    or g2254(n1346 ,n37[2] ,n37[3]);
    or g2255(n1345 ,n2[1] ,n2[0]);
    nor g2256(n1344 ,n38[0] ,n3[0]);
    or g2257(n1343 ,n39[2] ,n39[3]);
    or g2258(n1342 ,n2[3] ,n2[2]);
    or g2259(n1341 ,n35[0] ,n35[3]);
    or g2260(n1340 ,n36[2] ,n36[3]);
    or g2261(n1339 ,n37[0] ,n37[1]);
    or g2262(n1406 ,n943 ,n38[2]);
    or g2263(n1405 ,n945 ,n43[1]);
    nor g2264(n1403 ,n43[0] ,n43[1]);
    or g2265(n1402 ,n962 ,n38[3]);
    or g2266(n1401 ,n38[0] ,n38[2]);
    or g2267(n1400 ,n38[1] ,n38[3]);
    not g2268(n1338 ,n12[31]);
    not g2269(n1337 ,n14[0]);
    not g2270(n1336 ,n15[13]);
    not g2271(n1335 ,n5[18]);
    not g2272(n1334 ,n8[11]);
    not g2273(n1333 ,n3339);
    not g2274(n1332 ,n3298);
    not g2275(n1331 ,n3379);
    not g2276(n1330 ,n10[2]);
    not g2277(n1329 ,n14[1]);
    not g2278(n1328 ,n10[0]);
    not g2279(n1327 ,n3287);
    not g2280(n1326 ,n15[3]);
    not g2281(n1325 ,n15[12]);
    not g2282(n1324 ,n21[1]);
    not g2283(n1323 ,n8[2]);
    not g2284(n1322 ,n4[27]);
    not g2285(n1321 ,n3377);
    not g2286(n1320 ,n10[20]);
    not g2287(n1319 ,n5[11]);
    not g2288(n1318 ,n15[0]);
    not g2289(n1317 ,n10[26]);
    not g2290(n1316 ,n11[3]);
    not g2291(n1315 ,n13[7]);
    not g2292(n1314 ,n3376);
    not g2293(n1313 ,n8[15]);
    not g2294(n1312 ,n19[1]);
    not g2295(n1311 ,n3282);
    not g2296(n1310 ,n5[16]);
    not g2297(n1309 ,n3362);
    not g2298(n1308 ,n6[23]);
    not g2299(n1307 ,n3361);
    not g2300(n1306 ,n4[18]);
    not g2301(n1305 ,n3306);
    not g2302(n1304 ,n4[17]);
    not g2303(n1303 ,n3357);
    not g2304(n1302 ,n3356);
    not g2305(n1301 ,n8[28]);
    not g2306(n1300 ,n12[11]);
    not g2307(n1299 ,n9[31]);
    not g2308(n1298 ,n9[30]);
    not g2309(n1297 ,n10[9]);
    not g2310(n1296 ,n4[3]);
    not g2311(n1295 ,n5[28]);
    not g2312(n1294 ,n14[12]);
    not g2313(n1293 ,n15[6]);
    not g2314(n1292 ,n14[15]);
    not g2315(n1291 ,n11[12]);
    not g2316(n1290 ,n14[14]);
    not g2317(n1289 ,n5[1]);
    not g2318(n1288 ,n3346);
    not g2319(n1287 ,n13[12]);
    not g2320(n1286 ,n3283);
    not g2321(n1285 ,n6[27]);
    not g2322(n1284 ,n3295);
    not g2323(n1283 ,n16[8]);
    not g2324(n1282 ,n10[4]);
    not g2325(n1281 ,n10[22]);
    not g2326(n1280 ,n15[10]);
    not g2327(n1279 ,n8[24]);
    not g2328(n1278 ,n14[7]);
    not g2329(n1277 ,n5[20]);
    not g2330(n1276 ,n10[27]);
    not g2331(n1275 ,n12[30]);
    not g2332(n1274 ,n6[1]);
    not g2333(n1273 ,n8[29]);
    not g2334(n1272 ,n3358);
    not g2335(n1271 ,n7[8]);
    not g2336(n1270 ,n4[5]);
    not g2337(n1269 ,n8[14]);
    not g2338(n1268 ,n6[22]);
    not g2339(n1267 ,n3307);
    not g2340(n1266 ,n9[9]);
    not g2341(n1265 ,n16[5]);
    not g2342(n1264 ,n13[15]);
    not g2343(n1263 ,n10[18]);
    not g2344(n1262 ,n14[5]);
    not g2345(n1261 ,n6[16]);
    not g2346(n1260 ,n4[29]);
    not g2347(n1259 ,n3327);
    not g2348(n1258 ,n3348);
    not g2349(n1257 ,n11[19]);
    not g2350(n1256 ,n7[29]);
    not g2351(n1255 ,n49[6]);
    not g2352(n1254 ,n49[7]);
    not g2353(n1253 ,n42[1]);
    not g2354(n1252 ,n42[16]);
    not g2355(n1251 ,n25[30]);
    not g2356(n1250 ,n42[0]);
    not g2357(n1249 ,n25[31]);
    not g2358(n1248 ,n25[25]);
    not g2359(n1247 ,n40[25]);
    not g2360(n1246 ,n25[24]);
    not g2361(n1245 ,n26[2]);
    not g2362(n1244 ,n46[7]);
    not g2363(n1243 ,n48[2]);
    not g2364(n1242 ,n42[8]);
    not g2365(n1241 ,n25[12]);
    not g2366(n1240 ,n29[0]);
    not g2367(n1239 ,n26[0]);
    not g2368(n1238 ,n42[4]);
    not g2369(n1237 ,n26[17]);
    not g2370(n1236 ,n40[20]);
    not g2371(n1235 ,n25[11]);
    not g2372(n1234 ,n40[15]);
    not g2373(n1233 ,n40[2]);
    not g2374(n1232 ,n26[29]);
    not g2375(n1231 ,n32[3]);
    not g2376(n1230 ,n31[3]);
    not g2377(n1229 ,n40[10]);
    not g2378(n1228 ,n40[23]);
    not g2379(n1227 ,n31[7]);
    not g2380(n1226 ,n31[2]);
    not g2381(n1225 ,n40[7]);
    not g2382(n1224 ,n46[8]);
    not g2383(n1223 ,n49[5]);
    not g2384(n1222 ,n30[1]);
    not g2385(n1221 ,n26[18]);
    not g2386(n1220 ,n25[16]);
    not g2387(n1219 ,n29[1]);
    not g2388(n1218 ,n48[4]);
    not g2389(n1217 ,n31[4]);
    not g2390(n1216 ,n47[4]);
    not g2391(n1215 ,n25[14]);
    not g2392(n1214 ,n26[8]);
    not g2393(n1213 ,n40[31]);
    not g2394(n1212 ,n34[3]);
    not g2395(n1211 ,n26[23]);
    not g2396(n1210 ,n30[0]);
    not g2397(n1209 ,n40[13]);
    not g2398(n1208 ,n46[4]);
    not g2399(n1207 ,n34[9]);
    not g2400(n1206 ,n42[20]);
    not g2401(n1205 ,n30[3]);
    not g2402(n1204 ,n34[11]);
    not g2403(n1203 ,n34[10]);
    not g2404(n1202 ,n46[9]);
    not g2405(n1201 ,n25[9]);
    not g2406(n1200 ,n42[7]);
    not g2407(n1199 ,n42[17]);
    not g2408(n1198 ,n48[1]);
    not g2409(n1197 ,n27);
    not g2410(n1196 ,n48[3]);
    not g2411(n1195 ,n32[2]);
    not g2412(n1194 ,n34[8]);
    not g2413(n1193 ,n42[10]);
    not g2414(n1192 ,n34[7]);
    not g2415(n1191 ,n40[1]);
    not g2416(n1190 ,n26[26]);
    not g2417(n1189 ,n26[25]);
    not g2418(n1188 ,n42[11]);
    not g2419(n1187 ,n25[20]);
    not g2420(n1186 ,n34[6]);
    not g2421(n1185 ,n26[15]);
    not g2422(n1184 ,n25[8]);
    not g2423(n1183 ,n42[12]);
    not g2424(n1182 ,n26[16]);
    not g2425(n1181 ,n25[26]);
    not g2426(n1180 ,n42[2]);
    not g2427(n1179 ,n34[5]);
    not g2428(n1178 ,n25[22]);
    not g2429(n1177 ,n42[14]);
    not g2430(n1176 ,n31[5]);
    not g2431(n1175 ,n25[23]);
    not g2432(n1174 ,n31[1]);
    not g2433(n1173 ,n34[4]);
    not g2434(n1172 ,n42[13]);
    not g2435(n1171 ,n45[2]);
    not g2436(n1170 ,n46[2]);
    not g2437(n1169 ,n45[0]);
    not g2438(n1168 ,n45[1]);
    not g2439(n1167 ,n40[12]);
    not g2440(n1166 ,n40[28]);
    not g2441(n1165 ,n26[20]);
    not g2442(n1164 ,n40[6]);
    not g2443(n1163 ,n26[28]);
    not g2444(n1162 ,n40[30]);
    not g2445(n1161 ,n48[8]);
    not g2446(n1160 ,n34[2]);
    not g2447(n1159 ,n42[18]);
    not g2448(n1158 ,n40[0]);
    not g2449(n1157 ,n25[7]);
    not g2450(n1156 ,n49[3]);
    not g2451(n1155 ,n30[2]);
    not g2452(n1154 ,n42[19]);
    not g2453(n1153 ,n34[1]);
    not g2454(n1152 ,n42[31]);
    not g2455(n1151 ,n40[17]);
    not g2456(n1150 ,n26[7]);
    not g2457(n1149 ,n25[18]);
    not g2458(n1148 ,n40[24]);
    not g2459(n1147 ,n49[4]);
    not g2460(n1146 ,n48[9]);
    not g2461(n1145 ,n40[22]);
    not g2462(n1144 ,n40[14]);
    not g2463(n1143 ,n26[24]);
    not g2464(n1142 ,n31[0]);
    not g2465(n1141 ,n40[16]);
    not g2466(n1140 ,n47[5]);
    not g2467(n1139 ,n34[14]);
    not g2468(n1138 ,n26[14]);
    not g2469(n1137 ,n42[23]);
    not g2470(n1136 ,n40[21]);
    not g2471(n1135 ,n25[6]);
    not g2472(n1134 ,n40[27]);
    not g2473(n1133 ,n26[19]);
    not g2474(n1132 ,n26[12]);
    not g2475(n1131 ,n42[24]);
    not g2476(n1130 ,n42[5]);
    not g2477(n1129 ,n34[13]);
    not g2478(n1128 ,n25[19]);
    not g2479(n1127 ,n34[15]);
    not g2480(n1126 ,n25[29]);
    not g2481(n1125 ,n42[15]);
    not g2482(n1124 ,n49[9]);
    not g2483(n1123 ,n31[6]);
    not g2484(n1122 ,n42[26]);
    not g2485(n1121 ,n34[12]);
    not g2486(n1120 ,n25[2]);
    not g2487(n1119 ,n47[3]);
    not g2488(n1118 ,n42[30]);
    not g2489(n1117 ,n42[25]);
    not g2490(n1116 ,n42[3]);
    not g2491(n1115 ,n46[5]);
    not g2492(n1114 ,n25[21]);
    not g2493(n1113 ,n26[1]);
    not g2494(n1112 ,n49[2]);
    not g2495(n1111 ,n26[31]);
    not g2496(n1110 ,n25[28]);
    not g2497(n1109 ,n42[29]);
    not g2498(n1108 ,n40[9]);
    not g2499(n1107 ,n26[13]);
    not g2500(n1106 ,n40[18]);
    not g2501(n1105 ,n25[5]);
    not g2502(n1104 ,n40[11]);
    not g2503(n1103 ,n26[10]);
    not g2504(n1102 ,n46[1]);
    not g2505(n1101 ,n42[28]);
    not g2506(n1100 ,n25[10]);
    not g2507(n1099 ,n42[22]);
    not g2508(n1098 ,n48[5]);
    not g2509(n1097 ,n42[6]);
    not g2510(n1096 ,n26[9]);
    not g2511(n1095 ,n25[1]);
    not g2512(n1094 ,n26[11]);
    not g2513(n1093 ,n47[6]);
    not g2514(n1092 ,n32[0]);
    not g2515(n1091 ,n40[19]);
    not g2516(n1090 ,n26[22]);
    not g2517(n1089 ,n42[27]);
    not g2518(n1088 ,n25[4]);
    not g2519(n1087 ,n49[8]);
    not g2520(n1086 ,n40[3]);
    not g2521(n1085 ,n42[21]);
    not g2522(n1084 ,n40[29]);
    not g2523(n1083 ,n46[6]);
    not g2524(n1082 ,n25[15]);
    not g2525(n1081 ,n40[5]);
    not g2526(n1080 ,n40[4]);
    not g2527(n1079 ,n25[0]);
    not g2528(n1078 ,n48[7]);
    not g2529(n1077 ,n47[7]);
    not g2530(n1076 ,n25[3]);
    not g2531(n1075 ,n40[26]);
    not g2532(n1074 ,n25[27]);
    not g2533(n1073 ,n25[13]);
    not g2534(n1072 ,n26[27]);
    not g2535(n1071 ,n32[1]);
    not g2536(n1070 ,n46[3]);
    not g2537(n1069 ,n26[4]);
    not g2538(n1068 ,n28);
    not g2539(n1067 ,n47[2]);
    not g2540(n1066 ,n26[3]);
    not g2541(n1065 ,n26[5]);
    not g2542(n1064 ,n29[3]);
    not g2543(n1063 ,n47[1]);
    not g2544(n1062 ,n48[6]);
    not g2545(n1061 ,n29[2]);
    not g2546(n1060 ,n25[17]);
    not g2547(n1059 ,n49[1]);
    not g2548(n1058 ,n26[6]);
    not g2549(n1057 ,n26[30]);
    not g2550(n1056 ,n40[8]);
    not g2551(n1055 ,n42[9]);
    not g2552(n1054 ,n47[9]);
    not g2553(n1053 ,n47[8]);
    not g2554(n1052 ,n26[21]);
    not g2555(n1051 ,n37[2]);
    not g2556(n1050 ,n48[0]);
    not g2557(n1049 ,n36[0]);
    not g2558(n1048 ,n37[1]);
    not g2559(n1047 ,n36[3]);
    not g2560(n1046 ,n36[2]);
    not g2561(n1045 ,n47[0]);
    not g2562(n1044 ,n37[0]);
    not g2563(n1043 ,n49[0]);
    not g2564(n1042 ,n46[0]);
    not g2565(n1041 ,n36[1]);
    not g2566(n1040 ,n39[3]);
    not g2567(n1039 ,n37[3]);
    not g2568(n1038 ,n39[2]);
    not g2569(n1037 ,n39[0]);
    not g2570(n1036 ,n39[1]);
    not g2571(n1035 ,n50[5]);
    not g2572(n1034 ,n50[7]);
    not g2573(n1033 ,n51[8]);
    not g2574(n1032 ,n35[0]);
    not g2575(n1031 ,n53[8]);
    not g2576(n1030 ,n51[4]);
    not g2577(n1029 ,n52[5]);
    not g2578(n1028 ,n50[6]);
    not g2579(n1027 ,n44[0]);
    not g2580(n1026 ,n53[1]);
    not g2581(n1025 ,n50[12]);
    not g2582(n1024 ,n53[2]);
    not g2583(n1023 ,n53[3]);
    not g2584(n1022 ,n53[4]);
    not g2585(n1021 ,n53[5]);
    not g2586(n1020 ,n53[11]);
    not g2587(n1019 ,n53[6]);
    not g2588(n1018 ,n50[4]);
    not g2589(n1017 ,n53[7]);
    not g2590(n1016 ,n50[11]);
    not g2591(n1015 ,n51[7]);
    not g2592(n1014 ,n51[13]);
    not g2593(n1013 ,n51[9]);
    not g2594(n1012 ,n50[15]);
    not g2595(n1011 ,n53[10]);
    not g2596(n1010 ,n53[12]);
    not g2597(n1009 ,n51[10]);
    not g2598(n1008 ,n53[13]);
    not g2599(n1007 ,n53[14]);
    not g2600(n1006 ,n53[9]);
    not g2601(n1005 ,n53[15]);
    not g2602(n1004 ,n52[9]);
    not g2603(n1003 ,n52[7]);
    not g2604(n1002 ,n52[1]);
    not g2605(n1001 ,n52[2]);
    not g2606(n1000 ,n52[3]);
    not g2607(n999 ,n50[3]);
    not g2608(n998 ,n51[3]);
    not g2609(n997 ,n52[8]);
    not g2610(n996 ,n38[3]);
    not g2611(n995 ,n52[10]);
    not g2612(n994 ,n35[1]);
    not g2613(n993 ,n52[14]);
    not g2614(n992 ,n52[6]);
    not g2615(n991 ,n50[13]);
    not g2616(n990 ,n52[13]);
    not g2617(n989 ,n52[11]);
    not g2618(n988 ,n51[6]);
    not g2619(n987 ,n51[15]);
    not g2620(n986 ,n51[1]);
    not g2621(n985 ,n52[12]);
    not g2622(n984 ,n51[11]);
    not g2623(n983 ,n43[1]);
    not g2624(n982 ,n51[14]);
    not g2625(n981 ,n51[2]);
    not g2626(n980 ,n35[2]);
    not g2627(n979 ,n51[5]);
    not g2628(n978 ,n50[9]);
    not g2629(n977 ,n35[3]);
    not g2630(n976 ,n51[12]);
    not g2631(n975 ,n50[1]);
    not g2632(n974 ,n50[14]);
    not g2633(n973 ,n52[15]);
    not g2634(n972 ,n50[8]);
    not g2635(n971 ,n50[10]);
    not g2636(n970 ,n52[4]);
    not g2637(n969 ,n50[2]);
    not g2638(n968 ,n50[0]);
    not g2639(n967 ,n38[2]);
    not g2640(n966 ,n53[0]);
    not g2641(n965 ,n51[0]);
    not g2642(n964 ,n44[1]);
    not g2643(n963 ,n52[0]);
    not g2644(n962 ,n38[1]);
    not g2645(n961 ,n43[2]);
    not g2646(n960 ,n41[11]);
    not g2647(n959 ,n41[9]);
    not g2648(n958 ,n41[7]);
    not g2649(n957 ,n41[8]);
    not g2650(n956 ,n41[13]);
    not g2651(n955 ,n41[12]);
    not g2652(n954 ,n41[10]);
    not g2653(n953 ,n41[2]);
    not g2654(n952 ,n41[5]);
    not g2655(n951 ,n41[0]);
    not g2656(n950 ,n41[6]);
    not g2657(n949 ,n41[4]);
    not g2658(n948 ,n41[15]);
    not g2659(n947 ,n41[3]);
    not g2660(n946 ,n41[14]);
    not g2661(n945 ,n43[0]);
    not g2662(n944 ,n41[1]);
    not g2663(n943 ,n38[0]);
    not g2664(n942 ,n16[15]);
    not g2665(n941 ,n10[8]);
    not g2666(n940 ,n9[8]);
    not g2667(n939 ,n3319);
    not g2668(n938 ,n3317);
    not g2669(n937 ,n13[6]);
    not g2670(n936 ,n5[10]);
    not g2671(n935 ,n8[7]);
    not g2672(n934 ,n9[2]);
    not g2673(n933 ,n6[3]);
    not g2674(n932 ,n3280);
    not g2675(n931 ,n3331);
    not g2676(n930 ,n4[19]);
    not g2677(n929 ,n3330);
    not g2678(n928 ,n11[27]);
    not g2679(n927 ,n17[1]);
    not g2680(n926 ,n7[1]);
    not g2681(n925 ,n4[25]);
    not g2682(n924 ,n7[24]);
    not g2683(n923 ,n9[10]);
    not g2684(n922 ,n4[9]);
    not g2685(n921 ,n3303);
    not g2686(n920 ,n7[4]);
    not g2687(n919 ,n11[14]);
    not g2688(n918 ,n13[5]);
    not g2689(n917 ,n16[10]);
    not g2690(n916 ,n15[4]);
    not g2691(n915 ,n11[11]);
    not g2692(n914 ,n12[24]);
    not g2693(n913 ,n13[10]);
    not g2694(n912 ,n6[25]);
    not g2695(n911 ,n14[8]);
    not g2696(n910 ,n13[2]);
    not g2697(n909 ,n9[19]);
    not g2698(n908 ,n11[9]);
    not g2699(n907 ,n3286);
    not g2700(n906 ,n11[2]);
    not g2701(n905 ,n14[2]);
    not g2702(n904 ,n10[16]);
    not g2703(n903 ,n14[3]);
    not g2704(n902 ,n15[15]);
    not g2705(n901 ,n12[0]);
    not g2706(n900 ,n15[5]);
    not g2707(n899 ,n16[6]);
    not g2708(n898 ,n3281);
    not g2709(n897 ,n7[26]);
    not g2710(n896 ,n7[15]);
    not g2711(n895 ,n12[5]);
    not g2712(n894 ,n3365);
    not g2713(n893 ,n4[12]);
    not g2714(n892 ,n3318);
    not g2715(n891 ,n9[26]);
    not g2716(n890 ,n3294);
    not g2717(n889 ,n3347);
    not g2718(n888 ,n4[11]);
    not g2719(n887 ,n3309);
    not g2720(n886 ,n10[24]);
    not g2721(n885 ,n13[11]);
    not g2722(n884 ,n6[20]);
    not g2723(n883 ,n3276);
    not g2724(n882 ,n6[17]);
    not g2725(n881 ,n7[14]);
    not g2726(n880 ,n15[7]);
    not g2727(n879 ,n3332);
    not g2728(n878 ,n5[5]);
    not g2729(n877 ,n12[3]);
    not g2730(n876 ,n3370);
    not g2731(n875 ,n11[5]);
    not g2732(n874 ,n12[19]);
    not g2733(n873 ,n9[5]);
    not g2734(n872 ,n6[28]);
    not g2735(n871 ,n3308);
    not g2736(n870 ,n10[10]);
    not g2737(n869 ,n4[1]);
    not g2738(n868 ,n3311);
    not g2739(n867 ,n4[30]);
    not g2740(n866 ,n3314);
    not g2741(n865 ,n14[4]);
    not g2742(n864 ,n3363);
    not g2743(n863 ,n3382);
    not g2744(n862 ,n3329);
    not g2745(n861 ,n7[16]);
    not g2746(n860 ,n6[30]);
    not g2747(n859 ,n3310);
    not g2748(n858 ,n8[17]);
    not g2749(n857 ,n4[7]);
    not g2750(n856 ,n3359);
    not g2751(n855 ,n3320);
    not g2752(n854 ,n3374);
    not g2753(n853 ,n3277);
    not g2754(n852 ,n9[20]);
    not g2755(n851 ,n3354);
    not g2756(n850 ,n12[13]);
    not g2757(n849 ,n9[7]);
    not g2758(n848 ,n11[25]);
    not g2759(n847 ,n8[8]);
    not g2760(n846 ,n3323);
    not g2761(n845 ,n12[25]);
    not g2762(n844 ,n8[19]);
    not g2763(n843 ,n7[7]);
    not g2764(n842 ,n9[18]);
    not g2765(n841 ,n11[8]);
    not g2766(n840 ,n11[0]);
    not g2767(n839 ,n3326);
    not g2768(n838 ,n15[8]);
    not g2769(n837 ,n8[26]);
    not g2770(n836 ,n7[9]);
    not g2771(n835 ,n9[21]);
    not g2772(n834 ,n10[19]);
    not g2773(n833 ,n8[25]);
    not g2774(n832 ,n10[11]);
    not g2775(n831 ,n10[12]);
    not g2776(n830 ,n13[14]);
    not g2777(n829 ,n4[20]);
    not g2778(n828 ,n3[2]);
    not g2779(n827 ,n3366);
    not g2780(n826 ,n9[28]);
    not g2781(n825 ,n12[6]);
    not g2782(n824 ,n9[23]);
    not g2783(n823 ,n7[23]);
    not g2784(n822 ,n5[26]);
    not g2785(n821 ,n4[8]);
    not g2786(n820 ,n3304);
    not g2787(n819 ,n16[12]);
    not g2788(n818 ,n7[21]);
    not g2789(n817 ,n12[29]);
    not g2790(n816 ,n10[1]);
    not g2791(n815 ,n3274);
    not g2792(n814 ,n7[25]);
    not g2793(n813 ,n5[12]);
    not g2794(n812 ,n3328);
    not g2795(n811 ,n16[9]);
    not g2796(n810 ,n3302);
    not g2797(n809 ,n12[14]);
    not g2798(n808 ,n3345);
    not g2799(n807 ,n14[10]);
    not g2800(n806 ,n3296);
    not g2801(n805 ,n3341);
    not g2802(n804 ,n11[4]);
    not g2803(n803 ,n12[23]);
    not g2804(n802 ,n5[0]);
    not g2805(n801 ,n10[15]);
    not g2806(n800 ,n6[26]);
    not g2807(n799 ,n13[9]);
    not g2808(n798 ,n3334);
    not g2809(n797 ,n9[14]);
    not g2810(n796 ,n3352);
    not g2811(n795 ,n7[27]);
    not g2812(n794 ,n5[31]);
    not g2813(n793 ,n3360);
    not g2814(n792 ,n3344);
    not g2815(n791 ,n3297);
    not g2816(n790 ,n9[27]);
    not g2817(n789 ,n23[0]);
    not g2818(n788 ,n3380);
    not g2819(n787 ,n12[4]);
    not g2820(n786 ,n7[19]);
    not g2821(n785 ,n8[27]);
    not g2822(n784 ,n5[15]);
    not g2823(n783 ,n3305);
    not g2824(n782 ,n10[7]);
    not g2825(n781 ,n9[25]);
    not g2826(n780 ,n10[14]);
    not g2827(n779 ,n4[31]);
    not g2828(n778 ,n6[15]);
    not g2829(n777 ,n3284);
    not g2830(n776 ,n12[26]);
    not g2831(n775 ,n23[1]);
    not g2832(n774 ,n3325);
    not g2833(n773 ,n8[16]);
    not g2834(n772 ,n10[25]);
    not g2835(n771 ,n15[9]);
    not g2836(n770 ,n9[24]);
    not g2837(n769 ,n4[10]);
    not g2838(n768 ,n10[3]);
    not g2839(n767 ,n3371);
    not g2840(n766 ,n5[21]);
    not g2841(n765 ,n9[17]);
    not g2842(n764 ,n10[13]);
    not g2843(n763 ,n9[15]);
    not g2844(n762 ,n16[13]);
    not g2845(n761 ,n16[11]);
    not g2846(n760 ,n8[21]);
    not g2847(n759 ,n8[0]);
    not g2848(n758 ,n5[17]);
    not g2849(n757 ,n16[7]);
    not g2850(n756 ,n3299);
    not g2851(n755 ,n11[15]);
    not g2852(n754 ,n3293);
    not g2853(n753 ,n4[24]);
    not g2854(n752 ,n13[0]);
    not g2855(n751 ,n10[28]);
    not g2856(n750 ,n4[2]);
    not g2857(n749 ,n3292);
    not g2858(n748 ,n16[4]);
    not g2859(n747 ,n14[6]);
    not g2860(n746 ,n5[23]);
    not g2861(n745 ,n5[27]);
    not g2862(n744 ,n6[13]);
    not g2863(n743 ,n3290);
    not g2864(n742 ,n3338);
    not g2865(n741 ,n6[8]);
    not g2866(n740 ,n3272);
    not g2867(n739 ,n10[31]);
    not g2868(n738 ,n6[5]);
    not g2869(n737 ,n12[28]);
    not g2870(n736 ,n11[7]);
    not g2871(n735 ,n3369);
    not g2872(n734 ,n4[22]);
    not g2873(n733 ,n11[1]);
    not g2874(n732 ,n9[16]);
    not g2875(n731 ,n6[12]);
    not g2876(n730 ,n12[22]);
    not g2877(n729 ,n4[15]);
    not g2878(n728 ,n11[23]);
    not g2879(n727 ,n6[29]);
    not g2880(n726 ,n3300);
    not g2881(n725 ,n3350);
    not g2882(n724 ,n7[3]);
    not g2883(n723 ,n3315);
    not g2884(n722 ,n13[4]);
    not g2885(n721 ,n3343);
    not g2886(n720 ,n7[12]);
    not g2887(n719 ,n16[14]);
    not g2888(n718 ,n7[0]);
    not g2889(n717 ,n3313);
    not g2890(n716 ,n12[7]);
    not g2891(n715 ,n10[17]);
    not g2892(n714 ,n3364);
    not g2893(n713 ,n3288);
    not g2894(n712 ,n6[11]);
    not g2895(n711 ,n8[31]);
    not g2896(n710 ,n3279);
    not g2897(n709 ,n11[21]);
    not g2898(n708 ,n12[1]);
    not g2899(n707 ,n11[18]);
    not g2900(n706 ,n6[21]);
    not g2901(n705 ,n12[10]);
    not g2902(n704 ,n3351);
    not g2903(n703 ,n7[2]);
    not g2904(n702 ,n3271);
    not g2905(n701 ,n6[14]);
    not g2906(n700 ,n13[3]);
    not g2907(n699 ,n3291);
    not g2908(n698 ,n3301);
    not g2909(n697 ,n12[2]);
    not g2910(n696 ,n11[26]);
    not g2911(n695 ,n7[17]);
    not g2912(n694 ,n7[22]);
    not g2913(n693 ,n5[24]);
    not g2914(n692 ,n7[10]);
    not g2915(n691 ,n3336);
    not g2916(n690 ,n8[6]);
    not g2917(n689 ,n5[30]);
    not g2918(n688 ,n5[6]);
    not g2919(n687 ,n4[4]);
    not g2920(n686 ,n6[6]);
    not g2921(n685 ,n8[13]);
    not g2922(n684 ,n5[25]);
    not g2923(n683 ,n3337);
    not g2924(n682 ,n7[13]);
    not g2925(n681 ,n5[8]);
    not g2926(n680 ,n8[5]);
    not g2927(n679 ,n8[20]);
    not g2928(n678 ,n12[15]);
    not g2929(n677 ,n6[2]);
    not g2930(n676 ,n8[12]);
    not g2931(n675 ,n9[4]);
    not g2932(n674 ,n6[19]);
    not g2933(n673 ,n10[6]);
    not g2934(n672 ,n8[4]);
    not g2935(n671 ,n7[31]);
    not g2936(n670 ,n10[29]);
    not g2937(n669 ,n9[12]);
    not g2938(n668 ,n4[28]);
    not g2939(n667 ,n4[14]);
    not g2940(n666 ,n7[30]);
    not g2941(n665 ,n4[13]);
    not g2942(n664 ,n12[16]);
    not g2943(n663 ,n5[2]);
    not g2944(n662 ,n15[11]);
    not g2945(n661 ,n5[29]);
    not g2946(n660 ,n9[29]);
    not g2947(n659 ,n3372);
    not g2948(n658 ,n8[1]);
    not g2949(n657 ,n3373);
    not g2950(n656 ,n8[22]);
    not g2951(n655 ,n8[23]);
    not g2952(n654 ,n11[29]);
    not g2953(n653 ,n11[31]);
    not g2954(n652 ,n6[9]);
    not g2955(n651 ,n7[6]);
    not g2956(n650 ,n9[1]);
    not g2957(n649 ,n5[13]);
    not g2958(n648 ,n8[3]);
    not g2959(n647 ,n6[18]);
    not g2960(n646 ,n15[1]);
    not g2961(n645 ,n3335);
    not g2962(n644 ,n4[21]);
    not g2963(n643 ,n4[23]);
    not g2964(n642 ,n14[9]);
    not g2965(n641 ,n11[17]);
    not g2966(n640 ,n6[7]);
    not g2967(n639 ,n11[30]);
    not g2968(n638 ,n21[0]);
    not g2969(n637 ,n5[22]);
    not g2970(n636 ,n7[18]);
    not g2971(n635 ,n16[3]);
    not g2972(n634 ,n3349);
    not g2973(n633 ,n12[20]);
    not g2974(n632 ,n3285);
    not g2975(n631 ,n5[9]);
    not g2976(n630 ,n3[3]);
    not g2977(n629 ,n11[13]);
    not g2978(n628 ,n3273);
    not g2979(n627 ,n11[22]);
    not g2980(n626 ,n7[5]);
    not g2981(n625 ,n14[11]);
    not g2982(n624 ,n5[14]);
    not g2983(n623 ,n5[7]);
    not g2984(n622 ,n14[13]);
    not g2985(n621 ,n11[24]);
    not g2986(n620 ,n12[9]);
    not g2987(n619 ,n11[10]);
    not g2988(n618 ,n3381);
    not g2989(n617 ,n9[6]);
    not g2990(n616 ,n10[5]);
    not g2991(n615 ,n9[13]);
    not g2992(n614 ,n10[21]);
    not g2993(n613 ,n3355);
    not g2994(n612 ,n8[30]);
    not g2995(n611 ,n3289);
    not g2996(n610 ,n6[24]);
    not g2997(n609 ,n11[20]);
    not g2998(n608 ,n12[27]);
    not g2999(n607 ,n4[6]);
    not g3000(n606 ,n7[28]);
    not g3001(n605 ,n3278);
    not g3002(n604 ,n3375);
    not g3003(n603 ,n7[20]);
    not g3004(n602 ,n3378);
    not g3005(n601 ,n6[31]);
    not g3006(n600 ,n12[18]);
    not g3007(n599 ,n17[0]);
    not g3008(n598 ,n9[22]);
    not g3009(n597 ,n3340);
    not g3010(n596 ,n12[12]);
    not g3011(n595 ,n8[18]);
    not g3012(n594 ,n16[1]);
    not g3013(n593 ,n19[0]);
    not g3014(n592 ,n3275);
    not g3015(n591 ,n11[6]);
    not g3016(n590 ,n11[16]);
    not g3017(n589 ,n9[0]);
    not g3018(n588 ,n3333);
    not g3019(n587 ,n3316);
    not g3020(n586 ,n15[14]);
    not g3021(n585 ,n13[1]);
    not g3022(n584 ,n3342);
    not g3023(n583 ,n15[2]);
    not g3024(n582 ,n9[3]);
    not g3025(n581 ,n3368);
    not g3026(n580 ,n7[11]);
    not g3027(n579 ,n4[0]);
    not g3028(n578 ,n6[0]);
    not g3029(n577 ,n12[17]);
    not g3030(n576 ,n5[19]);
    not g3031(n575 ,n6[10]);
    not g3032(n574 ,n12[8]);
    not g3033(n573 ,n11[28]);
    not g3034(n572 ,n16[0]);
    not g3035(n571 ,n4[26]);
    not g3036(n570 ,n10[30]);
    not g3037(n569 ,n5[3]);
    not g3038(n568 ,n6[4]);
    not g3039(n567 ,n3312);
    not g3040(n566 ,n12[21]);
    not g3041(n565 ,n13[8]);
    not g3042(n564 ,n3353);
    not g3043(n563 ,n3322);
    not g3044(n562 ,n16[2]);
    not g3045(n561 ,n3321);
    not g3046(n560 ,n8[10]);
    not g3047(n559 ,n13[13]);
    not g3048(n558 ,n4[16]);
    not g3049(n557 ,n8[9]);
    not g3050(n556 ,n3324);
    not g3051(n555 ,n5[4]);
    not g3052(n554 ,n9[11]);
    not g3053(n553 ,n10[23]);
    not g3054(n552 ,n3261);
    not g3055(n551 ,n3259);
    not g3056(n550 ,n3260);
    not g3057(n549 ,n2[3]);
    not g3058(n548 ,n3383);
    not g3059(n547 ,n3386);
    not g3060(n546 ,n3384);
    not g3061(n545 ,n3385);
    not g3062(n544 ,n1);
    not g3063(n543 ,n1);
    not g3064(n542 ,n1);
    not g3065(n541 ,n1);
    not g3066(n540 ,n1);
    not g3067(n539 ,n1);
    not g3068(n538 ,n1);
    not g3069(n537 ,n1);
    or g3070(n3367 ,n18[1] ,n18[0]);
    or g3071(n3268 ,n57 ,n60);
    nor g3072(n60 ,n3269 ,n59);
    or g3073(n59 ,n56 ,n58);
    nor g3074(n58 ,n55 ,n20[1]);
    nor g3075(n57 ,n54 ,n3270);
    not g3076(n56 ,n20[0]);
    not g3077(n55 ,n3270);
    not g3078(n54 ,n20[1]);
    or g3079(n3265 ,n64 ,n67);
    nor g3080(n67 ,n3266 ,n66);
    or g3081(n66 ,n63 ,n65);
    nor g3082(n65 ,n62 ,n22[1]);
    nor g3083(n64 ,n61 ,n3267);
    not g3084(n63 ,n22[0]);
    not g3085(n62 ,n3267);
    not g3086(n61 ,n22[1]);
    or g3087(n3262 ,n71 ,n74);
    nor g3088(n74 ,n3263 ,n73);
    or g3089(n73 ,n70 ,n72);
    nor g3090(n72 ,n69 ,n24[1]);
    nor g3091(n71 ,n68 ,n3264);
    not g3092(n70 ,n24[0]);
    not g3093(n69 ,n3264);
    not g3094(n68 ,n24[1]);
    nor g3095(n3383 ,n81 ,n84);
    or g3096(n84 ,n76 ,n83);
    or g3097(n83 ,n82 ,n80);
    or g3098(n82 ,n79 ,n75);
    or g3099(n81 ,n77 ,n78);
    nor g3100(n80 ,n46[4] ,n46[3]);
    not g3101(n79 ,n46[9]);
    not g3102(n78 ,n46[5]);
    not g3103(n77 ,n46[6]);
    not g3104(n76 ,n46[7]);
    not g3105(n75 ,n46[8]);
    nor g3106(n3384 ,n91 ,n94);
    or g3107(n94 ,n86 ,n93);
    or g3108(n93 ,n92 ,n90);
    or g3109(n92 ,n89 ,n85);
    or g3110(n91 ,n87 ,n88);
    nor g3111(n90 ,n47[4] ,n47[3]);
    not g3112(n89 ,n47[9]);
    not g3113(n88 ,n47[5]);
    not g3114(n87 ,n47[6]);
    not g3115(n86 ,n47[7]);
    not g3116(n85 ,n47[8]);
    nor g3117(n3385 ,n101 ,n104);
    or g3118(n104 ,n96 ,n103);
    or g3119(n103 ,n102 ,n100);
    or g3120(n102 ,n99 ,n95);
    or g3121(n101 ,n97 ,n98);
    nor g3122(n100 ,n48[4] ,n48[3]);
    not g3123(n99 ,n48[9]);
    not g3124(n98 ,n48[5]);
    not g3125(n97 ,n48[6]);
    not g3126(n96 ,n48[7]);
    not g3127(n95 ,n48[8]);
    nor g3128(n3386 ,n111 ,n114);
    or g3129(n114 ,n106 ,n113);
    or g3130(n113 ,n112 ,n110);
    or g3131(n112 ,n109 ,n105);
    or g3132(n111 ,n107 ,n108);
    nor g3133(n110 ,n49[4] ,n49[3]);
    not g3134(n109 ,n49[9]);
    not g3135(n108 ,n49[5]);
    not g3136(n107 ,n49[6]);
    not g3137(n106 ,n49[7]);
    not g3138(n105 ,n49[8]);
    xor g3139(n3366 ,n50[15] ,n170);
    nor g3140(n3365 ,n169 ,n170);
    nor g3141(n170 ,n126 ,n168);
    nor g3142(n169 ,n50[14] ,n167);
    nor g3143(n3364 ,n166 ,n167);
    not g3144(n168 ,n167);
    nor g3145(n167 ,n116 ,n165);
    nor g3146(n166 ,n50[13] ,n164);
    nor g3147(n3363 ,n163 ,n164);
    not g3148(n165 ,n164);
    nor g3149(n164 ,n129 ,n162);
    nor g3150(n163 ,n50[12] ,n161);
    nor g3151(n3362 ,n160 ,n161);
    not g3152(n162 ,n161);
    nor g3153(n161 ,n125 ,n159);
    nor g3154(n160 ,n50[11] ,n158);
    nor g3155(n3361 ,n157 ,n158);
    not g3156(n159 ,n158);
    nor g3157(n158 ,n127 ,n156);
    nor g3158(n157 ,n50[10] ,n155);
    nor g3159(n3360 ,n154 ,n155);
    not g3160(n156 ,n155);
    nor g3161(n155 ,n124 ,n153);
    nor g3162(n154 ,n50[9] ,n152);
    nor g3163(n3359 ,n151 ,n152);
    not g3164(n153 ,n152);
    nor g3165(n152 ,n121 ,n150);
    nor g3166(n151 ,n50[8] ,n149);
    nor g3167(n3358 ,n148 ,n149);
    not g3168(n150 ,n149);
    nor g3169(n149 ,n122 ,n147);
    nor g3170(n148 ,n50[7] ,n146);
    nor g3171(n3357 ,n145 ,n146);
    not g3172(n147 ,n146);
    nor g3173(n146 ,n115 ,n144);
    nor g3174(n145 ,n50[6] ,n143);
    nor g3175(n3356 ,n142 ,n143);
    not g3176(n144 ,n143);
    nor g3177(n143 ,n120 ,n141);
    nor g3178(n142 ,n50[5] ,n140);
    nor g3179(n3355 ,n139 ,n140);
    not g3180(n141 ,n140);
    nor g3181(n140 ,n118 ,n138);
    nor g3182(n139 ,n50[4] ,n137);
    nor g3183(n3354 ,n136 ,n137);
    not g3184(n138 ,n137);
    nor g3185(n137 ,n117 ,n135);
    nor g3186(n136 ,n50[3] ,n134);
    nor g3187(n3353 ,n133 ,n134);
    not g3188(n135 ,n134);
    nor g3189(n134 ,n119 ,n132);
    nor g3190(n133 ,n50[2] ,n131);
    nor g3191(n3352 ,n131 ,n130);
    not g3192(n132 ,n131);
    nor g3193(n131 ,n123 ,n128);
    nor g3194(n130 ,n50[1] ,n50[0]);
    not g3195(n129 ,n50[12]);
    not g3196(n128 ,n50[0]);
    not g3197(n127 ,n50[10]);
    not g3198(n126 ,n50[14]);
    not g3199(n125 ,n50[11]);
    not g3200(n124 ,n50[9]);
    not g3201(n123 ,n50[1]);
    not g3202(n122 ,n50[7]);
    not g3203(n121 ,n50[8]);
    not g3204(n120 ,n50[5]);
    not g3205(n119 ,n50[2]);
    not g3206(n118 ,n50[4]);
    not g3207(n117 ,n50[3]);
    not g3208(n116 ,n50[13]);
    not g3209(n115 ,n50[6]);
    xor g3210(n3351 ,n51[15] ,n226);
    nor g3211(n3350 ,n225 ,n226);
    nor g3212(n226 ,n182 ,n224);
    nor g3213(n225 ,n51[14] ,n223);
    nor g3214(n3349 ,n222 ,n223);
    not g3215(n224 ,n223);
    nor g3216(n223 ,n172 ,n221);
    nor g3217(n222 ,n51[13] ,n220);
    nor g3218(n3348 ,n219 ,n220);
    not g3219(n221 ,n220);
    nor g3220(n220 ,n185 ,n218);
    nor g3221(n219 ,n51[12] ,n217);
    nor g3222(n3347 ,n216 ,n217);
    not g3223(n218 ,n217);
    nor g3224(n217 ,n181 ,n215);
    nor g3225(n216 ,n51[11] ,n214);
    nor g3226(n3346 ,n213 ,n214);
    not g3227(n215 ,n214);
    nor g3228(n214 ,n183 ,n212);
    nor g3229(n213 ,n51[10] ,n211);
    nor g3230(n3345 ,n210 ,n211);
    not g3231(n212 ,n211);
    nor g3232(n211 ,n180 ,n209);
    nor g3233(n210 ,n51[9] ,n208);
    nor g3234(n3344 ,n207 ,n208);
    not g3235(n209 ,n208);
    nor g3236(n208 ,n177 ,n206);
    nor g3237(n207 ,n51[8] ,n205);
    nor g3238(n3343 ,n204 ,n205);
    not g3239(n206 ,n205);
    nor g3240(n205 ,n178 ,n203);
    nor g3241(n204 ,n51[7] ,n202);
    nor g3242(n3342 ,n201 ,n202);
    not g3243(n203 ,n202);
    nor g3244(n202 ,n171 ,n200);
    nor g3245(n201 ,n51[6] ,n199);
    nor g3246(n3341 ,n198 ,n199);
    not g3247(n200 ,n199);
    nor g3248(n199 ,n176 ,n197);
    nor g3249(n198 ,n51[5] ,n196);
    nor g3250(n3340 ,n195 ,n196);
    not g3251(n197 ,n196);
    nor g3252(n196 ,n174 ,n194);
    nor g3253(n195 ,n51[4] ,n193);
    nor g3254(n3339 ,n192 ,n193);
    not g3255(n194 ,n193);
    nor g3256(n193 ,n173 ,n191);
    nor g3257(n192 ,n51[3] ,n190);
    nor g3258(n3338 ,n189 ,n190);
    not g3259(n191 ,n190);
    nor g3260(n190 ,n175 ,n188);
    nor g3261(n189 ,n51[2] ,n187);
    nor g3262(n3337 ,n187 ,n186);
    not g3263(n188 ,n187);
    nor g3264(n187 ,n179 ,n184);
    nor g3265(n186 ,n51[1] ,n51[0]);
    not g3266(n185 ,n51[12]);
    not g3267(n184 ,n51[0]);
    not g3268(n183 ,n51[10]);
    not g3269(n182 ,n51[14]);
    not g3270(n181 ,n51[11]);
    not g3271(n180 ,n51[9]);
    not g3272(n179 ,n51[1]);
    not g3273(n178 ,n51[7]);
    not g3274(n177 ,n51[8]);
    not g3275(n176 ,n51[5]);
    not g3276(n175 ,n51[2]);
    not g3277(n174 ,n51[4]);
    not g3278(n173 ,n51[3]);
    not g3279(n172 ,n51[13]);
    not g3280(n171 ,n51[6]);
    xor g3281(n3336 ,n52[15] ,n282);
    nor g3282(n3335 ,n281 ,n282);
    nor g3283(n282 ,n238 ,n280);
    nor g3284(n281 ,n52[14] ,n279);
    nor g3285(n3334 ,n278 ,n279);
    not g3286(n280 ,n279);
    nor g3287(n279 ,n228 ,n277);
    nor g3288(n278 ,n52[13] ,n276);
    nor g3289(n3333 ,n275 ,n276);
    not g3290(n277 ,n276);
    nor g3291(n276 ,n241 ,n274);
    nor g3292(n275 ,n52[12] ,n273);
    nor g3293(n3332 ,n272 ,n273);
    not g3294(n274 ,n273);
    nor g3295(n273 ,n237 ,n271);
    nor g3296(n272 ,n52[11] ,n270);
    nor g3297(n3331 ,n269 ,n270);
    not g3298(n271 ,n270);
    nor g3299(n270 ,n239 ,n268);
    nor g3300(n269 ,n52[10] ,n267);
    nor g3301(n3330 ,n266 ,n267);
    not g3302(n268 ,n267);
    nor g3303(n267 ,n236 ,n265);
    nor g3304(n266 ,n52[9] ,n264);
    nor g3305(n3329 ,n263 ,n264);
    not g3306(n265 ,n264);
    nor g3307(n264 ,n233 ,n262);
    nor g3308(n263 ,n52[8] ,n261);
    nor g3309(n3328 ,n260 ,n261);
    not g3310(n262 ,n261);
    nor g3311(n261 ,n234 ,n259);
    nor g3312(n260 ,n52[7] ,n258);
    nor g3313(n3327 ,n257 ,n258);
    not g3314(n259 ,n258);
    nor g3315(n258 ,n227 ,n256);
    nor g3316(n257 ,n52[6] ,n255);
    nor g3317(n3326 ,n254 ,n255);
    not g3318(n256 ,n255);
    nor g3319(n255 ,n232 ,n253);
    nor g3320(n254 ,n52[5] ,n252);
    nor g3321(n3325 ,n251 ,n252);
    not g3322(n253 ,n252);
    nor g3323(n252 ,n230 ,n250);
    nor g3324(n251 ,n52[4] ,n249);
    nor g3325(n3324 ,n248 ,n249);
    not g3326(n250 ,n249);
    nor g3327(n249 ,n229 ,n247);
    nor g3328(n248 ,n52[3] ,n246);
    nor g3329(n3323 ,n245 ,n246);
    not g3330(n247 ,n246);
    nor g3331(n246 ,n231 ,n244);
    nor g3332(n245 ,n52[2] ,n243);
    nor g3333(n3322 ,n243 ,n242);
    not g3334(n244 ,n243);
    nor g3335(n243 ,n235 ,n240);
    nor g3336(n242 ,n52[1] ,n52[0]);
    not g3337(n241 ,n52[12]);
    not g3338(n240 ,n52[0]);
    not g3339(n239 ,n52[10]);
    not g3340(n238 ,n52[14]);
    not g3341(n237 ,n52[11]);
    not g3342(n236 ,n52[9]);
    not g3343(n235 ,n52[1]);
    not g3344(n234 ,n52[7]);
    not g3345(n233 ,n52[8]);
    not g3346(n232 ,n52[5]);
    not g3347(n231 ,n52[2]);
    not g3348(n230 ,n52[4]);
    not g3349(n229 ,n52[3]);
    not g3350(n228 ,n52[13]);
    not g3351(n227 ,n52[6]);
    xor g3352(n3321 ,n53[15] ,n338);
    nor g3353(n3320 ,n337 ,n338);
    nor g3354(n338 ,n294 ,n336);
    nor g3355(n337 ,n53[14] ,n335);
    nor g3356(n3319 ,n334 ,n335);
    not g3357(n336 ,n335);
    nor g3358(n335 ,n284 ,n333);
    nor g3359(n334 ,n53[13] ,n332);
    nor g3360(n3318 ,n331 ,n332);
    not g3361(n333 ,n332);
    nor g3362(n332 ,n297 ,n330);
    nor g3363(n331 ,n53[12] ,n329);
    nor g3364(n3317 ,n328 ,n329);
    not g3365(n330 ,n329);
    nor g3366(n329 ,n293 ,n327);
    nor g3367(n328 ,n53[11] ,n326);
    nor g3368(n3316 ,n325 ,n326);
    not g3369(n327 ,n326);
    nor g3370(n326 ,n295 ,n324);
    nor g3371(n325 ,n53[10] ,n323);
    nor g3372(n3315 ,n322 ,n323);
    not g3373(n324 ,n323);
    nor g3374(n323 ,n292 ,n321);
    nor g3375(n322 ,n53[9] ,n320);
    nor g3376(n3314 ,n319 ,n320);
    not g3377(n321 ,n320);
    nor g3378(n320 ,n289 ,n318);
    nor g3379(n319 ,n53[8] ,n317);
    nor g3380(n3313 ,n316 ,n317);
    not g3381(n318 ,n317);
    nor g3382(n317 ,n290 ,n315);
    nor g3383(n316 ,n53[7] ,n314);
    nor g3384(n3312 ,n313 ,n314);
    not g3385(n315 ,n314);
    nor g3386(n314 ,n283 ,n312);
    nor g3387(n313 ,n53[6] ,n311);
    nor g3388(n3311 ,n310 ,n311);
    not g3389(n312 ,n311);
    nor g3390(n311 ,n288 ,n309);
    nor g3391(n310 ,n53[5] ,n308);
    nor g3392(n3310 ,n307 ,n308);
    not g3393(n309 ,n308);
    nor g3394(n308 ,n286 ,n306);
    nor g3395(n307 ,n53[4] ,n305);
    nor g3396(n3309 ,n304 ,n305);
    not g3397(n306 ,n305);
    nor g3398(n305 ,n285 ,n303);
    nor g3399(n304 ,n53[3] ,n302);
    nor g3400(n3308 ,n301 ,n302);
    not g3401(n303 ,n302);
    nor g3402(n302 ,n287 ,n300);
    nor g3403(n301 ,n53[2] ,n299);
    nor g3404(n3307 ,n299 ,n298);
    not g3405(n300 ,n299);
    nor g3406(n299 ,n291 ,n296);
    nor g3407(n298 ,n53[1] ,n53[0]);
    not g3408(n297 ,n53[12]);
    not g3409(n296 ,n53[0]);
    not g3410(n295 ,n53[10]);
    not g3411(n294 ,n53[14]);
    not g3412(n293 ,n53[11]);
    not g3413(n292 ,n53[9]);
    not g3414(n291 ,n53[1]);
    not g3415(n290 ,n53[7]);
    not g3416(n289 ,n53[8]);
    not g3417(n288 ,n53[5]);
    not g3418(n287 ,n53[2]);
    not g3419(n286 ,n53[4]);
    not g3420(n285 ,n53[3]);
    not g3421(n284 ,n53[13]);
    not g3422(n283 ,n53[6]);
    xor g3423(n3306 ,n46[9] ,n370);
    nor g3424(n3305 ,n369 ,n370);
    nor g3425(n370 ,n345 ,n368);
    nor g3426(n369 ,n46[8] ,n367);
    nor g3427(n3304 ,n366 ,n367);
    not g3428(n368 ,n367);
    nor g3429(n367 ,n341 ,n365);
    nor g3430(n366 ,n46[7] ,n364);
    nor g3431(n3303 ,n363 ,n364);
    not g3432(n365 ,n364);
    nor g3433(n364 ,n342 ,n362);
    nor g3434(n363 ,n46[6] ,n361);
    nor g3435(n3302 ,n360 ,n361);
    not g3436(n362 ,n361);
    nor g3437(n361 ,n339 ,n359);
    nor g3438(n360 ,n46[5] ,n358);
    nor g3439(n3301 ,n357 ,n358);
    not g3440(n359 ,n358);
    nor g3441(n358 ,n346 ,n356);
    nor g3442(n357 ,n46[4] ,n355);
    nor g3443(n3300 ,n354 ,n355);
    not g3444(n356 ,n355);
    nor g3445(n355 ,n347 ,n353);
    nor g3446(n354 ,n46[3] ,n352);
    nor g3447(n3299 ,n351 ,n352);
    not g3448(n353 ,n352);
    nor g3449(n352 ,n340 ,n350);
    nor g3450(n351 ,n46[2] ,n349);
    nor g3451(n3298 ,n349 ,n348);
    not g3452(n350 ,n349);
    nor g3453(n349 ,n343 ,n344);
    nor g3454(n348 ,n46[1] ,n46[0]);
    not g3455(n347 ,n46[3]);
    not g3456(n346 ,n46[4]);
    not g3457(n345 ,n46[8]);
    not g3458(n344 ,n46[0]);
    not g3459(n343 ,n46[1]);
    not g3460(n342 ,n46[6]);
    not g3461(n341 ,n46[7]);
    not g3462(n340 ,n46[2]);
    not g3463(n339 ,n46[5]);
    xor g3464(n3297 ,n47[9] ,n402);
    nor g3465(n3296 ,n401 ,n402);
    nor g3466(n402 ,n377 ,n400);
    nor g3467(n401 ,n47[8] ,n399);
    nor g3468(n3295 ,n398 ,n399);
    not g3469(n400 ,n399);
    nor g3470(n399 ,n373 ,n397);
    nor g3471(n398 ,n47[7] ,n396);
    nor g3472(n3294 ,n395 ,n396);
    not g3473(n397 ,n396);
    nor g3474(n396 ,n374 ,n394);
    nor g3475(n395 ,n47[6] ,n393);
    nor g3476(n3293 ,n392 ,n393);
    not g3477(n394 ,n393);
    nor g3478(n393 ,n371 ,n391);
    nor g3479(n392 ,n47[5] ,n390);
    nor g3480(n3292 ,n389 ,n390);
    not g3481(n391 ,n390);
    nor g3482(n390 ,n378 ,n388);
    nor g3483(n389 ,n47[4] ,n387);
    nor g3484(n3291 ,n386 ,n387);
    not g3485(n388 ,n387);
    nor g3486(n387 ,n379 ,n385);
    nor g3487(n386 ,n47[3] ,n384);
    nor g3488(n3290 ,n383 ,n384);
    not g3489(n385 ,n384);
    nor g3490(n384 ,n372 ,n382);
    nor g3491(n383 ,n47[2] ,n381);
    nor g3492(n3289 ,n381 ,n380);
    not g3493(n382 ,n381);
    nor g3494(n381 ,n375 ,n376);
    nor g3495(n380 ,n47[1] ,n47[0]);
    not g3496(n379 ,n47[3]);
    not g3497(n378 ,n47[4]);
    not g3498(n377 ,n47[8]);
    not g3499(n376 ,n47[0]);
    not g3500(n375 ,n47[1]);
    not g3501(n374 ,n47[6]);
    not g3502(n373 ,n47[7]);
    not g3503(n372 ,n47[2]);
    not g3504(n371 ,n47[5]);
    xor g3505(n3288 ,n48[9] ,n434);
    nor g3506(n3287 ,n433 ,n434);
    nor g3507(n434 ,n409 ,n432);
    nor g3508(n433 ,n48[8] ,n431);
    nor g3509(n3286 ,n430 ,n431);
    not g3510(n432 ,n431);
    nor g3511(n431 ,n405 ,n429);
    nor g3512(n430 ,n48[7] ,n428);
    nor g3513(n3285 ,n427 ,n428);
    not g3514(n429 ,n428);
    nor g3515(n428 ,n406 ,n426);
    nor g3516(n427 ,n48[6] ,n425);
    nor g3517(n3284 ,n424 ,n425);
    not g3518(n426 ,n425);
    nor g3519(n425 ,n403 ,n423);
    nor g3520(n424 ,n48[5] ,n422);
    nor g3521(n3283 ,n421 ,n422);
    not g3522(n423 ,n422);
    nor g3523(n422 ,n410 ,n420);
    nor g3524(n421 ,n48[4] ,n419);
    nor g3525(n3282 ,n418 ,n419);
    not g3526(n420 ,n419);
    nor g3527(n419 ,n411 ,n417);
    nor g3528(n418 ,n48[3] ,n416);
    nor g3529(n3281 ,n415 ,n416);
    not g3530(n417 ,n416);
    nor g3531(n416 ,n404 ,n414);
    nor g3532(n415 ,n48[2] ,n413);
    nor g3533(n3280 ,n413 ,n412);
    not g3534(n414 ,n413);
    nor g3535(n413 ,n407 ,n408);
    nor g3536(n412 ,n48[1] ,n48[0]);
    not g3537(n411 ,n48[3]);
    not g3538(n410 ,n48[4]);
    not g3539(n409 ,n48[8]);
    not g3540(n408 ,n48[0]);
    not g3541(n407 ,n48[1]);
    not g3542(n406 ,n48[6]);
    not g3543(n405 ,n48[7]);
    not g3544(n404 ,n48[2]);
    not g3545(n403 ,n48[5]);
    xor g3546(n3279 ,n49[9] ,n466);
    nor g3547(n3278 ,n465 ,n466);
    nor g3548(n466 ,n441 ,n464);
    nor g3549(n465 ,n49[8] ,n463);
    nor g3550(n3277 ,n462 ,n463);
    not g3551(n464 ,n463);
    nor g3552(n463 ,n437 ,n461);
    nor g3553(n462 ,n49[7] ,n460);
    nor g3554(n3276 ,n459 ,n460);
    not g3555(n461 ,n460);
    nor g3556(n460 ,n438 ,n458);
    nor g3557(n459 ,n49[6] ,n457);
    nor g3558(n3275 ,n456 ,n457);
    not g3559(n458 ,n457);
    nor g3560(n457 ,n435 ,n455);
    nor g3561(n456 ,n49[5] ,n454);
    nor g3562(n3274 ,n453 ,n454);
    not g3563(n455 ,n454);
    nor g3564(n454 ,n442 ,n452);
    nor g3565(n453 ,n49[4] ,n451);
    nor g3566(n3273 ,n450 ,n451);
    not g3567(n452 ,n451);
    nor g3568(n451 ,n443 ,n449);
    nor g3569(n450 ,n49[3] ,n448);
    nor g3570(n3272 ,n447 ,n448);
    not g3571(n449 ,n448);
    nor g3572(n448 ,n436 ,n446);
    nor g3573(n447 ,n49[2] ,n445);
    nor g3574(n3271 ,n445 ,n444);
    not g3575(n446 ,n445);
    nor g3576(n445 ,n439 ,n440);
    nor g3577(n444 ,n49[1] ,n49[0]);
    not g3578(n443 ,n49[3]);
    not g3579(n442 ,n49[4]);
    not g3580(n441 ,n49[8]);
    not g3581(n440 ,n49[0]);
    not g3582(n439 ,n49[1]);
    not g3583(n438 ,n49[6]);
    not g3584(n437 ,n49[7]);
    not g3585(n436 ,n49[2]);
    not g3586(n435 ,n49[5]);
    xor g3587(n3368 ,n34[15] ,n522);
    nor g3588(n3369 ,n521 ,n522);
    nor g3589(n522 ,n478 ,n520);
    nor g3590(n521 ,n34[14] ,n519);
    nor g3591(n3370 ,n518 ,n519);
    not g3592(n520 ,n519);
    nor g3593(n519 ,n468 ,n517);
    nor g3594(n518 ,n34[13] ,n516);
    nor g3595(n3371 ,n515 ,n516);
    not g3596(n517 ,n516);
    nor g3597(n516 ,n481 ,n514);
    nor g3598(n515 ,n34[12] ,n513);
    nor g3599(n3372 ,n512 ,n513);
    not g3600(n514 ,n513);
    nor g3601(n513 ,n477 ,n511);
    nor g3602(n512 ,n34[11] ,n510);
    nor g3603(n3373 ,n509 ,n510);
    not g3604(n511 ,n510);
    nor g3605(n510 ,n479 ,n508);
    nor g3606(n509 ,n34[10] ,n507);
    nor g3607(n3374 ,n506 ,n507);
    not g3608(n508 ,n507);
    nor g3609(n507 ,n476 ,n505);
    nor g3610(n506 ,n34[9] ,n504);
    nor g3611(n3375 ,n503 ,n504);
    not g3612(n505 ,n504);
    nor g3613(n504 ,n473 ,n502);
    nor g3614(n503 ,n34[8] ,n501);
    nor g3615(n3376 ,n500 ,n501);
    not g3616(n502 ,n501);
    nor g3617(n501 ,n474 ,n499);
    nor g3618(n500 ,n34[7] ,n498);
    nor g3619(n3377 ,n497 ,n498);
    not g3620(n499 ,n498);
    nor g3621(n498 ,n467 ,n496);
    nor g3622(n497 ,n34[6] ,n495);
    nor g3623(n3378 ,n494 ,n495);
    not g3624(n496 ,n495);
    nor g3625(n495 ,n472 ,n493);
    nor g3626(n494 ,n34[5] ,n492);
    nor g3627(n3379 ,n491 ,n492);
    not g3628(n493 ,n492);
    nor g3629(n492 ,n470 ,n490);
    nor g3630(n491 ,n34[4] ,n489);
    nor g3631(n3380 ,n488 ,n489);
    not g3632(n490 ,n489);
    nor g3633(n489 ,n469 ,n487);
    nor g3634(n488 ,n34[3] ,n486);
    nor g3635(n3381 ,n485 ,n486);
    not g3636(n487 ,n486);
    nor g3637(n486 ,n471 ,n484);
    nor g3638(n485 ,n34[2] ,n483);
    nor g3639(n3382 ,n483 ,n482);
    not g3640(n484 ,n483);
    nor g3641(n483 ,n475 ,n480);
    nor g3642(n482 ,n34[1] ,n34[0]);
    not g3643(n481 ,n34[12]);
    not g3644(n480 ,n34[0]);
    not g3645(n479 ,n34[10]);
    not g3646(n478 ,n34[14]);
    not g3647(n477 ,n34[11]);
    not g3648(n476 ,n34[9]);
    not g3649(n475 ,n34[1]);
    not g3650(n474 ,n34[7]);
    not g3651(n473 ,n34[8]);
    not g3652(n472 ,n34[5]);
    not g3653(n471 ,n34[2]);
    not g3654(n470 ,n34[4]);
    not g3655(n469 ,n34[3]);
    not g3656(n468 ,n34[13]);
    not g3657(n467 ,n34[6]);
    buf g3658(n3252 ,n3270);
endmodule
