module top (n0, n1, n3, n4, n5, n6, n8, n9, n2, n7, n10, n11, n12, n13, n14, n15, n16, n17);
    input n0, n1, n2;
    input [31:0] n3, n4, n5;
    input [3:0] n6, n7;
    input [1:0] n8;
    input [7:0] n9;
    output [3:0] n10;
    output [31:0] n11, n12, n13, n14;
    output [15:0] n15, n16;
    output [7:0] n17;
    wire n0, n1, n2;
    wire [31:0] n3, n4, n5;
    wire [3:0] n6, n7;
    wire [1:0] n8;
    wire [7:0] n9;
    wire [3:0] n10;
    wire [31:0] n11, n12, n13, n14;
    wire [15:0] n15, n16;
    wire [7:0] n17;
    wire [1:0] n18;
    wire [31:0] n19;
    wire [31:0] n20;
    wire [31:0] n21;
    wire [7:0] n22;
    wire [3:0] n23;
    wire [31:0] n24;
    wire [31:0] n25;
    wire [31:0] n26;
    wire [3:0] n27;
    wire [31:0] n28;
    wire [31:0] n29;
    wire [31:0] n30;
    wire [31:0] n31;
    wire [31:0] n32;
    wire [31:0] n33;
    wire [31:0] n34;
    wire [31:0] n35;
    wire [3:0] n36;
    wire n37, n38, n39, n40, n41, n42, n43, n44;
    wire n45, n46, n47, n48, n49, n50, n51, n52;
    wire n53, n54, n55, n56, n57, n58, n59, n60;
    wire n61, n62, n63, n64, n65, n66, n67, n68;
    wire n69, n70, n71, n72, n73, n74, n75, n76;
    wire n77, n78, n79, n80, n81, n82, n83, n84;
    wire n85, n86, n87, n88, n89, n90, n91, n92;
    wire n93, n94, n95, n96, n97, n98, n99, n100;
    wire n101, n102, n103, n104, n105, n106, n107, n108;
    wire n109, n110, n111, n112, n113, n114, n115, n116;
    wire n117, n118, n119, n120, n121, n122, n123, n124;
    wire n125, n126, n127, n128, n129, n130, n131, n132;
    wire n133, n134, n135, n136, n137, n138, n139, n140;
    wire n141, n142, n143, n144, n145, n146, n147, n148;
    wire n149, n150, n151, n152, n153, n154, n155, n156;
    wire n157, n158, n159, n160, n161, n162, n163, n164;
    wire n165, n166, n167, n168, n169, n170, n171, n172;
    wire n173, n174, n175, n176, n177, n178, n179, n180;
    wire n181, n182, n183, n184, n185, n186, n187, n188;
    wire n189, n190, n191, n192, n193, n194, n195, n196;
    wire n197, n198, n199, n200, n201, n202, n203, n204;
    wire n205, n206, n207, n208, n209, n210, n211, n212;
    wire n213, n214, n215, n216, n217, n218, n219, n220;
    wire n221, n222, n223, n224, n225, n226, n227, n228;
    wire n229, n230, n231, n232, n233, n234, n235, n236;
    wire n237, n238, n239, n240, n241, n242, n243, n244;
    wire n245, n246, n247, n248, n249, n250, n251, n252;
    wire n253, n254, n255, n256, n257, n258, n259, n260;
    wire n261, n262, n263, n264, n265, n266, n267, n268;
    wire n269, n270, n271, n272, n273, n274, n275, n276;
    wire n277, n278, n279, n280, n281, n282, n283, n284;
    wire n285, n286, n287, n288, n289, n290, n291, n292;
    wire n293, n294, n295, n296, n297, n298, n299, n300;
    wire n301, n302, n303, n304, n305, n306, n307, n308;
    wire n309, n310, n311, n312, n313, n314, n315, n316;
    wire n317, n318, n319, n320, n321, n322, n323, n324;
    wire n325, n326, n327, n328, n329, n330, n331, n332;
    wire n333, n334, n335, n336, n337, n338, n339, n340;
    wire n341, n342, n343, n344, n345, n346, n347, n348;
    wire n349, n350, n351, n352, n353, n354, n355, n356;
    wire n357, n358, n359, n360, n361, n362, n363, n364;
    wire n365, n366, n367, n368, n369, n370, n371, n372;
    wire n373, n374, n375, n376, n377, n378, n379, n380;
    wire n381, n382, n383, n384, n385, n386, n387, n388;
    wire n389, n390, n391, n392, n393, n394, n395, n396;
    wire n397, n398, n399, n400, n401, n402, n403, n404;
    wire n405, n406, n407, n408, n409, n410, n411, n412;
    wire n413, n414, n415, n416, n417, n418, n419, n420;
    wire n421, n422, n423, n424, n425, n426, n427, n428;
    wire n429, n430, n431, n432, n433, n434, n435, n436;
    wire n437, n438, n439, n440, n441, n442, n443, n444;
    wire n445, n446, n447, n448, n449, n450, n451, n452;
    wire n453, n454, n455, n456, n457, n458, n459, n460;
    wire n461, n462, n463, n464, n465, n466, n467, n468;
    wire n469, n470, n471, n472, n473, n474, n475, n476;
    wire n477, n478, n479, n480, n481, n482, n483, n484;
    wire n485, n486, n487, n488, n489, n490, n491, n492;
    wire n493, n494, n495, n496, n497, n498, n499, n500;
    wire n501, n502, n503, n504, n505, n506, n507, n508;
    wire n509, n510, n511, n512, n513, n514, n515, n516;
    wire n517, n518, n519, n520, n521, n522, n523, n524;
    wire n525, n526, n527, n528, n529, n530, n531, n532;
    wire n533, n534, n535, n536, n537, n538, n539, n540;
    wire n541, n542, n543, n544, n545, n546, n547, n548;
    wire n549, n550, n551, n552, n553, n554, n555, n556;
    wire n557, n558, n559, n560, n561, n562, n563, n564;
    wire n565, n566, n567, n568, n569, n570, n571, n572;
    wire n573, n574, n575, n576, n577, n578, n579, n580;
    wire n581, n582, n583, n584, n585, n586, n587, n588;
    wire n589, n590, n591, n592, n593, n594, n595, n596;
    wire n597, n598, n599, n600, n601, n602, n603, n604;
    wire n605, n606, n607, n608, n609, n610, n611, n612;
    wire n613, n614, n615, n616, n617, n618, n619, n620;
    wire n621, n622, n623, n624, n625, n626, n627, n628;
    wire n629, n630, n631, n632, n633, n634, n635, n636;
    wire n637, n638, n639, n640, n641, n642, n643, n644;
    wire n645, n646, n647, n648, n649, n650, n651, n652;
    wire n653, n654, n655, n656, n657, n658, n659, n660;
    wire n661, n662, n663, n664, n665, n666, n667, n668;
    wire n669, n670, n671, n672, n673, n674, n675, n676;
    wire n677, n678, n679, n680, n681, n682, n683, n684;
    wire n685, n686, n687, n688, n689, n690, n691, n692;
    wire n693, n694, n695, n696, n697, n698, n699, n700;
    wire n701, n702, n703, n704, n705, n706, n707, n708;
    wire n709, n710, n711, n712, n713, n714, n715, n716;
    wire n717, n718, n719, n720, n721, n722, n723, n724;
    wire n725, n726, n727, n728, n729, n730, n731, n732;
    wire n733, n734, n735, n736, n737, n738, n739, n740;
    wire n741, n742, n743, n744, n745, n746, n747, n748;
    wire n749, n750, n751, n752, n753, n754, n755, n756;
    wire n757, n758, n759, n760, n761, n762, n763, n764;
    wire n765, n766, n767, n768, n769, n770, n771, n772;
    wire n773, n774, n775, n776, n777, n778, n779, n780;
    wire n781, n782, n783, n784, n785, n786, n787, n788;
    wire n789, n790, n791, n792, n793, n794, n795, n796;
    wire n797, n798, n799, n800, n801, n802, n803, n804;
    wire n805, n806, n807, n808, n809, n810, n811, n812;
    wire n813, n814, n815, n816, n817, n818, n819, n820;
    wire n821, n822, n823, n824, n825, n826, n827, n828;
    wire n829, n830, n831, n832, n833, n834, n835, n836;
    wire n837, n838, n839, n840, n841, n842, n843, n844;
    wire n845, n846, n847, n848, n849, n850, n851, n852;
    wire n853, n854, n855, n856, n857, n858, n859, n860;
    wire n861, n862, n863, n864, n865, n866, n867, n868;
    wire n869, n870, n871, n872, n873, n874, n875, n876;
    wire n877, n878, n879, n880, n881, n882, n883, n884;
    wire n885, n886, n887, n888, n889, n890, n891, n892;
    wire n893, n894, n895, n896, n897, n898, n899, n900;
    wire n901, n902, n903, n904, n905, n906, n907, n908;
    wire n909, n910, n911, n912, n913, n914, n915, n916;
    wire n917, n918, n919, n920, n921, n922, n923, n924;
    wire n925, n926, n927, n928, n929, n930, n931, n932;
    wire n933, n934, n935, n936, n937, n938, n939, n940;
    wire n941, n942, n943, n944, n945, n946, n947, n948;
    wire n949, n950, n951, n952, n953, n954, n955, n956;
    wire n957, n958, n959, n960, n961, n962, n963, n964;
    wire n965, n966, n967, n968, n969, n970, n971, n972;
    wire n973, n974, n975, n976, n977, n978, n979, n980;
    wire n981, n982, n983, n984, n985, n986, n987, n988;
    wire n989, n990, n991, n992, n993, n994, n995, n996;
    wire n997, n998, n999, n1000, n1001, n1002, n1003, n1004;
    wire n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
    wire n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
    wire n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028;
    wire n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
    wire n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
    wire n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
    wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
    wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
    wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084;
    wire n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092;
    wire n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100;
    wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
    wire n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116;
    wire n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124;
    wire n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132;
    wire n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140;
    wire n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
    wire n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156;
    wire n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
    wire n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172;
    wire n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180;
    wire n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188;
    wire n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196;
    wire n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204;
    wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212;
    wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
    wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
    wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
    wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
    wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
    wire n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260;
    wire n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268;
    wire n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276;
    wire n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284;
    wire n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292;
    wire n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300;
    wire n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
    wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
    wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
    wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332;
    wire n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340;
    wire n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348;
    wire n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356;
    wire n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364;
    wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
    wire n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380;
    wire n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388;
    wire n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
    wire n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404;
    wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
    wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
    wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
    wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
    wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
    wire n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452;
    wire n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460;
    wire n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468;
    wire n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476;
    wire n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484;
    wire n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492;
    wire n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500;
    wire n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508;
    wire n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516;
    wire n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524;
    wire n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532;
    wire n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540;
    wire n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548;
    wire n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556;
    wire n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564;
    wire n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572;
    wire n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
    wire n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588;
    wire n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596;
    wire n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604;
    wire n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612;
    wire n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620;
    wire n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628;
    wire n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636;
    wire n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644;
    wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
    wire n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660;
    wire n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668;
    wire n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676;
    wire n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684;
    wire n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692;
    wire n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
    wire n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708;
    wire n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716;
    wire n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724;
    wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
    wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
    wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
    wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
    wire n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764;
    wire n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772;
    wire n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
    wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
    wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
    wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
    wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
    wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
    wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
    wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
    wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
    wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
    wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
    wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
    wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
    wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
    wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
    wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
    wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
    wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
    wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
    wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
    wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
    wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
    wire n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956;
    wire n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964;
    wire n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972;
    wire n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980;
    wire n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
    wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
    wire n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
    wire n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012;
    wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
    wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
    wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
    wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
    wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
    wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
    wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
    wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076;
    wire n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084;
    wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
    wire n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100;
    wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
    wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
    wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
    wire n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
    wire n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;
    wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
    wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
    wire n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164;
    wire n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172;
    wire n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180;
    wire n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188;
    wire n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196;
    wire n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204;
    wire n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
    wire n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220;
    wire n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228;
    wire n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236;
    wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
    wire n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252;
    wire n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260;
    wire n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268;
    wire n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276;
    wire n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284;
    wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
    wire n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300;
    wire n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308;
    wire n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316;
    wire n2317, n2318, n2319, n2320, n2321, n2322;
    not g0(n270 ,n9[4]);
    not g1(n224 ,n13[6]);
    or g2(n1997 ,n1053 ,n1591);
    not g3(n267 ,n4[31]);
    not g4(n497 ,n31[7]);
    or g5(n2101 ,n1429 ,n1625);
    dff g6(.RN(n1), .SN(1'b1), .CK(n0), .D(n2223), .Q(n27[0]));
    not g7(n2249 ,n19[7]);
    nor g8(n1473 ,n553 ,n816);
    not g9(n618 ,n35[21]);
    buf g10(n16[15], 1'b0);
    nor g11(n988 ,n671 ,n69);
    xnor g12(n764 ,n511 ,n86);
    nor g13(n1558 ,n613 ,n45);
    dff g14(.RN(n1), .SN(1'b1), .CK(n0), .D(n1912), .Q(n31[12]));
    dff g15(.RN(n1), .SN(1'b1), .CK(n0), .D(n2145), .Q(n13[31]));
    nor g16(n1291 ,n401 ,n67);
    dff g17(.RN(n1), .SN(1'b1), .CK(n0), .D(n2000), .Q(n30[20]));
    nor g18(n1532 ,n108 ,n45);
    nor g19(n961 ,n707 ,n63);
    dff g20(.RN(n1), .SN(1'b1), .CK(n0), .D(n1977), .Q(n21[26]));
    xnor g21(n668 ,n158 ,n395);
    xnor g22(n789 ,n76 ,n86);
    or g23(n1869 ,n1247 ,n1100);
    nor g24(n1103 ,n93 ,n59);
    not g25(n212 ,n29[23]);
    xnor g26(n710 ,n26[21] ,n33[17]);
    not g27(n258 ,n35[26]);
    xnor g28(n684 ,n550 ,n179);
    not g29(n145 ,n32[15]);
    not g30(n305 ,n4[6]);
    not g31(n294 ,n4[23]);
    xnor g32(n808 ,n26[7] ,n33[3]);
    or g33(n2177 ,n1292 ,n1007);
    or g34(n1889 ,n1267 ,n1107);
    xnor g35(n669 ,n171 ,n481);
    not g36(n527 ,n28[17]);
    nor g37(n1208 ,n478 ,n61);
    dff g38(.RN(n1), .SN(1'b1), .CK(n0), .D(n2022), .Q(n30[14]));
    not g39(n495 ,n29[26]);
    nor g40(n943 ,n685 ,n64);
    nor g41(n1472 ,n618 ,n68);
    dff g42(.RN(n1), .SN(1'b1), .CK(n0), .D(n1789), .Q(n11[7]));
    nor g43(n1096 ,n367 ,n59);
    dff g44(.RN(n1), .SN(1'b1), .CK(n0), .D(n1940), .Q(n35[8]));
    nor g45(n1457 ,n213 ,n43);
    nor g46(n1453 ,n141 ,n50);
    or g47(n1896 ,n1278 ,n1110);
    nor g48(n1188 ,n112 ,n57);
    nor g49(n1626 ,n341 ,n49);
    or g50(n2089 ,n1080 ,n1606);
    or g51(n2293 ,n2280 ,n2264);
    or g52(n2171 ,n1493 ,n1115);
    nor g53(n1160 ,n430 ,n43);
    not g54(n171 ,n34[18]);
    not g55(n493 ,n31[9]);
    xnor g56(n634 ,n534 ,n116);
    nor g57(n853 ,n722 ,n48);
    nor g58(n1728 ,n466 ,n66);
    nor g59(n1074 ,n360 ,n51);
    not g60(n611 ,n35[14]);
    nor g61(n1529 ,n463 ,n48);
    nor g62(n1636 ,n276 ,n52);
    dff g63(.RN(n1), .SN(1'b1), .CK(n0), .D(n1774), .Q(n26[31]));
    not g64(n494 ,n29[27]);
    nor g65(n1216 ,n140 ,n57);
    not g66(n455 ,n26[29]);
    or g67(n2270 ,n2256 ,n24[4]);
    nor g68(n1126 ,n411 ,n43);
    xnor g69(n751 ,n21[15] ,n24[15]);
    nor g70(n1705 ,n145 ,n63);
    dff g71(.RN(n1), .SN(1'b1), .CK(n0), .D(n1760), .Q(n11[28]));
    not g72(n375 ,n21[23]);
    dff g73(.RN(n1), .SN(1'b1), .CK(n0), .D(n2059), .Q(n30[5]));
    dff g74(.RN(n1), .SN(1'b1), .CK(n0), .D(n2109), .Q(n24[17]));
    not g75(n472 ,n29[8]);
    or g76(n2271 ,n2255 ,n19[4]);
    dff g77(.RN(n1), .SN(1'b1), .CK(n0), .D(n2174), .Q(n15[10]));
    nor g78(n1707 ,n448 ,n63);
    dff g79(.RN(n1), .SN(1'b1), .CK(n0), .D(n1786), .Q(n11[10]));
    nor g80(n58 ,n37 ,n41);
    not g81(n94 ,n21[17]);
    xnor g82(n685 ,n195 ,n408);
    xnor g83(n640 ,n26[25] ,n33[21]);
    or g84(n1836 ,n1227 ,n1090);
    dff g85(.RN(n1), .SN(1'b1), .CK(n0), .D(n2184), .Q(n25[28]));
    not g86(n364 ,n21[30]);
    or g87(n1781 ,n1159 ,n1541);
    or g88(n1980 ,n1353 ,n1688);
    nor g89(n1259 ,n189 ,n53);
    nor g90(n1358 ,n196 ,n54);
    not g91(n296 ,n5[13]);
    dff g92(.RN(n1), .SN(1'b1), .CK(n0), .D(n1873), .Q(n28[17]));
    dff g93(.RN(n1), .SN(1'b1), .CK(n0), .D(n2004), .Q(n34[3]));
    not g94(n559 ,n15[9]);
    nor g95(n2205 ,n788 ,n1008);
    nor g96(n1313 ,n207 ,n53);
    nor g97(n1546 ,n449 ,n47);
    or g98(n2309 ,n2298 ,n2293);
    dff g99(.RN(n1), .SN(1'b1), .CK(n0), .D(n2088), .Q(n24[28]));
    or g100(n1803 ,n1187 ,n873);
    nor g101(n1329 ,n537 ,n68);
    dff g102(.RN(n1), .SN(1'b1), .CK(n0), .D(n2060), .Q(n21[12]));
    dff g103(.RN(n1), .SN(1'b1), .CK(n0), .D(n2162), .Q(n29[23]));
    nor g104(n1553 ,n226 ,n48);
    not g105(n2245 ,n20[3]);
    or g106(n1938 ,n1404 ,n1733);
    not g107(n165 ,n35[5]);
    nor g108(n1147 ,n220 ,n44);
    not g109(n402 ,n33[20]);
    buf g110(n17[6], 1'b0);
    nor g111(n955 ,n697 ,n63);
    dff g112(.RN(n1), .SN(1'b1), .CK(n0), .D(n1981), .Q(n26[7]));
    or g113(n1963 ,n1341 ,n1671);
    not g114(n343 ,n5[25]);
    dff g115(.RN(n1), .SN(1'b1), .CK(n0), .D(n1991), .Q(n34[9]));
    or g116(n2151 ,n1470 ,n840);
    dff g117(.RN(n1), .SN(1'b1), .CK(n0), .D(n2025), .Q(n33[25]));
    or g118(n1876 ,n1253 ,n1102);
    not g119(n491 ,n29[21]);
    dff g120(.RN(n1), .SN(1'b1), .CK(n0), .D(n2196), .Q(n15[6]));
    nor g121(n1387 ,n465 ,n51);
    dff g122(.RN(n1), .SN(1'b1), .CK(n0), .D(n1751), .Q(n12[29]));
    not g123(n159 ,n28[5]);
    or g124(n2094 ,n1425 ,n1618);
    not g125(n72 ,n22[3]);
    xnor g126(n771 ,n92 ,n104);
    nor g127(n992 ,n675 ,n69);
    nor g128(n1461 ,n494 ,n61);
    not g129(n344 ,n4[4]);
    or g130(n2202 ,n1414 ,n975);
    dff g131(.RN(n1), .SN(1'b1), .CK(n0), .D(n1810), .Q(n29[4]));
    not g132(n253 ,n13[8]);
    not g133(n2239 ,n21[29]);
    not g134(n544 ,n34[2]);
    not g135(n297 ,n4[3]);
    dff g136(.RN(n1), .SN(1'b1), .CK(n0), .D(n2125), .Q(n29[30]));
    dff g137(.RN(n1), .SN(1'b1), .CK(n0), .D(n1918), .Q(n31[10]));
    nor g138(n1565 ,n618 ,n47);
    or g139(n2033 ,n1140 ,n1565);
    nor g140(n1095 ,n375 ,n60);
    buf g141(n16[5], n15[1]);
    nor g142(n1593 ,n329 ,n49);
    dff g143(.RN(n1), .SN(1'b1), .CK(n0), .D(n2002), .Q(n26[5]));
    not g144(n482 ,n34[7]);
    not g145(n291 ,n5[22]);
    nor g146(n986 ,n669 ,n69);
    dff g147(.RN(n1), .SN(1'b1), .CK(n0), .D(n2113), .Q(n21[3]));
    nor g148(n835 ,n762 ,n47);
    dff g149(.RN(n1), .SN(1'b1), .CK(n0), .D(n1807), .Q(n26[28]));
    dff g150(.RN(n1), .SN(1'b1), .CK(n0), .D(n1932), .Q(n35[14]));
    buf g151(n16[10], n15[6]);
    nor g152(n1084 ,n98 ,n48);
    dff g153(.RN(n1), .SN(1'b1), .CK(n0), .D(n2080), .Q(n10[0]));
    xnor g154(n694 ,n178 ,n431);
    or g155(n2041 ,n1389 ,n1570);
    or g156(n2053 ,n1490 ,n1575);
    nor g157(n1676 ,n112 ,n63);
    nor g158(n1364 ,n441 ,n61);
    dff g159(.RN(n1), .SN(1'b1), .CK(n0), .D(n822), .Q(n17[1]));
    or g160(n2135 ,n1453 ,n1654);
    dff g161(.RN(n1), .SN(1'b1), .CK(n0), .D(n1816), .Q(n26[25]));
    dff g162(.RN(n1), .SN(1'b1), .CK(n0), .D(n1842), .Q(n32[8]));
    not g163(n103 ,n33[11]);
    nor g164(n1414 ,n573 ,n65);
    not g165(n459 ,n24[14]);
    nor g166(n1622 ,n313 ,n49);
    nor g167(n883 ,n742 ,n60);
    dff g168(.RN(n1), .SN(1'b1), .CK(n0), .D(n2108), .Q(n22[1]));
    dff g169(.RN(n1), .SN(1'b1), .CK(n0), .D(n1747), .Q(n15[5]));
    nor g170(n1010 ,n350 ,n818);
    or g171(n2214 ,n1318 ,n2209);
    not g172(n418 ,n24[22]);
    nor g173(n1591 ,n294 ,n49);
    nor g174(n1221 ,n544 ,n53);
    or g175(n2027 ,n1378 ,n1563);
    nor g176(n1391 ,n454 ,n44);
    or g177(n2168 ,n1492 ,n964);
    dff g178(.RN(n1), .SN(1'b1), .CK(n0), .D(n1797), .Q(n29[7]));
    dff g179(.RN(n1), .SN(1'b1), .CK(n0), .D(n1772), .Q(n29[11]));
    dff g180(.RN(n1), .SN(1'b1), .CK(n0), .D(n2031), .Q(n33[22]));
    or g181(n822 ,n17[1] ,n820);
    nor g182(n953 ,n806 ,n63);
    not g183(n530 ,n28[21]);
    not g184(n429 ,n30[26]);
    not g185(n322 ,n4[30]);
    not g186(n498 ,n31[13]);
    xnor g187(n646 ,n494 ,n452);
    or g188(n1915 ,n1301 ,n934);
    not g189(n181 ,n34[6]);
    nor g190(n1253 ,n515 ,n57);
    xnor g191(n20[0] ,n2227 ,n18[0]);
    not g192(n211 ,n35[3]);
    dff g193(.RN(n1), .SN(1'b1), .CK(n0), .D(n2028), .Q(n33[23]));
    or g194(n2083 ,n1421 ,n1609);
    nor g195(n1304 ,n452 ,n61);
    dff g196(.RN(n1), .SN(1'b1), .CK(n0), .D(n2180), .Q(n13[10]));
    nor g197(n1290 ,n159 ,n57);
    nor g198(n1485 ,n595 ,n68);
    nor g199(n1031 ,n77 ,n818);
    or g200(n1921 ,n1302 ,n1003);
    nor g201(n1505 ,n260 ,n816);
    xnor g202(n735 ,n21[29] ,n24[29]);
    not g203(n511 ,n29[0]);
    not g204(n81 ,n21[6]);
    xnor g205(n743 ,n547 ,n368);
    nor g206(n1616 ,n292 ,n52);
    not g207(n197 ,n28[15]);
    dff g208(.RN(n1), .SN(1'b1), .CK(n0), .D(n1757), .Q(n11[29]));
    nor g209(n1352 ,n529 ,n54);
    or g210(n2288 ,n2233 ,n2240);
    or g211(n2055 ,n1400 ,n1576);
    not g212(n421 ,n24[3]);
    nor g213(n1228 ,n420 ,n57);
    nor g214(n829 ,n766 ,n47);
    nor g215(n1337 ,n487 ,n53);
    nor g216(n1100 ,n90 ,n59);
    dff g217(.RN(n1), .SN(1'b1), .CK(n0), .D(n2063), .Q(n30[4]));
    nor g218(n889 ,n747 ,n63);
    dff g219(.RN(n1), .SN(1'b1), .CK(n0), .D(n2096), .Q(n24[24]));
    nor g220(n1637 ,n296 ,n49);
    not g221(n496 ,n34[30]);
    dff g222(.RN(n1), .SN(1'b1), .CK(n0), .D(n1819), .Q(n29[2]));
    not g223(n175 ,n28[18]);
    nor g224(n1195 ,n415 ,n57);
    dff g225(.RN(n1), .SN(1'b1), .CK(n0), .D(n1792), .Q(n26[30]));
    not g226(n448 ,n32[13]);
    dff g227(.RN(n1), .SN(1'b1), .CK(n0), .D(n1990), .Q(n21[24]));
    or g228(n2030 ,n1042 ,n1597);
    or g229(n1873 ,n1249 ,n1101);
    nor g230(n1419 ,n433 ,n51);
    dff g231(.RN(n1), .SN(1'b1), .CK(n0), .D(n2143), .Q(n14[0]));
    not g232(n453 ,n30[12]);
    not g233(n204 ,n28[25]);
    or g234(n1773 ,n1153 ,n1535);
    or g235(n2023 ,n1375 ,n1561);
    nor g236(n1218 ,n448 ,n58);
    or g237(n2077 ,n1412 ,n1120);
    or g238(n1908 ,n1290 ,n1113);
    buf g239(n12[5], n11[5]);
    xnor g240(n680 ,n544 ,n208);
    nor g241(n1500 ,n239 ,n43);
    nor g242(n974 ,n792 ,n66);
    nor g243(n838 ,n761 ,n45);
    not g244(n574 ,n13[16]);
    dff g245(.RN(n1), .SN(1'b1), .CK(n0), .D(n2163), .Q(n13[20]));
    not g246(n503 ,n34[26]);
    dff g247(.RN(n1), .SN(1'b1), .CK(n0), .D(n1848), .Q(n32[5]));
    or g248(n1937 ,n1319 ,n947);
    nor g249(n1471 ,n184 ,n61);
    dff g250(.RN(n1), .SN(1'b1), .CK(n0), .D(n1956), .Q(n34[30]));
    nor g251(n863 ,n802 ,n48);
    nor g252(n1136 ,n249 ,n65);
    dff g253(.RN(n1), .SN(1'b1), .CK(n0), .D(n1935), .Q(n31[6]));
    nor g254(n1540 ,n462 ,n47);
    dff g255(.RN(n1), .SN(1'b1), .CK(n0), .D(n2084), .Q(n22[7]));
    or g256(n1768 ,n1149 ,n1532);
    nor g257(n895 ,n752 ,n60);
    buf g258(n16[11], n15[7]);
    nor g259(n1592 ,n274 ,n49);
    nor g260(n1335 ,n485 ,n54);
    nor g261(n1319 ,n166 ,n53);
    or g262(n2196 ,n1517 ,n1028);
    nor g263(n1132 ,n231 ,n816);
    xor g264(n19[3] ,n21[3] ,n22[3]);
    not g265(n615 ,n11[4]);
    nor g266(n2210 ,n59 ,n1744);
    nor g267(n1675 ,n408 ,n63);
    or g268(n1859 ,n1031 ,n1579);
    not g269(n168 ,n31[26]);
    dff g270(.RN(n1), .SN(1'b1), .CK(n0), .D(n2024), .Q(n30[13]));
    dff g271(.RN(n1), .SN(1'b1), .CK(n0), .D(n1882), .Q(n28[14]));
    nor g272(n1257 ,n405 ,n67);
    dff g273(.RN(n1), .SN(1'b1), .CK(n0), .D(n2128), .Q(n24[4]));
    nor g274(n852 ,n720 ,n47);
    dff g275(.RN(n1), .SN(1'b1), .CK(n0), .D(n1983), .Q(n30[24]));
    nor g276(n832 ,n781 ,n47);
    dff g277(.RN(n1), .SN(1'b1), .CK(n0), .D(n2073), .Q(n33[0]));
    not g278(n371 ,n21[26]);
    nor g279(n2199 ,n173 ,n1282);
    not g280(n463 ,n26[25]);
    or g281(n1968 ,n1342 ,n1676);
    nor g282(n1638 ,n300 ,n49);
    not g283(n342 ,n9[7]);
    buf g284(n16[14], 1'b0);
    nor g285(n914 ,n642 ,n56);
    dff g286(.RN(n1), .SN(1'b1), .CK(n0), .D(n1821), .Q(n32[20]));
    not g287(n276 ,n5[14]);
    nor g288(n869 ,n733 ,n59);
    nor g289(n1235 ,n404 ,n65);
    dff g290(.RN(n1), .SN(1'b1), .CK(n0), .D(n1892), .Q(n28[9]));
    xnor g291(n19[1] ,n2225 ,n18[1]);
    dff g292(.RN(n1), .SN(1'b1), .CK(n0), .D(n2111), .Q(n22[0]));
    or g293(n1830 ,n1210 ,n1720);
    or g294(n1795 ,n1176 ,n1553);
    dff g295(.RN(n1), .SN(1'b1), .CK(n0), .D(n2112), .Q(n24[15]));
    not g296(n415 ,n32[25]);
    not g297(n535 ,n28[26]);
    or g298(n2068 ,n1070 ,n1602);
    nor g299(n54 ,n38 ,n41);
    nor g300(n1112 ,n81 ,n59);
    nor g301(n1305 ,n493 ,n53);
    nor g302(n1508 ,n558 ,n46);
    not g303(n423 ,n32[11]);
    dff g304(.RN(n1), .SN(1'b1), .CK(n0), .D(n1906), .Q(n35[29]));
    or g305(n1855 ,n1236 ,n1095);
    dff g306(.RN(n1), .SN(1'b1), .CK(n0), .D(n2070), .Q(n26[2]));
    dff g307(.RN(n1), .SN(1'b1), .CK(n0), .D(n2006), .Q(n34[2]));
    nor g308(n1374 ,n131 ,n51);
    not g309(n2246 ,n24[16]);
    not g310(n239 ,n13[12]);
    or g311(n1780 ,n1150 ,n1021);
    dff g312(.RN(n1), .SN(1'b1), .CK(n0), .D(n2136), .Q(n18[1]));
    not g313(n356 ,n21[2]);
    dff g314(.RN(n1), .SN(1'b1), .CK(n0), .D(n2179), .Q(n29[19]));
    xnor g315(n629 ,n185 ,n388);
    xnor g316(n36[2] ,n2322 ,n25[30]);
    dff g317(.RN(n1), .SN(1'b1), .CK(n0), .D(n1825), .Q(n32[17]));
    nor g318(n1263 ,n522 ,n53);
    or g319(n1850 ,n1232 ,n1093);
    nor g320(n1451 ,n139 ,n51);
    nor g321(n957 ,n726 ,n64);
    not g322(n620 ,n11[11]);
    not g323(n454 ,n33[14]);
    or g324(n2088 ,n1394 ,n1612);
    or g325(n2280 ,n2258 ,n24[29]);
    not g326(n213 ,n14[1]);
    or g327(n2218 ,n70 ,n2211);
    xnor g328(n716 ,n26[22] ,n33[18]);
    nor g329(n902 ,n767 ,n59);
    dff g330(.RN(n1), .SN(1'b1), .CK(n0), .D(n2046), .Q(n33[14]));
    dff g331(.RN(n1), .SN(1'b1), .CK(n0), .D(n2016), .Q(n33[30]));
    nor g332(n926 ,n656 ,n56);
    or g333(n1949 ,n1317 ,n1734);
    or g334(n1901 ,n1285 ,n1112);
    dff g335(.RN(n1), .SN(1'b1), .CK(n0), .D(n1843), .Q(n28[27]));
    dff g336(.RN(n1), .SN(1'b1), .CK(n0), .D(n1845), .Q(n26[20]));
    not g337(n283 ,n4[25]);
    nor g338(n1247 ,n175 ,n57);
    or g339(n2215 ,n1324 ,n2210);
    not g340(n447 ,n33[17]);
    or g341(n1961 ,n1336 ,n1672);
    nor g342(n1502 ,n559 ,n65);
    nor g343(n1431 ,n460 ,n50);
    dff g344(.RN(n1), .SN(1'b1), .CK(n0), .D(n1874), .Q(n26[17]));
    not g345(n474 ,n28[12]);
    xnor g346(n749 ,n21[17] ,n24[17]);
    nor g347(n1171 ,n216 ,n43);
    dff g348(.RN(n1), .SN(1'b1), .CK(n0), .D(n1926), .Q(n35[17]));
    buf g349(n12[4], n11[4]);
    buf g350(n14[19], n11[19]);
    or g351(n1916 ,n1459 ,n982);
    nor g352(n1038 ,n355 ,n50);
    dff g353(.RN(n1), .SN(1'b1), .CK(n0), .D(n2107), .Q(n24[18]));
    dff g354(.RN(n1), .SN(1'b1), .CK(n0), .D(n1791), .Q(n11[6]));
    dff g355(.RN(n1), .SN(1'b1), .CK(n0), .D(n1885), .Q(n31[22]));
    dff g356(.RN(n1), .SN(1'b1), .CK(n0), .D(n2062), .Q(n33[5]));
    nor g357(n1435 ,n459 ,n818);
    nor g358(n1417 ,n560 ,n819);
    nor g359(n1004 ,n631 ,n69);
    buf g360(n14[18], n11[18]);
    or g361(n1874 ,n1257 ,n1727);
    buf g362(n14[6], n11[30]);
    not g363(n109 ,n32[26]);
    dff g364(.RN(n1), .SN(1'b1), .CK(n0), .D(n1958), .Q(n21[30]));
    nor g365(n1121 ,n98 ,n69);
    or g366(n1943 ,n1325 ,n993);
    not g367(n127 ,n32[31]);
    or g368(n2130 ,n1449 ,n1650);
    not g369(n146 ,n24[13]);
    nor g370(n1678 ,n456 ,n55);
    or g371(n1785 ,n1163 ,n1544);
    not g372(n614 ,n13[15]);
    not g373(n293 ,n5[3]);
    not g374(n422 ,n32[27]);
    not g375(n538 ,n28[27]);
    xnor g376(n807 ,n485 ,n523);
    nor g377(n1486 ,n539 ,n62);
    xnor g378(n774 ,n21[26] ,n24[26]);
    not g379(n164 ,n31[30]);
    or g380(n1845 ,n1235 ,n1724);
    nor g381(n843 ,n708 ,n47);
    not g382(n2204 ,n2203);
    nor g383(n1401 ,n142 ,n44);
    not g384(n336 ,n4[15]);
    not g385(n416 ,n30[17]);
    not g386(n316 ,n5[27]);
    nor g387(n1317 ,n449 ,n67);
    not g388(n384 ,n32[7]);
    not g389(n124 ,n32[17]);
    nor g390(n1653 ,n317 ,n49);
    not g391(n540 ,n29[2]);
    dff g392(.RN(n1), .SN(1'b1), .CK(n0), .D(n2182), .Q(n13[9]));
    xnor g393(n647 ,n495 ,n429);
    dff g394(.RN(n1), .SN(1'b1), .CK(n0), .D(n2181), .Q(n15[9]));
    not g395(n272 ,n9[5]);
    nor g396(n1093 ,n358 ,n59);
    xnor g397(n802 ,n26[6] ,n33[2]);
    or g398(n2015 ,n1064 ,n1594);
    or g399(n1835 ,n1222 ,n899);
    nor g400(n1617 ,n270 ,n49);
    nor g401(n1361 ,n211 ,n68);
    dff g402(.RN(n1), .SN(1'b1), .CK(n0), .D(n1857), .Q(n28[22]));
    nor g403(n1017 ,n349 ,n47);
    dff g404(.RN(n1), .SN(1'b1), .CK(n0), .D(n1830), .Q(n26[24]));
    not g405(n571 ,n13[27]);
    or g406(n2159 ,n1478 ,n844);
    nor g407(n1397 ,n450 ,n61);
    dff g408(.RN(n1), .SN(1'b1), .CK(n0), .D(n2021), .Q(n33[27]));
    nor g409(n1564 ,n215 ,n45);
    buf g410(n12[24], n11[24]);
    dff g411(.RN(n1), .SN(1'b1), .CK(n0), .D(n1934), .Q(n35[12]));
    or g412(n2029 ,n1379 ,n1661);
    or g413(n1770 ,n1146 ,n1020);
    dff g414(.RN(n1), .SN(1'b1), .CK(n0), .D(n2121), .Q(n24[10]));
    nor g415(n848 ,n693 ,n45);
    xnor g416(n803 ,n350 ,n370);
    nor g417(n1735 ,n101 ,n66);
    dff g418(.RN(n1), .SN(1'b1), .CK(n0), .D(n2066), .Q(n33[3]));
    nor g419(n1026 ,n73 ,n66);
    nor g420(n1647 ,n281 ,n52);
    dff g421(.RN(n1), .SN(1'b1), .CK(n0), .D(n1779), .Q(n29[10]));
    nor g422(n975 ,n793 ,n66);
    nor g423(n1580 ,n287 ,n817);
    not g424(n335 ,n5[16]);
    dff g425(.RN(n1), .SN(1'b1), .CK(n0), .D(n1853), .Q(n32[3]));
    dff g426(.RN(n1), .SN(1'b1), .CK(n0), .D(n2035), .Q(n30[10]));
    dff g427(.RN(n1), .SN(1'b1), .CK(n0), .D(n2187), .Q(n29[17]));
    nor g428(n1523 ,n385 ,n48);
    not g429(n573 ,n26[1]);
    not g430(n458 ,n26[19]);
    not g431(n334 ,n5[9]);
    nor g432(n1143 ,n555 ,n46);
    xnor g433(n679 ,n26[13] ,n33[9]);
    not g434(n369 ,n21[8]);
    nor g435(n1528 ,n107 ,n45);
    not g436(n299 ,n4[0]);
    nor g437(n1338 ,n503 ,n54);
    nor g438(n1201 ,n396 ,n58);
    not g439(n2259 ,n21[10]);
    dff g440(.RN(n1), .SN(1'b1), .CK(n0), .D(n2072), .Q(n30[2]));
    not g441(n288 ,n5[10]);
    not g442(n394 ,n24[10]);
    nor g443(n1741 ,n103 ,n66);
    xnor g444(n796 ,n74 ,n362);
    nor g445(n1288 ,n613 ,n819);
    buf g446(n14[25], n11[25]);
    not g447(n499 ,n28[0]);
    dff g448(.RN(n1), .SN(1'b1), .CK(n0), .D(n1752), .Q(n29[14]));
    nor g449(n1217 ,n209 ,n57);
    nor g450(n1116 ,n82 ,n66);
    nor g451(n1354 ,n203 ,n53);
    nor g452(n1377 ,n152 ,n62);
    nor g453(n1721 ,n102 ,n66);
    or g454(n2004 ,n1233 ,n903);
    not g455(n537 ,n35[2]);
    or g456(n1778 ,n1158 ,n1540);
    nor g457(n1054 ,n380 ,n818);
    or g458(n2301 ,n2260 ,n2273);
    xor g459(n19[5] ,n21[5] ,n22[5]);
    dff g460(.RN(n1), .SN(1'b1), .CK(n0), .D(n1809), .Q(n32[26]));
    or g461(n1987 ,n1060 ,n1589);
    nor g462(n1545 ,n446 ,n47);
    nor g463(n1436 ,n146 ,n818);
    nor g464(n1667 ,n109 ,n64);
    not g465(n480 ,n34[5]);
    or g466(n2049 ,n1510 ,n1577);
    or g467(n2152 ,n1471 ,n960);
    not g468(n268 ,n4[7]);
    not g469(n529 ,n34[15]);
    nor g470(n1484 ,n232 ,n43);
    not g471(n214 ,n11[9]);
    not g472(n539 ,n29[22]);
    not g473(n326 ,n9[0]);
    nor g474(n1418 ,n497 ,n53);
    not g475(n432 ,n30[30]);
    nor g476(n1677 ,n403 ,n56);
    nor g477(n1349 ,n585 ,n67);
    nor g478(n1671 ,n438 ,n56);
    nor g479(n1016 ,n348 ,n45);
    or g480(n2098 ,n1426 ,n1621);
    or g481(n2024 ,n1377 ,n1707);
    xnor g482(n650 ,n212 ,n456);
    buf g483(n12[19], n11[19]);
    not g484(n1282 ,n1281);
    dff g485(.RN(n1), .SN(1'b1), .CK(n0), .D(n2085), .Q(n24[29]));
    nor g486(n1205 ,n132 ,n57);
    or g487(n1947 ,n1361 ,n996);
    xnor g488(n658 ,n473 ,n416);
    not g489(n567 ,n35[29]);
    not g490(n392 ,n30[11]);
    nor g491(n1090 ,n97 ,n59);
    buf g492(n14[4], n11[28]);
    not g493(n298 ,n4[8]);
    not g494(n581 ,n11[29]);
    nor g495(n1059 ,n364 ,n51);
    not g496(n556 ,n15[5]);
    nor g497(n1005 ,n639 ,n69);
    dff g498(.RN(n1), .SN(1'b1), .CK(n0), .D(n2191), .Q(n13[5]));
    nor g499(n1189 ,n524 ,n61);
    not g500(n560 ,n10[3]);
    buf g501(n12[2], n11[30]);
    buf g502(n12[26], n11[26]);
    nor g503(n1571 ,n611 ,n47);
    or g504(n2034 ,n1384 ,n1566);
    nor g505(n951 ,n805 ,n64);
    not g506(n512 ,n31[19]);
    xnor g507(n801 ,n516 ,n199);
    nor g508(n827 ,n783 ,n48);
    xnor g509(n2226 ,n21[0] ,n22[0]);
    nor g510(n1480 ,n212 ,n62);
    or g511(n2063 ,n1406 ,n949);
    xnor g512(n663 ,n157 ,n453);
    not g513(n365 ,n21[29]);
    xnor g514(n2225 ,n21[1] ,n22[1]);
    dff g515(.RN(n1), .SN(1'b1), .CK(n0), .D(n1782), .Q(n11[13]));
    nor g516(n1623 ,n291 ,n817);
    nor g517(n1362 ,n147 ,n61);
    nor g518(n1495 ,n614 ,n44);
    nor g519(n1240 ,n458 ,n65);
    nor g520(n1241 ,n475 ,n58);
    dff g521(.RN(n1), .SN(1'b1), .CK(n0), .D(n1787), .Q(n11[9]));
    not g522(n92 ,n36[0]);
    or g523(n2066 ,n1408 ,n833);
    not g524(n596 ,n35[19]);
    not g525(n116 ,n30[4]);
    nor g526(n1149 ,n244 ,n44);
    nor g527(n1302 ,n223 ,n819);
    nor g528(n1610 ,n315 ,n817);
    xnor g529(n699 ,n202 ,n423);
    nor g530(n870 ,n636 ,n63);
    not g531(n280 ,n5[23]);
    or g532(n2078 ,n1413 ,n1121);
    xnor g533(n765 ,n21[6] ,n24[6]);
    dff g534(.RN(n1), .SN(1'b1), .CK(n0), .D(n2087), .Q(n22[6]));
    dff g535(.RN(n1), .SN(1'b1), .CK(n0), .D(n2114), .Q(n24[14]));
    not g536(n388 ,n30[9]);
    not g537(n257 ,n35[9]);
    dff g538(.RN(n1), .SN(1'b1), .CK(n0), .D(n2030), .Q(n21[17]));
    nor g539(n1578 ,n617 ,n45);
    xnor g540(n804 ,n72 ,n357);
    nor g541(n1407 ,n468 ,n816);
    not g542(n247 ,n13[30]);
    not g543(n424 ,n24[9]);
    nor g544(n934 ,n799 ,n60);
    or g545(n1912 ,n1296 ,n931);
    nor g546(n1170 ,n233 ,n43);
    or g547(n2161 ,n1481 ,n846);
    dff g548(.RN(n1), .SN(1'b1), .CK(n0), .D(n1989), .Q(n34[10]));
    dff g549(.RN(n1), .SN(1'b1), .CK(n0), .D(n1827), .Q(n32[15]));
    dff g550(.RN(n1), .SN(1'b1), .CK(n0), .D(n1939), .Q(n35[9]));
    dff g551(.RN(n1), .SN(1'b1), .CK(n0), .D(n2194), .Q(n29[16]));
    or g552(n1771 ,n1152 ,n1534);
    not g553(n467 ,n26[7]);
    dff g554(.RN(n1), .SN(1'b1), .CK(n0), .D(n1858), .Q(n32[0]));
    nor g555(n1685 ,n416 ,n56);
    nor g556(n1309 ,n575 ,n68);
    or g557(n2155 ,n1473 ,n841);
    dff g558(.RN(n1), .SN(1'b1), .CK(n0), .D(n1788), .Q(n11[8]));
    buf g559(n12[8], n11[8]);
    or g560(n1864 ,n1034 ,n1582);
    nor g561(n1021 ,n349 ,n66);
    nor g562(n1340 ,n471 ,n54);
    not g563(n582 ,n14[2]);
    dff g564(.RN(n1), .SN(1'b1), .CK(n0), .D(n2003), .Q(n30[19]));
    not g565(n819 ,n69);
    nor g566(n1000 ,n787 ,n69);
    not g567(n2233 ,n24[27]);
    nor g568(n1483 ,n387 ,n44);
    xnor g569(n812 ,n26[10] ,n33[6]);
    xnor g570(n676 ,n181 ,n502);
    or g571(n2134 ,n1452 ,n1653);
    nor g572(n897 ,n794 ,n55);
    not g573(n471 ,n34[24]);
    xnor g574(n2224 ,n23[1] ,n24[1]);
    or g575(n2147 ,n1464 ,n837);
    nor g576(n1619 ,n320 ,n52);
    nor g577(n1140 ,n470 ,n43);
    not g578(n50 ,n52);
    not g579(n199 ,n31[29]);
    nor g580(n1649 ,n327 ,n49);
    not g581(n553 ,n13[26]);
    not g582(n265 ,n4[27]);
    dff g583(.RN(n1), .SN(1'b1), .CK(n0), .D(n2015), .Q(n21[20]));
    nor g584(n976 ,n680 ,n69);
    or g585(n2200 ,n1348 ,n1684);
    nor g586(n1184 ,n127 ,n57);
    not g587(n568 ,n11[21]);
    nor g588(n1060 ,n358 ,n50);
    not g589(n153 ,n24[7]);
    dff g590(.RN(n1), .SN(1'b1), .CK(n0), .D(n2144), .Q(n29[27]));
    or g591(n2219 ,n621 ,n2216);
    nor g592(n861 ,n809 ,n45);
    dff g593(.RN(n1), .SN(1'b1), .CK(n0), .D(n2135), .Q(n24[0]));
    not g594(n244 ,n11[22]);
    nor g595(n1609 ,n345 ,n52);
    nor g596(n1475 ,n557 ,n816);
    or g597(n2320 ,n2317 ,n2318);
    not g598(n516 ,n34[29]);
    not g599(n61 ,n64);
    or g600(n2170 ,n1495 ,n851);
    or g601(n1909 ,n1488 ,n1114);
    dff g602(.RN(n1), .SN(1'b1), .CK(n0), .D(n1896), .Q(n28[8]));
    or g603(n1750 ,n1129 ,n1524);
    or g604(n2321 ,n2319 ,n2316);
    not g605(n301 ,n4[28]);
    not g606(n282 ,n6[1]);
    or g607(n2149 ,n1465 ,n959);
    nor g608(n1372 ,n110 ,n62);
    nor g609(n1394 ,n144 ,n51);
    xnor g610(n757 ,n21[7] ,n24[7]);
    dff g611(.RN(n1), .SN(1'b1), .CK(n0), .D(n1849), .Q(n26[21]));
    not g612(n180 ,n29[24]);
    nor g613(n1124 ,n554 ,n816);
    nor g614(n1316 ,n572 ,n68);
    nor g615(n1627 ,n297 ,n49);
    or g616(n1865 ,n1241 ,n1098);
    not g617(n2235 ,n21[27]);
    dff g618(.RN(n1), .SN(1'b1), .CK(n0), .D(n2158), .Q(n29[24]));
    not g619(n312 ,n5[7]);
    nor g620(n1215 ,n511 ,n61);
    not g621(n99 ,n26[5]);
    not g622(n250 ,n15[1]);
    or g623(n1827 ,n1214 ,n894);
    not g624(n325 ,n5[28]);
    xnor g625(n777 ,n355 ,n141);
    not g626(n525 ,n29[19]);
    not g627(n228 ,n13[31]);
    dff g628(.RN(n1), .SN(1'b1), .CK(n0), .D(n1769), .Q(n11[21]));
    nor g629(n876 ,n737 ,n60);
    not g630(n338 ,n4[18]);
    buf g631(n16[0], n15[8]);
    nor g632(n1006 ,n715 ,n69);
    nor g633(n1646 ,n324 ,n49);
    dff g634(.RN(n1), .SN(1'b1), .CK(n0), .D(n1919), .Q(n35[21]));
    not g635(n114 ,n32[28]);
    or g636(n2040 ,n1276 ,n1569);
    not g637(n185 ,n29[9]);
    or g638(n1954 ,n1334 ,n1669);
    nor g639(n1739 ,n393 ,n66);
    xnor g640(n36[0] ,n2322 ,n25[28]);
    not g641(n363 ,n21[10]);
    xnor g642(n740 ,n21[25] ,n24[25]);
    not g643(n577 ,n13[7]);
    dff g644(.RN(n1), .SN(1'b1), .CK(n0), .D(n1945), .Q(n35[5]));
    or g645(n1791 ,n1171 ,n1549);
    or g646(n1840 ,n1226 ,n901);
    nor g647(n907 ,n759 ,n60);
    dff g648(.RN(n1), .SN(1'b1), .CK(n0), .D(n2149), .Q(n29[26]));
    buf g649(n14[15], n11[15]);
    or g650(n2117 ,n1359 ,n955);
    xnor g651(n632 ,n474 ,n439);
    dff g652(.RN(n1), .SN(1'b1), .CK(n0), .D(n1900), .Q(n31[15]));
    not g653(n304 ,n5[29]);
    dff g654(.RN(n1), .SN(1'b1), .CK(n0), .D(n2014), .Q(n33[31]));
    nor g655(n1334 ,n183 ,n54);
    not g656(n132 ,n32[20]);
    not g657(n548 ,n29[20]);
    dff g658(.RN(n1), .SN(1'b1), .CK(n0), .D(n1966), .Q(n26[8]));
    or g659(n2016 ,n1209 ,n1558);
    nor g660(n1499 ,n609 ,n43);
    dff g661(.RN(n1), .SN(1'b1), .CK(n0), .D(n2169), .Q(n13[16]));
    or g662(n1813 ,n1197 ,n881);
    nor g663(n2209 ,n59 ,n1975);
    not g664(n372 ,n21[12]);
    or g665(n1794 ,n1174 ,n1552);
    nor g666(n1258 ,n435 ,n67);
    nor g667(n1690 ,n152 ,n55);
    or g668(n2198 ,n1295 ,n1685);
    or g669(n2176 ,n1500 ,n854);
    nor g670(n1029 ,n351 ,n66);
    nor g671(n962 ,n712 ,n64);
    or g672(n2291 ,n2237 ,n24[8]);
    buf g673(n14[9], n11[9]);
    dff g674(.RN(n1), .SN(1'b1), .CK(n0), .D(n1955), .Q(n21[31]));
    or g675(n1751 ,n1132 ,n1525);
    buf g676(n14[16], n11[16]);
    nor g677(n1434 ,n428 ,n818);
    xnor g678(n36[1] ,n2322 ,n25[29]);
    not g679(n215 ,n35[22]);
    xnor g680(n752 ,n21[14] ,n24[14]);
    not g681(n2241 ,n21[25]);
    or g682(n1935 ,n1315 ,n938);
    dff g683(.RN(n1), .SN(1'b1), .CK(n0), .D(n1799), .Q(n26[29]));
    dff g684(.RN(n1), .SN(1'b1), .CK(n0), .D(n2130), .Q(n24[3]));
    dff g685(.RN(n1), .SN(1'b1), .CK(n0), .D(n2151), .Q(n13[27]));
    nor g686(n1641 ,n288 ,n52);
    xnor g687(n693 ,n26[23] ,n33[19]);
    not g688(n77 ,n23[3]);
    nor g689(n1114 ,n366 ,n60);
    not g690(n169 ,n29[3]);
    or g691(n1826 ,n1212 ,n892);
    dff g692(.RN(n1), .SN(1'b1), .CK(n0), .D(n1904), .Q(n26[13]));
    nor g693(n1549 ,n440 ,n47);
    dff g694(.RN(n1), .SN(1'b1), .CK(n0), .D(n2189), .Q(n13[6]));
    or g695(n1008 ,n7[3] ,n821);
    not g696(n477 ,n34[21]);
    or g697(n1904 ,n1283 ,n1731);
    not g698(n2234 ,n21[23]);
    nor g699(n1531 ,n123 ,n45);
    dff g700(.RN(n1), .SN(1'b1), .CK(n0), .D(n2055), .Q(n33[8]));
    dff g701(.RN(n1), .SN(1'b1), .CK(n0), .D(n2032), .Q(n30[11]));
    nor g702(n859 ,n812 ,n45);
    dff g703(.RN(n1), .SN(1'b1), .CK(n0), .D(n1834), .Q(n28[30]));
    nor g704(n1321 ,n612 ,n68);
    or g705(n1984 ,n1354 ,n1691);
    xnor g706(n683 ,n207 ,n498);
    dff g707(.RN(n1), .SN(1'b1), .CK(n0), .D(n2175), .Q(n13[13]));
    dff g708(.RN(n1), .SN(1'b1), .CK(n0), .D(n1996), .Q(n34[7]));
    not g709(n603 ,n35[27]);
    or g710(n2272 ,n2243 ,n24[6]);
    nor g711(n1720 ,n397 ,n66);
    or g712(n1762 ,n1136 ,n1019);
    dff g713(.RN(n1), .SN(1'b1), .CK(n0), .D(n1899), .Q(n28[7]));
    not g714(n174 ,n31[20]);
    or g715(n2136 ,n1039 ,n1655);
    or g716(n2123 ,n1442 ,n1643);
    nor g717(n1684 ,n148 ,n56);
    or g718(n1805 ,n1189 ,n875);
    or g719(n2167 ,n1491 ,n826);
    or g720(n1906 ,n1289 ,n979);
    dff g721(.RN(n1), .SN(1'b1), .CK(n0), .D(n1954), .Q(n34[31]));
    dff g722(.RN(n1), .SN(1'b1), .CK(n0), .D(n1880), .Q(n31[25]));
    nor g723(n1272 ,n542 ,n57);
    not g724(n379 ,n30[3]);
    not g725(n437 ,n24[17]);
    or g726(n1030 ,n347 ,n821);
    nor g727(n1144 ,n157 ,n61);
    xnor g728(n785 ,n350 ,n488);
    not g729(n358 ,n21[25]);
    nor g730(n1234 ,n162 ,n57);
    buf g731(n16[13], 1'b0);
    not g732(n206 ,n35[6]);
    not g733(n141 ,n24[0]);
    nor g734(n927 ,n658 ,n56);
    dff g735(.RN(n1), .SN(1'b1), .CK(n0), .D(n2192), .Q(n13[4]));
    dff g736(.RN(n1), .SN(1'b1), .CK(n0), .D(n1995), .Q(n30[21]));
    not g737(n564 ,n11[24]);
    not g738(n76 ,n23[0]);
    not g739(n2244 ,n24[22]);
    or g740(n2306 ,n2290 ,n2289);
    dff g741(.RN(n1), .SN(1'b1), .CK(n0), .D(n2056), .Q(n21[13]));
    or g742(n1806 ,n1190 ,n876);
    or g743(n2035 ,n1385 ,n1710);
    nor g744(n1602 ,n273 ,n49);
    or g745(n2112 ,n1434 ,n1635);
    nor g746(n1191 ,n422 ,n58);
    or g747(n2110 ,n1365 ,n1633);
    or g748(n1939 ,n1320 ,n991);
    not g749(n580 ,n25[31]);
    or g750(n2051 ,n1395 ,n1573);
    xnor g751(n633 ,n549 ,n413);
    nor g752(n969 ,n810 ,n55);
    dff g753(.RN(n1), .SN(1'b1), .CK(n0), .D(n2012), .Q(n21[21]));
    dff g754(.RN(n1), .SN(1'b1), .CK(n0), .D(n1846), .Q(n32[6]));
    nor g755(n885 ,n743 ,n63);
    not g756(n193 ,n28[28]);
    nor g757(n820 ,n626 ,n624);
    dff g758(.RN(n1), .SN(1'b1), .CK(n0), .D(n1988), .Q(n34[25]));
    or g759(n2292 ,n2291 ,n2265);
    dff g760(.RN(n1), .SN(1'b1), .CK(n0), .D(n1865), .Q(n28[20]));
    not g761(n112 ,n32[29]);
    dff g762(.RN(n1), .SN(1'b1), .CK(n0), .D(n2071), .Q(n33[1]));
    or g763(n1776 ,n1155 ,n1538);
    not g764(n411 ,n33[18]);
    nor g765(n1665 ,n114 ,n64);
    nor g766(n1672 ,n127 ,n63);
    dff g767(.RN(n1), .SN(1'b1), .CK(n0), .D(n1776), .Q(n11[17]));
    or g768(n1787 ,n1167 ,n1546);
    dff g769(.RN(n1), .SN(1'b1), .CK(n0), .D(n1961), .Q(n30[31]));
    xnor g770(n745 ,n21[20] ,n24[20]);
    dff g771(.RN(n1), .SN(1'b1), .CK(n0), .D(n2100), .Q(n22[3]));
    nor g772(n1536 ,n563 ,n45);
    nor g773(n1470 ,n571 ,n816);
    nor g774(n940 ,n763 ,n56);
    or g775(n2294 ,n2285 ,n2263);
    or g776(n2160 ,n1479 ,n845);
    or g777(n1862 ,n1240 ,n1725);
    nor g778(n1376 ,n179 ,n53);
    dff g779(.RN(n1), .SN(1'b1), .CK(n0), .D(n2029), .Q(n30[12]));
    nor g780(n1256 ,n168 ,n53);
    xnor g781(n767 ,n21[8] ,n24[8]);
    or g782(n1884 ,n1262 ,n1105);
    xnor g783(n670 ,n543 ,n500);
    or g784(n1801 ,n1184 ,n869);
    nor g785(n1607 ,n323 ,n49);
    dff g786(.RN(n1), .SN(1'b1), .CK(n0), .D(n2017), .Q(n30[15]));
    nor g787(n1207 ,n105 ,n57);
    not g788(n163 ,n29[6]);
    dff g789(.RN(n1), .SN(1'b1), .CK(n0), .D(n2219), .Q(n27[2]));
    or g790(n1994 ,n1358 ,n1663);
    nor g791(n994 ,n689 ,n69);
    dff g792(.RN(n1), .SN(1'b1), .CK(n0), .D(n1840), .Q(n32[9]));
    xnor g793(n723 ,n160 ,n136);
    or g794(n2122 ,n1441 ,n1642);
    not g795(n469 ,n26[13]);
    nor g796(n1738 ,n143 ,n66);
    nor g797(n935 ,n704 ,n63);
    dff g798(.RN(n1), .SN(1'b1), .CK(n0), .D(n1876), .Q(n28[16]));
    nor g799(n1222 ,n423 ,n57);
    dff g800(.RN(n1), .SN(1'b1), .CK(n0), .D(n2164), .Q(n13[19]));
    nor g801(n1432 ,n386 ,n50);
    or g802(n2018 ,n1373 ,n1559);
    nor g803(n947 ,n674 ,n55);
    not g804(n393 ,n33[3]);
    dff g805(.RN(n1), .SN(1'b1), .CK(n0), .D(n1925), .Q(n35[18]));
    or g806(n2118 ,n1439 ,n1640);
    nor g807(n1085 ,n82 ,n48);
    not g808(n166 ,n31[5]);
    or g809(n2052 ,n1396 ,n1574);
    buf g810(n15[15], 1'b0);
    nor g811(n1225 ,n413 ,n57);
    dff g812(.RN(n1), .SN(1'b1), .CK(n0), .D(n1861), .Q(n28[21]));
    dff g813(.RN(n1), .SN(1'b1), .CK(n0), .D(n1905), .Q(n35[30]));
    or g814(n2114 ,n1435 ,n1636);
    nor g815(n1410 ,n588 ,n68);
    dff g816(.RN(n1), .SN(1'b1), .CK(n0), .D(n1820), .Q(n26[26]));
    nor g817(n1175 ,n400 ,n816);
    nor g818(n1055 ,n371 ,n818);
    xnor g819(n665 ,n510 ,n134);
    or g820(n1854 ,n1280 ,n909);
    nor g821(n2212 ,n106 ,n2204);
    or g822(n1759 ,n1131 ,n1018);
    nor g823(n1102 ,n88 ,n59);
    nor g824(n847 ,n714 ,n48);
    dff g825(.RN(n1), .SN(1'b1), .CK(n0), .D(n1928), .Q(n28[2]));
    buf g826(n12[7], n11[7]);
    dff g827(.RN(n1), .SN(1'b1), .CK(n0), .D(n1826), .Q(n32[16]));
    xnor g828(n701 ,n190 ,n512);
    not g829(n395 ,n30[31]);
    xnor g830(n667 ,n508 ,n174);
    dff g831(.RN(n1), .SN(1'b1), .CK(n0), .D(n1783), .Q(n11[12]));
    or g832(n1852 ,n1234 ,n1094);
    nor g833(n1620 ,n344 ,n52);
    nor g834(n1559 ,n567 ,n45);
    nor g835(n854 ,n724 ,n48);
    or g836(n1843 ,n1229 ,n1091);
    or g837(n1842 ,n1228 ,n902);
    nor g838(n2208 ,n27[0] ,n2205);
    nor g839(n623 ,n347 ,n2);
    dff g840(.RN(n1), .SN(1'b1), .CK(n0), .D(n1938), .Q(n26[10]));
    buf g841(n16[2], n15[10]);
    dff g842(.RN(n1), .SN(1'b1), .CK(n0), .D(n1930), .Q(n35[15]));
    dff g843(.RN(n1), .SN(1'b1), .CK(n0), .D(n1878), .Q(n26[15]));
    or g844(n1817 ,n1201 ,n884);
    nor g845(n1724 ,n402 ,n66);
    or g846(n2109 ,n1433 ,n1632);
    or g847(n1928 ,n1427 ,n936);
    or g848(n2003 ,n1364 ,n1700);
    not g849(n490 ,n31[31]);
    dff g850(.RN(n1), .SN(1'b1), .CK(n0), .D(n1870), .Q(n31[29]));
    xnor g851(n811 ,n26[9] ,n33[5]);
    xnor g852(n783 ,n348 ,n537);
    nor g853(n1392 ,n407 ,n816);
    or g854(n1756 ,n1135 ,n1085);
    not g855(n207 ,n34[13]);
    nor g856(n1039 ,n354 ,n50);
    or g857(n1812 ,n1194 ,n1717);
    dff g858(.RN(n1), .SN(1'b1), .CK(n0), .D(n1867), .Q(n31[30]));
    nor g859(n1353 ,n520 ,n54);
    xnor g860(n652 ,n491 ,n457);
    or g861(n814 ,n182 ,n38);
    nor g862(n1041 ,n88 ,n50);
    nor g863(n1197 ,n406 ,n57);
    not g864(n53 ,n56);
    xor g865(n19[6] ,n21[6] ,n22[6]);
    xnor g866(n666 ,n531 ,n521);
    not g867(n332 ,n4[14]);
    nor g868(n960 ,n705 ,n64);
    nor g869(n1014 ,n350 ,n47);
    nor g870(n911 ,n777 ,n60);
    nor g871(n1115 ,n95 ,n66);
    buf g872(n15[14], 1'b0);
    or g873(n823 ,n17[0] ,n820);
    nor g874(n1052 ,n83 ,n57);
    xnor g875(n746 ,n21[19] ,n24[19]);
    buf g876(n12[27], n11[27]);
    nor g877(n1138 ,n507 ,n61);
    xnor g878(n657 ,n509 ,n493);
    or g879(n1872 ,n1250 ,n916);
    nor g880(n891 ,n749 ,n59);
    dff g881(.RN(n1), .SN(1'b1), .CK(n0), .D(n2116), .Q(n24[12]));
    nor g882(n1110 ,n369 ,n60);
    not g883(n201 ,n34[11]);
    xnor g884(n726 ,n193 ,n114);
    dff g885(.RN(n1), .SN(1'b1), .CK(n0), .D(n1813), .Q(n32[24]));
    or g886(n1892 ,n1272 ,n1109);
    nor g887(n1023 ,n75 ,n51);
    buf g888(n14[12], n11[12]);
    nor g889(n890 ,n748 ,n60);
    not g890(n600 ,n14[3]);
    or g891(n2268 ,n2253 ,n24[15]);
    nor g892(n1603 ,n275 ,n817);
    xnor g893(n729 ,n26[4] ,n33[0]);
    nor g894(n922 ,n651 ,n55);
    not g895(n63 ,n62);
    or g896(n2084 ,n1023 ,n1608);
    buf g897(n14[27], n11[27]);
    or g898(n1782 ,n1416 ,n1542);
    nor g899(n837 ,n770 ,n48);
    nor g900(n1146 ,n250 ,n65);
    nor g901(n1585 ,n264 ,n52);
    or g902(n2036 ,n1386 ,n1567);
    nor g903(n996 ,n684 ,n69);
    not g904(n566 ,n11[15]);
    nor g905(n1193 ,n534 ,n61);
    nor g906(n1572 ,n248 ,n47);
    nor g907(n1454 ,n176 ,n62);
    nor g908(n1579 ,n286 ,n49);
    nor g909(n880 ,n740 ,n60);
    or g910(n1747 ,n1516 ,n1029);
    not g911(n387 ,n33[15]);
    or g912(n2297 ,n2286 ,n2261);
    or g913(n2091 ,n1423 ,n1614);
    not g914(n182 ,n7[0]);
    not g915(n2228 ,n21[22]);
    or g916(n2264 ,n24[31] ,n24[30]);
    not g917(n69 ,n68);
    dff g918(.RN(n1), .SN(1'b1), .CK(n0), .D(n1803), .Q(n32[30]));
    nor g919(n1300 ,n215 ,n68);
    xnor g920(n736 ,n159 ,n374);
    dff g921(.RN(n1), .SN(1'b1), .CK(n0), .D(n1957), .Q(n31[0]));
    not g922(n508 ,n34[20]);
    dff g923(.RN(n1), .SN(1'b1), .CK(n0), .D(n2064), .Q(n33[4]));
    dff g924(.RN(n1), .SN(1'b1), .CK(n0), .D(n2134), .Q(n24[1]));
    xnor g925(n700 ,n187 ,n486);
    nor g926(n1521 ,n598 ,n44);
    not g927(n427 ,n26[4]);
    dff g928(.RN(n1), .SN(1'b1), .CK(n0), .D(n1927), .Q(n31[8]));
    dff g929(.RN(n1), .SN(1'b1), .CK(n0), .D(n1959), .Q(n34[28]));
    nor g930(n1541 ,n442 ,n45);
    not g931(n597 ,n25[28]);
    or g932(n1878 ,n1275 ,n1730);
    or g933(n2096 ,n1387 ,n1619);
    or g934(n1811 ,n1195 ,n880);
    not g935(n273 ,n4[10]);
    buf g936(n16[12], 1'b0);
    nor g937(n862 ,n808 ,n48);
    or g938(n2185 ,n1511 ,n857);
    nor g939(n1077 ,n377 ,n61);
    not g940(n255 ,n11[31]);
    buf g941(n16[3], n15[11]);
    nor g942(n1242 ,n482 ,n54);
    dff g943(.RN(n1), .SN(1'b1), .CK(n0), .D(n1869), .Q(n28[18]));
    not g944(n279 ,n4[20]);
    xnor g945(n630 ,n528 ,n448);
    nor g946(n1255 ,n197 ,n57);
    not g947(n135 ,n30[14]);
    nor g948(n948 ,n797 ,n64);
    not g949(n501 ,n35[7]);
    not g950(n155 ,n24[30]);
    nor g951(n1691 ,n453 ,n55);
    buf g952(n14[5], n11[29]);
    xnor g953(n728 ,n76 ,n355);
    or g954(n1757 ,n1137 ,n1084);
    nor g955(n1311 ,n496 ,n54);
    or g956(n2081 ,n1078 ,n1605);
    xnor g957(n36[3] ,n2322 ,n25[31]);
    or g958(n1823 ,n1207 ,n890);
    not g959(n449 ,n26[9]);
    xnor g960(n786 ,n349 ,n505);
    not g961(n361 ,n21[14]);
    not g962(n125 ,n32[21]);
    not g963(n129 ,n24[6]);
    xnor g964(n780 ,n75 ,n501);
    nor g965(n1425 ,n113 ,n818);
    not g966(n534 ,n29[4]);
    not g967(n610 ,n11[17]);
    or g968(n2172 ,n1497 ,n852);
    nor g969(n910 ,n776 ,n59);
    dff g970(.RN(n1), .SN(1'b1), .CK(n0), .D(n2110), .Q(n24[16]));
    nor g971(n1507 ,n498 ,n53);
    nor g972(n1370 ,n414 ,n62);
    or g973(n2097 ,n1025 ,n1617);
    nor g974(n1548 ,n467 ,n48);
    dff g975(.RN(n1), .SN(1'b1), .CK(n0), .D(n2115), .Q(n24[13]));
    or g976(n1951 ,n1474 ,n977);
    nor g977(n1070 ,n363 ,n818);
    nor g978(n1405 ,n143 ,n44);
    not g979(n60 ,n58);
    nor g980(n1064 ,n382 ,n51);
    dff g981(.RN(n1), .SN(1'b1), .CK(n0), .D(n1887), .Q(n31[21]));
    dff g982(.RN(n1), .SN(1'b1), .CK(n0), .D(n1773), .Q(n11[19]));
    xnor g983(n806 ,n349 ,n83);
    nor g984(n1326 ,n165 ,n68);
    or g985(n1868 ,n1243 ,n1099);
    nor g986(n968 ,n677 ,n63);
    not g987(n2229 ,n21[11]);
    or g988(n2026 ,n1043 ,n1596);
    nor g989(n1365 ,n150 ,n51);
    dff g990(.RN(n1), .SN(1'b1), .CK(n0), .D(n2142), .Q(n14[1]));
    not g991(n563 ,n35[23]);
    or g992(n1847 ,n1230 ,n1092);
    nor g993(n1076 ,n89 ,n816);
    or g994(n1815 ,n1198 ,n882);
    nor g995(n1450 ,n580 ,n50);
    xnor g996(n759 ,n21[4] ,n24[4]);
    or g997(n2067 ,n1071 ,n950);
    not g998(n198 ,n29[14]);
    xnor g999(n782 ,n351 ,n165);
    nor g1000(n936 ,n800 ,n59);
    dff g1001(.RN(n1), .SN(1'b1), .CK(n0), .D(n2198), .Q(n34[17]));
    or g1002(n1871 ,n1245 ,n1726);
    or g1003(n1902 ,n1485 ,n978);
    buf g1004(n12[6], n11[6]);
    or g1005(n2174 ,n1496 ,n1116);
    xnor g1006(n788 ,n27[1] ,n106);
    or g1007(n2000 ,n1362 ,n1662);
    nor g1008(n1355 ,n456 ,n62);
    not g1009(n456 ,n30[23]);
    dff g1010(.RN(n1), .SN(1'b1), .CK(n0), .D(n2118), .Q(n24[11]));
    not g1011(n117 ,n30[25]);
    nor g1012(n1443 ,n194 ,n62);
    nor g1013(n1717 ,n400 ,n66);
    dff g1014(.RN(n1), .SN(1'b1), .CK(n0), .D(n1893), .Q(n31[18]));
    nor g1015(n1501 ,n525 ,n61);
    not g1016(n133 ,n24[4]);
    not g1017(n443 ,n33[30]);
    nor g1018(n1710 ,n413 ,n64);
    nor g1019(n1533 ,n138 ,n45);
    not g1020(n289 ,n4[16]);
    not g1021(n331 ,n5[17]);
    buf g1022(n12[25], n11[25]);
    not g1023(n440 ,n26[6]);
    nor g1024(n1447 ,n133 ,n50);
    not g1025(n446 ,n26[10]);
    xnor g1026(n702 ,n156 ,n112);
    or g1027(n2175 ,n1499 ,n853);
    nor g1028(n1056 ,n87 ,n818);
    not g1029(n579 ,n13[2]);
    nor g1030(n964 ,n717 ,n63);
    dff g1031(.RN(n1), .SN(1'b1), .CK(n0), .D(n2049), .Q(n33[12]));
    not g1032(n2248 ,n21[13]);
    or g1033(n2180 ,n1505 ,n825);
    xnor g1034(n779 ,n74 ,n206);
    xnor g1035(n787 ,n186 ,n533);
    or g1036(n2129 ,n1038 ,n1645);
    or g1037(n1941 ,n1411 ,n939);
    nor g1038(n1594 ,n279 ,n817);
    nor g1039(n913 ,n760 ,n55);
    not g1040(n85 ,n21[19]);
    nor g1041(n920 ,n649 ,n56);
    not g1042(n330 ,n4[24]);
    nor g1043(n849 ,n716 ,n47);
    or g1044(n627 ,n106 ,n7[3]);
    nor g1045(n1011 ,n72 ,n818);
    nor g1046(n1082 ,n366 ,n51);
    or g1047(n1841 ,n1223 ,n1722);
    nor g1048(n1065 ,n93 ,n51);
    not g1049(n397 ,n33[24]);
    or g1050(n1918 ,n1448 ,n958);
    nor g1051(n1482 ,n245 ,n51);
    buf g1052(n14[17], n11[17]);
    nor g1053(n1269 ,n174 ,n53);
    nor g1054(n1238 ,n480 ,n54);
    not g1055(n616 ,n13[5]);
    dff g1056(.RN(n1), .SN(1'b1), .CK(n0), .D(n1921), .Q(n35[20]));
    nor g1057(n1111 ,n381 ,n59);
    nor g1058(n912 ,n668 ,n56);
    nor g1059(n887 ,n745 ,n60);
    nor g1060(n1534 ,n404 ,n48);
    xnor g1061(n673 ,n203 ,n536);
    xnor g1062(n772 ,n21[22] ,n24[22]);
    not g1063(n261 ,n11[2]);
    xnor g1064(n797 ,n351 ,n374);
    nor g1065(n1442 ,n434 ,n51);
    dff g1066(.RN(n1), .SN(1'b1), .CK(n0), .D(n1999), .Q(n34[5]));
    nor g1067(n941 ,n702 ,n63);
    dff g1068(.RN(n1), .SN(1'b1), .CK(n0), .D(n1822), .Q(n32[19]));
    nor g1069(n1347 ,n467 ,n67);
    dff g1070(.RN(n1), .SN(1'b1), .CK(n0), .D(n2178), .Q(n13[11]));
    nor g1071(n1498 ,n548 ,n62);
    not g1072(n241 ,n11[8]);
    not g1073(n221 ,n11[10]);
    nor g1074(n1245 ,n137 ,n65);
    nor g1075(n1379 ,n453 ,n62);
    or g1076(n2045 ,n1388 ,n1739);
    dff g1077(.RN(n1), .SN(1'b1), .CK(n0), .D(n1784), .Q(n29[9]));
    nor g1078(n1330 ,n188 ,n54);
    not g1079(n414 ,n30[16]);
    dff g1080(.RN(n1), .SN(1'b1), .CK(n0), .D(n2171), .Q(n15[11]));
    nor g1081(n1469 ,n607 ,n819);
    nor g1082(n1692 ,n392 ,n56);
    dff g1083(.RN(n1), .SN(1'b1), .CK(n0), .D(n1890), .Q(n28[10]));
    dff g1084(.RN(n1), .SN(1'b1), .CK(n0), .D(n1767), .Q(n29[12]));
    not g1085(n360 ,n21[9]);
    nor g1086(n840 ,n653 ,n47);
    not g1087(n98 ,n36[1]);
    nor g1088(n942 ,n630 ,n64);
    nor g1089(n68 ,n40 ,n42);
    nor g1090(n622 ,n346 ,n2);
    nor g1091(n1466 ,n518 ,n53);
    nor g1092(n1382 ,n154 ,n46);
    dff g1093(.RN(n1), .SN(1'b1), .CK(n0), .D(n1833), .Q(n32[12]));
    nor g1094(n1089 ,n365 ,n60);
    or g1095(n1930 ,n1420 ,n987);
    not g1096(n816 ,n45);
    not g1097(n266 ,n5[8]);
    dff g1098(.RN(n1), .SN(1'b1), .CK(n0), .D(n1974), .Q(n34[20]));
    nor g1099(n1514 ,n224 ,n816);
    not g1100(n345 ,n5[30]);
    not g1101(n285 ,n4[1]);
    nor g1102(n972 ,n661 ,n64);
    or g1103(n1844 ,n1045 ,n904);
    nor g1104(n952 ,n803 ,n63);
    not g1105(n195 ,n28[30]);
    xnor g1106(n747 ,n200 ,n370);
    or g1107(n1950 ,n1329 ,n976);
    nor g1108(n1403 ,n425 ,n44);
    or g1109(n1789 ,n1170 ,n1548);
    or g1110(n1899 ,n1279 ,n1111);
    dff g1111(.RN(n1), .SN(1'b1), .CK(n0), .D(n2185), .Q(n13[8]));
    not g1112(n2251 ,n21[12]);
    not g1113(n234 ,n15[10]);
    dff g1114(.RN(n1), .SN(1'b1), .CK(n0), .D(n2048), .Q(n30[7]));
    dff g1115(.RN(n1), .SN(1'b1), .CK(n0), .D(n1920), .Q(n26[12]));
    nor g1116(n1066 ,n361 ,n50);
    not g1117(n461 ,n30[22]);
    nor g1118(n981 ,n641 ,n69);
    not g1119(n520 ,n34[14]);
    nor g1120(n1458 ,n578 ,n50);
    not g1121(n120 ,n24[11]);
    or g1122(n1979 ,n1286 ,n1664);
    dff g1123(.RN(n1), .SN(1'b1), .CK(n0), .D(n2054), .Q(n30[6]));
    or g1124(n624 ,n347 ,n70);
    or g1125(n1956 ,n1311 ,n1670);
    dff g1126(.RN(n1), .SN(1'b1), .CK(n0), .D(n1872), .Q(n31[28]));
    or g1127(n2032 ,n1383 ,n1708);
    nor g1128(n1131 ,n217 ,n65);
    or g1129(n2022 ,n1173 ,n1706);
    nor g1130(n1173 ,n135 ,n61);
    not g1131(n56 ,n54);
    not g1132(n378 ,n21[11]);
    or g1133(n1927 ,n1307 ,n954);
    dff g1134(.RN(n1), .SN(1'b1), .CK(n0), .D(n2044), .Q(n21[15]));
    dff g1135(.RN(n1), .SN(1'b1), .CK(n0), .D(n2091), .Q(n24[27]));
    nor g1136(n959 ,n662 ,n64);
    or g1137(n2275 ,n21[31] ,n21[30]);
    nor g1138(n1503 ,n254 ,n46);
    or g1139(n2192 ,n1519 ,n861);
    nor g1140(n858 ,n687 ,n47);
    or g1141(n2313 ,n2306 ,n2304);
    nor g1142(n919 ,n648 ,n55);
    nor g1143(n1120 ,n82 ,n69);
    xnor g1144(n660 ,n210 ,n110);
    nor g1145(n1596 ,n338 ,n52);
    not g1146(n406 ,n32[24]);
    not g1147(n2230 ,n21[21]);
    or g1148(n1911 ,n1297 ,n1006);
    nor g1149(n1003 ,n667 ,n69);
    not g1150(n444 ,n30[24]);
    dff g1151(.RN(n1), .SN(1'b1), .CK(n0), .D(n1770), .Q(n15[1]));
    nor g1152(n868 ,n696 ,n64);
    or g1153(n2020 ,n1044 ,n1595);
    nor g1154(n1445 ,n129 ,n50);
    nor g1155(n1439 ,n120 ,n818);
    or g1156(n2307 ,n2278 ,n2277);
    not g1157(n173 ,n7[2]);
    not g1158(n451 ,n33[26]);
    nor g1159(n1730 ,n387 ,n66);
    xnor g1160(n713 ,n26[26] ,n33[22]);
    nor g1161(n1496 ,n234 ,n67);
    nor g1162(n828 ,n785 ,n48);
    nor g1163(n993 ,n676 ,n69);
    dff g1164(.RN(n1), .SN(1'b1), .CK(n0), .D(n2007), .Q(n30[18]));
    xnor g1165(n628 ,n191 ,n140);
    not g1166(n2238 ,n20[2]);
    not g1167(n542 ,n28[9]);
    buf g1168(n14[20], n11[20]);
    nor g1169(n1554 ,n238 ,n47);
    or g1170(n1942 ,n1381 ,n992);
    dff g1171(.RN(n1), .SN(1'b1), .CK(n0), .D(n2009), .Q(n34[1]));
    or g1172(n2179 ,n1501 ,n967);
    not g1173(n105 ,n32[18]);
    nor g1174(n1404 ,n446 ,n65);
    nor g1175(n1537 ,n137 ,n45);
    nor g1176(n1271 ,n512 ,n53);
    not g1177(n352 ,n23[1]);
    nor g1178(n1048 ,n376 ,n57);
    or g1179(n1009 ,n17[2] ,n820);
    not g1180(n546 ,n28[23]);
    nor g1181(n1339 ,n532 ,n61);
    nor g1182(n1277 ,n486 ,n53);
    nor g1183(n1524 ,n410 ,n45);
    not g1184(n602 ,n10[2]);
    dff g1185(.RN(n1), .SN(1'b1), .CK(n0), .D(n2051), .Q(n33[11]));
    not g1186(n152 ,n30[13]);
    nor g1187(n999 ,n670 ,n69);
    dff g1188(.RN(n1), .SN(1'b1), .CK(n0), .D(n2090), .Q(n30[1]));
    or g1189(n1824 ,n1208 ,n889);
    or g1190(n1894 ,n1258 ,n1728);
    nor g1191(n1068 ,n372 ,n818);
    nor g1192(n1264 ,n442 ,n67);
    nor g1193(n1280 ,n368 ,n57);
    xnor g1194(n744 ,n21[21] ,n24[21]);
    not g1195(n100 ,n33[29]);
    not g1196(n88 ,n21[16]);
    or g1197(n2298 ,n2269 ,n2275);
    dff g1198(.RN(n1), .SN(1'b1), .CK(n0), .D(n1824), .Q(n29[1]));
    or g1199(n2262 ,n19[1] ,n19[0]);
    nor g1200(n1569 ,n604 ,n47);
    buf g1201(n12[22], n11[22]);
    dff g1202(.RN(n1), .SN(1'b1), .CK(n0), .D(n1823), .Q(n32[18]));
    xnor g1203(n715 ,n503 ,n168);
    nor g1204(n1094 ,n380 ,n59);
    nor g1205(n1119 ,n95 ,n69);
    nor g1206(n916 ,n644 ,n56);
    nor g1207(n1468 ,n605 ,n816);
    xnor g1208(n642 ,n194 ,n432);
    or g1209(n2281 ,n2241 ,n21[24]);
    nor g1210(n1315 ,n502 ,n53);
    nor g1211(n1642 ,n334 ,n817);
    nor g1212(n1268 ,n479 ,n53);
    dff g1213(.RN(n1), .SN(1'b1), .CK(n0), .D(n1936), .Q(n35[11]));
    nor g1214(n1199 ,n445 ,n57);
    not g1215(n510 ,n29[10]);
    nor g1216(n1013 ,n349 ,n818);
    buf g1217(n14[8], n11[8]);
    xnor g1218(n2227 ,n23[0] ,n24[0]);
    nor g1219(n1383 ,n392 ,n61);
    not g1220(n426 ,n24[26]);
    nor g1221(n1007 ,n807 ,n69);
    not g1222(n111 ,n26[8]);
    not g1223(n593 ,n15[7]);
    or g1224(n2002 ,n1367 ,n1738);
    or g1225(n1925 ,n1306 ,n986);
    or g1226(n1910 ,n1294 ,n980);
    dff g1227(.RN(n1), .SN(1'b1), .CK(n0), .D(n1998), .Q(n34[6]));
    or g1228(n1748 ,n1127 ,n824);
    or g1229(n1786 ,n1166 ,n1545);
    or g1230(n2028 ,n1380 ,n1536);
    not g1231(n44 ,n45);
    dff g1232(.RN(n1), .SN(1'b1), .CK(n0), .D(n2172), .Q(n13[14]));
    or g1233(n1822 ,n1206 ,n888);
    dff g1234(.RN(n1), .SN(1'b1), .CK(n0), .D(n1863), .Q(n23[1]));
    nor g1235(n1625 ,n314 ,n49);
    nor g1236(n1700 ,n136 ,n64);
    nor g1237(n1072 ,n96 ,n43);
    or g1238(n1779 ,n1157 ,n867);
    nor g1239(n1575 ,n257 ,n47);
    or g1240(n2125 ,n1443 ,n943);
    nor g1241(n1631 ,n326 ,n817);
    nor g1242(n1489 ,n235 ,n44);
    or g1243(n2266 ,n19[3] ,n19[2]);
    nor g1244(n1477 ,n229 ,n816);
    nor g1245(n1051 ,n370 ,n58);
    not g1246(n122 ,n33[12]);
    nor g1247(n1230 ,n535 ,n57);
    dff g1248(.RN(n1), .SN(1'b1), .CK(n0), .D(n1911), .Q(n35[26]));
    not g1249(n420 ,n32[8]);
    or g1250(n2050 ,n1066 ,n1600);
    dff g1251(.RN(n1), .SN(1'b1), .CK(n0), .D(n2020), .Q(n21[19]));
    dff g1252(.RN(n1), .SN(1'b1), .CK(n0), .D(n1946), .Q(n35[4]));
    not g1253(n405 ,n26[17]);
    or g1254(n1784 ,n1164 ,n868);
    not g1255(n232 ,n13[20]);
    or g1256(n2273 ,n2246 ,n24[17]);
    not g1257(n2255 ,n19[5]);
    not g1258(n341 ,n5[20]);
    nor g1259(n1415 ,n439 ,n57);
    nor g1260(n1530 ,n130 ,n48);
    xnor g1261(n795 ,n75 ,n384);
    or g1262(n2315 ,n2307 ,n2300);
    not g1263(n2254 ,n21[15]);
    nor g1264(n1444 ,n153 ,n50);
    xnor g1265(n709 ,n26[27] ,n33[23]);
    not g1266(n321 ,n5[2]);
    or g1267(n1973 ,n1345 ,n1665);
    or g1268(n2289 ,n2230 ,n2236);
    not g1269(n52 ,n51);
    or g1270(n2148 ,n1467 ,n838);
    or g1271(n2060 ,n1068 ,n1659);
    nor g1272(n1522 ,n579 ,n46);
    xnor g1273(n731 ,n513 ,n384);
    nor g1274(n1706 ,n140 ,n64);
    not g1275(n220 ,n11[23]);
    dff g1276(.RN(n1), .SN(1'b1), .CK(n0), .D(n2037), .Q(n33[18]));
    dff g1277(.RN(n1), .SN(1'b1), .CK(n0), .D(n2001), .Q(n34[4]));
    dff g1278(.RN(n1), .SN(1'b1), .CK(n0), .D(n2156), .Q(n13[25]));
    dff g1279(.RN(n1), .SN(1'b1), .CK(n0), .D(n1923), .Q(n35[19]));
    not g1280(n227 ,n15[0]);
    dff g1281(.RN(n1), .SN(1'b1), .CK(n0), .D(n2069), .Q(n33[2]));
    not g1282(n570 ,n10[1]);
    or g1283(n2284 ,n2244 ,n24[23]);
    nor g1284(n1416 ,n237 ,n46);
    not g1285(n601 ,n11[18]);
    xnor g1286(n815 ,n26[12] ,n33[8]);
    not g1287(n584 ,n13[19]);
    xnor g1288(n732 ,n492 ,n362);
    nor g1289(n1047 ,n374 ,n58);
    nor g1290(n1356 ,n201 ,n53);
    nor g1291(n1053 ,n375 ,n51);
    or g1292(n1993 ,n1351 ,n1737);
    xor g1293(n19[7] ,n21[7] ,n22[7]);
    nor g1294(n836 ,n779 ,n45);
    or g1295(n1856 ,n1051 ,n910);
    buf g1296(n16[1], n15[9]);
    or g1297(n1885 ,n1265 ,n922);
    not g1298(n179 ,n31[3]);
    xnor g1299(n721 ,n487 ,n517);
    nor g1300(n2221 ,n2208 ,n2218);
    nor g1301(n1343 ,n205 ,n53);
    nor g1302(n1423 ,n115 ,n51);
    or g1303(n1946 ,n1327 ,n998);
    nor g1304(n1651 ,n321 ,n52);
    dff g1305(.RN(n1), .SN(1'b1), .CK(n0), .D(n2150), .Q(n13[28]));
    or g1306(n1953 ,n1333 ,n997);
    nor g1307(n1624 ,n339 ,n49);
    nor g1308(n923 ,n652 ,n56);
    dff g1309(.RN(n1), .SN(1'b1), .CK(n0), .D(n2043), .Q(n33[15]));
    not g1310(n412 ,n26[11]);
    or g1311(n2182 ,n1508 ,n856);
    or g1312(n1982 ,n1313 ,n1690);
    dff g1313(.RN(n1), .SN(1'b1), .CK(n0), .D(n2157), .Q(n13[24]));
    nor g1314(n1673 ,n452 ,n56);
    or g1315(n2133 ,n1450 ,n1646);
    nor g1316(n1346 ,n508 ,n53);
    not g1317(n74 ,n22[6]);
    not g1318(n290 ,n3[29]);
    dff g1319(.RN(n1), .SN(1'b1), .CK(n0), .D(n1871), .Q(n26[18]));
    or g1320(n2047 ,n1392 ,n1572);
    nor g1321(n1275 ,n462 ,n67);
    dff g1322(.RN(n1), .SN(1'b1), .CK(n0), .D(n1908), .Q(n28[5]));
    dff g1323(.RN(n1), .SN(1'b1), .CK(n0), .D(n1862), .Q(n26[19]));
    or g1324(n2099 ,n1428 ,n1623);
    or g1325(n2008 ,n1177 ,n1740);
    not g1326(n93 ,n21[15]);
    xnor g1327(n674 ,n524 ,n389);
    nor g1328(n1393 ,n431 ,n61);
    nor g1329(n1279 ,n513 ,n57);
    nor g1330(n1176 ,n592 ,n43);
    not g1331(n613 ,n35[30]);
    nor g1332(n1449 ,n421 ,n50);
    dff g1333(.RN(n1), .SN(1'b1), .CK(n0), .D(n2126), .Q(n24[6]));
    nor g1334(n1237 ,n167 ,n58);
    nor g1335(n1674 ,n429 ,n56);
    not g1336(n552 ,n11[26]);
    dff g1337(.RN(n1), .SN(1'b1), .CK(n0), .D(n2202), .Q(n26[1]));
    nor g1338(n903 ,n791 ,n55);
    nor g1339(n1568 ,n561 ,n48);
    or g1340(n2006 ,n1221 ,n897);
    not g1341(n555 ,n11[25]);
    nor g1342(n1002 ,n700 ,n69);
    nor g1343(n1332 ,n111 ,n67);
    or g1344(n2187 ,n1515 ,n970);
    or g1345(n1917 ,n1300 ,n983);
    or g1346(n2319 ,n2313 ,n2315);
    nor g1347(n1551 ,n603 ,n45);
    nor g1348(n1563 ,n607 ,n45);
    xnor g1349(n724 ,n26[16] ,n33[12]);
    not g1350(n314 ,n5[21]);
    nor g1351(n1656 ,n284 ,n52);
    nor g1352(n1737 ,n425 ,n66);
    nor g1353(n1740 ,n468 ,n66);
    or g1354(n1887 ,n1268 ,n923);
    nor g1355(n1733 ,n409 ,n66);
    nor g1356(n1389 ,n466 ,n44);
    nor g1357(n1492 ,n491 ,n61);
    nor g1358(n2220 ,n2207 ,n2217);
    nor g1359(n1462 ,n597 ,n818);
    not g1360(n246 ,n13[29]);
    dff g1361(.RN(n1), .SN(1'b1), .CK(n0), .D(n2023), .Q(n33[26]));
    nor g1362(n1390 ,n398 ,n62);
    or g1363(n2137 ,n1040 ,n1656);
    not g1364(n572 ,n35[12]);
    xnor g1365(n719 ,n26[19] ,n33[15]);
    dff g1366(.RN(n1), .SN(1'b1), .CK(n0), .D(n1944), .Q(n31[3]));
    dff g1367(.RN(n1), .SN(1'b1), .CK(n0), .D(n2057), .Q(n33[7]));
    nor g1368(n1042 ,n94 ,n50);
    not g1369(n407 ,n33[13]);
    dff g1370(.RN(n1), .SN(1'b1), .CK(n0), .D(n2077), .Q(n10[2]));
    dff g1371(.RN(n1), .SN(1'b1), .CK(n0), .D(n2222), .Q(n27[1]));
    nor g1372(n967 ,n723 ,n64);
    nor g1373(n1448 ,n533 ,n53);
    nor g1374(n1220 ,n195 ,n58);
    nor g1375(n1438 ,n526 ,n61);
    dff g1376(.RN(n1), .SN(1'b1), .CK(n0), .D(n1962), .Q(n34[26]));
    nor g1377(n1318 ,n200 ,n57);
    dff g1378(.RN(n1), .SN(1'b1), .CK(n0), .D(n2155), .Q(n13[26]));
    dff g1379(.RN(n1), .SN(1'b1), .CK(n0), .D(n1968), .Q(n30[29]));
    nor g1380(n1252 ,n461 ,n61);
    or g1381(n2039 ,n1041 ,n1598);
    nor g1382(n621 ,n71 ,n2);
    or g1383(n2061 ,n1403 ,n836);
    or g1384(n2071 ,n1072 ,n828);
    not g1385(n281 ,n5[6]);
    dff g1386(.RN(n1), .SN(1'b1), .CK(n0), .D(n1818), .Q(n32[21]));
    dff g1387(.RN(n1), .SN(1'b1), .CK(n0), .D(n1972), .Q(n34[21]));
    nor g1388(n844 ,n709 ,n48);
    or g1389(n2186 ,n1513 ,n858);
    or g1390(n1970 ,n1057 ,n1586);
    not g1391(n2252 ,n24[12]);
    dff g1392(.RN(n1), .SN(1'b1), .CK(n0), .D(n1982), .Q(n34[13]));
    not g1393(n575 ,n35[16]);
    nor g1394(n931 ,n663 ,n56);
    nor g1395(n1582 ,n277 ,n52);
    nor g1396(n1251 ,n509 ,n53);
    nor g1397(n1519 ,n219 ,n43);
    not g1398(n346 ,n27[1]);
    not g1399(n617 ,n35[15]);
    nor g1400(n1153 ,n583 ,n44);
    or g1401(n1793 ,n1172 ,n1550);
    dff g1402(.RN(n1), .SN(1'b1), .CK(n0), .D(n1847), .Q(n28[26]));
    or g1403(n1922 ,n1305 ,n956);
    dff g1404(.RN(n1), .SN(1'b1), .CK(n0), .D(n2167), .Q(n13[17]));
    nor g1405(n977 ,n686 ,n69);
    not g1406(n75 ,n22[7]);
    nor g1407(n1584 ,n267 ,n49);
    buf g1408(n12[14], n11[14]);
    xnor g1409(n769 ,n21[16] ,n24[16]);
    nor g1410(n872 ,n732 ,n63);
    not g1411(n131 ,n24[20]);
    not g1412(n2231 ,n21[17]);
    dff g1413(.RN(n1), .SN(1'b1), .CK(n0), .D(n2154), .Q(n25[29]));
    xnor g1414(n645 ,n26[29] ,n33[25]);
    or g1415(n1849 ,n1231 ,n1723);
    nor g1416(n1161 ,n385 ,n67);
    nor g1417(n1360 ,n457 ,n61);
    nor g1418(n1098 ,n382 ,n60);
    nor g1419(n1433 ,n437 ,n818);
    not g1420(n144 ,n24[28]);
    dff g1421(.RN(n1), .SN(1'b1), .CK(n0), .D(n1796), .Q(n11[2]));
    nor g1422(n1322 ,n161 ,n53);
    nor g1423(n963 ,n690 ,n63);
    dff g1424(.RN(n1), .SN(1'b1), .CK(n0), .D(n1841), .Q(n26[22]));
    dff g1425(.RN(n1), .SN(1'b1), .CK(n0), .D(n1953), .Q(n35[0]));
    not g1426(n465 ,n24[24]);
    not g1427(n310 ,n4[17]);
    nor g1428(n1734 ,n417 ,n66);
    dff g1429(.RN(n1), .SN(1'b1), .CK(n0), .D(n1907), .Q(n31[13]));
    not g1430(n260 ,n13[10]);
    nor g1431(n1663 ,n398 ,n56);
    dff g1432(.RN(n1), .SN(1'b1), .CK(n0), .D(n1831), .Q(n32[13]));
    dff g1433(.RN(n1), .SN(1'b1), .CK(n0), .D(n2045), .Q(n26[3]));
    nor g1434(n1267 ,n202 ,n57);
    dff g1435(.RN(n1), .SN(1'b1), .CK(n0), .D(n1976), .Q(n34[16]));
    not g1436(n435 ,n26[16]);
    or g1437(n2282 ,n2235 ,n21[26]);
    nor g1438(n1687 ,n110 ,n56);
    not g1439(n95 ,n36[3]);
    nor g1440(n1080 ,n81 ,n818);
    dff g1441(.RN(n1), .SN(1'b1), .CK(n0), .D(n1971), .Q(n34[22]));
    dff g1442(.RN(n1), .SN(1'b1), .CK(n0), .D(n2076), .Q(n10[3]));
    nor g1443(n946 ,n730 ,n55);
    dff g1444(.RN(n1), .SN(1'b1), .CK(n0), .D(n2078), .Q(n10[1]));
    nor g1445(n1113 ,n91 ,n60);
    dff g1446(.RN(n1), .SN(1'b1), .CK(n0), .D(n1914), .Q(n31[11]));
    or g1447(n2193 ,n1521 ,n862);
    not g1448(n48 ,n46);
    buf g1449(n17[4], 1'b0);
    not g1450(n517 ,n31[27]);
    nor g1451(n1276 ,n447 ,n43);
    nor g1452(n1618 ,n343 ,n49);
    nor g1453(n1576 ,n612 ,n45);
    not g1454(n2257 ,n19[6]);
    nor g1455(n1289 ,n567 ,n819);
    dff g1456(.RN(n1), .SN(1'b1), .CK(n0), .D(n1997), .Q(n21[23]));
    nor g1457(n908 ,n775 ,n60);
    not g1458(n108 ,n26[22]);
    nor g1459(n1301 ,n172 ,n57);
    nor g1460(n1652 ,n318 ,n49);
    buf g1461(n14[30], n12[30]);
    not g1462(n531 ,n34[22]);
    nor g1463(n1045 ,n384 ,n57);
    not g1464(n374 ,n32[5]);
    dff g1465(.RN(n1), .SN(1'b1), .CK(n0), .D(n2101), .Q(n24[21]));
    nor g1466(n1351 ,n440 ,n67);
    dff g1467(.RN(n1), .SN(1'b1), .CK(n0), .D(n2190), .Q(n15[7]));
    or g1468(n1924 ,n1303 ,n1741);
    not g1469(n598 ,n13[3]);
    dff g1470(.RN(n1), .SN(1'b1), .CK(n0), .D(n2131), .Q(n29[29]));
    or g1471(n2087 ,n1024 ,n1610);
    not g1472(n191 ,n28[14]);
    or g1473(n2111 ,n1013 ,n1631);
    nor g1474(n1719 ,n430 ,n66);
    or g1475(n2144 ,n1461 ,n935);
    nor g1476(n924 ,n654 ,n55);
    or g1477(n1769 ,n1151 ,n1533);
    dff g1478(.RN(n1), .SN(1'b1), .CK(n0), .D(n1895), .Q(n31[17]));
    xnor g1479(n821 ,n27[2] ,n173);
    or g1480(n2305 ,n2288 ,n2279);
    not g1481(n134 ,n30[10]);
    or g1482(n1967 ,n1340 ,n1709);
    not g1483(n158 ,n29[31]);
    or g1484(n2019 ,n1182 ,n1560);
    nor g1485(n1270 ,n549 ,n57);
    dff g1486(.RN(n1), .SN(1'b1), .CK(n0), .D(n1828), .Q(n29[0]));
    nor g1487(n1406 ,n116 ,n61);
    xnor g1488(n761 ,n98 ,n100);
    nor g1489(n1399 ,n589 ,n68);
    nor g1490(n1019 ,n348 ,n66);
    not g1491(n436 ,n26[27]);
    not g1492(n313 ,n9[3]);
    nor g1493(n1028 ,n74 ,n66);
    nor g1494(n1099 ,n85 ,n60);
    not g1495(n487 ,n34[27]);
    not g1496(n231 ,n12[29]);
    buf g1497(n12[10], n11[10]);
    dff g1498(.RN(n1), .SN(1'b1), .CK(n0), .D(n1754), .Q(n12[28]));
    or g1499(n2190 ,n1742 ,n1027);
    not g1500(n428 ,n24[15]);
    dff g1501(.RN(n1), .SN(1'b1), .CK(n0), .D(n2033), .Q(n33[21]));
    not g1502(n140 ,n32[14]);
    nor g1503(n954 ,n688 ,n55);
    buf g1504(n16[9], n15[5]);
    nor g1505(n1250 ,n523 ,n53);
    not g1506(n2243 ,n24[7]);
    nor g1507(n1293 ,n543 ,n53);
    nor g1508(n1600 ,n332 ,n49);
    not g1509(n357 ,n32[3]);
    dff g1510(.RN(n1), .SN(1'b1), .CK(n0), .D(n2086), .Q(n21[27]));
    xnor g1511(n763 ,n540 ,n373);
    dff g1512(.RN(n1), .SN(1'b1), .CK(n0), .D(n1800), .Q(n11[0]));
    dff g1513(.RN(n1), .SN(1'b1), .CK(n0), .D(n1794), .Q(n11[4]));
    buf g1514(n12[21], n11[21]);
    nor g1515(n1035 ,n80 ,n51);
    xnor g1516(n662 ,n535 ,n109);
    xnor g1517(n641 ,n205 ,n189);
    or g1518(n1893 ,n1274 ,n926);
    nor g1519(n1670 ,n432 ,n55);
    not g1520(n348 ,n22[2]);
    or g1521(n2128 ,n1447 ,n1649);
    dff g1522(.RN(n1), .SN(1'b1), .CK(n0), .D(n1785), .Q(n11[11]));
    not g1523(n605 ,n13[28]);
    nor g1524(n1061 ,n84 ,n50);
    not g1525(n97 ,n21[28]);
    dff g1526(.RN(n1), .SN(1'b1), .CK(n0), .D(n2095), .Q(n26[0]));
    not g1527(n481 ,n31[18]);
    xnor g1528(n649 ,n180 ,n444);
    not g1529(n170 ,n31[0]);
    dff g1530(.RN(n1), .SN(1'b1), .CK(n0), .D(n1775), .Q(n11[18]));
    xnor g1531(n739 ,n545 ,n376);
    nor g1532(n1408 ,n393 ,n816);
    or g1533(n2265 ,n24[11] ,n24[10]);
    nor g1534(n1168 ,n472 ,n61);
    nor g1535(n1058 ,n365 ,n51);
    nor g1536(n833 ,n784 ,n45);
    not g1537(n238 ,n26[2]);
    nor g1538(n939 ,n634 ,n56);
    nor g1539(n1708 ,n423 ,n63);
    nor g1540(n1517 ,n243 ,n65);
    buf g1541(n16[6], n15[2]);
    nor g1542(n1162 ,n586 ,n44);
    or g1543(n1851 ,n1048 ,n907);
    not g1544(n354 ,n18[1]);
    nor g1545(n1181 ,n455 ,n67);
    dff g1546(.RN(n1), .SN(1'b1), .CK(n0), .D(n1877), .Q(n31[26]));
    dff g1547(.RN(n1), .SN(1'b1), .CK(n0), .D(n1780), .Q(n15[0]));
    nor g1548(n1506 ,n240 ,n65);
    xnor g1549(n714 ,n26[24] ,n33[20]);
    or g1550(n2169 ,n1494 ,n850);
    nor g1551(n1200 ,n107 ,n65);
    nor g1552(n1661 ,n439 ,n64);
    nor g1553(n1348 ,n171 ,n53);
    not g1554(n274 ,n4[22]);
    dff g1555(.RN(n1), .SN(1'b1), .CK(n0), .D(n2133), .Q(n25[31]));
    dff g1556(.RN(n1), .SN(1'b1), .CK(n0), .D(n1933), .Q(n35[13]));
    not g1557(n489 ,n31[24]);
    nor g1558(n1071 ,n379 ,n61);
    xnor g1559(n639 ,n196 ,n504);
    xnor g1560(n682 ,n477 ,n479);
    nor g1561(n966 ,n796 ,n63);
    nor g1562(n1359 ,n158 ,n62);
    not g1563(n161 ,n34[23]);
    dff g1564(.RN(n1), .SN(1'b1), .CK(n0), .D(n2079), .Q(n30[0]));
    or g1565(n1800 ,n1183 ,n1556);
    not g1566(n433 ,n24[31]);
    or g1567(n1848 ,n1047 ,n906);
    or g1568(n2120 ,n1037 ,n1639);
    dff g1569(.RN(n1), .SN(1'b1), .CK(n0), .D(n2050), .Q(n21[14]));
    not g1570(n118 ,n32[16]);
    dff g1571(.RN(n1), .SN(1'b1), .CK(n0), .D(n2153), .Q(n35[24]));
    nor g1572(n1130 ,n198 ,n62);
    nor g1573(n1198 ,n169 ,n61);
    xnor g1574(n19[0] ,n2226 ,n18[0]);
    or g1575(n1879 ,n1255 ,n1103);
    dff g1576(.RN(n1), .SN(1'b1), .CK(n0), .D(n1804), .Q(n32[29]));
    not g1577(n83 ,n32[0]);
    dff g1578(.RN(n1), .SN(1'b1), .CK(n0), .D(n1790), .Q(n29[8]));
    dff g1579(.RN(n1), .SN(1'b1), .CK(n0), .D(n2013), .Q(n30[16]));
    dff g1580(.RN(n1), .SN(1'b1), .CK(n0), .D(n2083), .Q(n24[30]));
    not g1581(n275 ,n4[9]);
    nor g1582(n1281 ,n627 ,n814);
    not g1583(n350 ,n22[1]);
    or g1584(n1948 ,n1328 ,n940);
    nor g1585(n1037 ,n353 ,n818);
    or g1586(n2300 ,n2266 ,n2262);
    nor g1587(n1254 ,n181 ,n53);
    nor g1588(n1639 ,n285 ,n52);
    not g1589(n550 ,n34[3]);
    not g1590(n558 ,n13[9]);
    not g1591(n249 ,n15[2]);
    xnor g1592(n755 ,n21[10] ,n24[10]);
    not g1593(n147 ,n30[20]);
    not g1594(n382 ,n21[20]);
    not g1595(n513 ,n28[7]);
    not g1596(n329 ,n4[21]);
    or g1597(n2116 ,n1368 ,n1638);
    or g1598(n2311 ,n2303 ,n2299);
    dff g1599(.RN(n1), .SN(1'b1), .CK(n0), .D(n2061), .Q(n33[6]));
    or g1600(n1775 ,n1154 ,n1537);
    nor g1601(n1409 ,n464 ,n46);
    nor g1602(n1187 ,n408 ,n57);
    dff g1603(.RN(n1), .SN(1'b1), .CK(n0), .D(n2168), .Q(n29[21]));
    not g1604(n524 ,n29[5]);
    nor g1605(n886 ,n744 ,n59);
    dff g1606(.RN(n1), .SN(1'b1), .CK(n0), .D(n2105), .Q(n21[4]));
    nor g1607(n1097 ,n383 ,n59);
    not g1608(n47 ,n46);
    nor g1609(n1697 ,n431 ,n55);
    not g1610(n502 ,n31[6]);
    or g1611(n1853 ,n1049 ,n908);
    nor g1612(n984 ,n682 ,n69);
    xnor g1613(n672 ,n163 ,n450);
    not g1614(n217 ,n15[3]);
    xor g1615(n1975 ,n727 ,n18[1]);
    or g1616(n1818 ,n1203 ,n886);
    dff g1617(.RN(n1), .SN(1'b1), .CK(n0), .D(n1764), .Q(n11[25]));
    not g1618(n403 ,n30[28]);
    or g1619(n2121 ,n1440 ,n1641);
    not g1620(n519 ,n35[4]);
    xnor g1621(n784 ,n72 ,n211);
    nor g1622(n1135 ,n587 ,n816);
    or g1623(n2086 ,n1056 ,n1587);
    not g1624(n464 ,n33[2]);
    nor g1625(n1118 ,n92 ,n66);
    nor g1626(n1158 ,n566 ,n43);
    buf g1627(n14[31], n12[31]);
    not g1628(n106 ,n7[1]);
    dff g1629(.RN(n1), .SN(1'b1), .CK(n0), .D(n1812), .Q(n26[27]));
    or g1630(n1895 ,n1277 ,n927);
    buf g1631(n12[9], n11[9]);
    or g1632(n1976 ,n1293 ,n1686);
    dff g1633(.RN(n1), .SN(1'b1), .CK(n0), .D(n2139), .Q(n29[28]));
    or g1634(n1820 ,n1200 ,n1718);
    or g1635(n2108 ,n1010 ,n1629);
    dff g1636(.RN(n1), .SN(1'b1), .CK(n0), .D(n2166), .Q(n13[18]));
    dff g1637(.RN(n1), .SN(1'b1), .CK(n0), .D(n1947), .Q(n35[3]));
    not g1638(n385 ,n26[31]);
    buf g1639(n12[23], n11[23]);
    xnor g1640(n638 ,n197 ,n145);
    nor g1641(n1043 ,n90 ,n50);
    or g1642(n2274 ,n2254 ,n21[14]);
    xor g1643(n1744 ,n728 ,n18[0]);
    nor g1644(n1325 ,n206 ,n68);
    nor g1645(n1204 ,n540 ,n61);
    or g1646(n2115 ,n1436 ,n1637);
    not g1647(n121 ,n32[9]);
    nor g1648(n1688 ,n135 ,n56);
    or g1649(n1833 ,n1415 ,n898);
    or g1650(n2296 ,n2268 ,n2267);
    dff g1651(.RN(n1), .SN(1'b1), .CK(n0), .D(n1987), .Q(n21[25]));
    not g1652(n2250 ,n24[25]);
    nor g1653(n1681 ,n422 ,n64);
    dff g1654(.RN(n1), .SN(1'b1), .CK(n0), .D(n2173), .Q(n29[20]));
    or g1655(n2143 ,n1460 ,n1017);
    not g1656(n509 ,n34[9]);
    or g1657(n1797 ,n1178 ,n871);
    or g1658(n2194 ,n1520 ,n972);
    not g1659(n102 ,n33[23]);
    or g1660(n1760 ,n1139 ,n1086);
    not g1661(n110 ,n30[15]);
    not g1662(n328 ,n4[13]);
    nor g1663(n1209 ,n443 ,n43);
    xnor g1664(n681 ,n483 ,n170);
    or g1665(n2158 ,n1476 ,n961);
    dff g1666(.RN(n1), .SN(1'b1), .CK(n0), .D(n2165), .Q(n29[22]));
    not g1667(n200 ,n28[1]);
    nor g1668(n1629 ,n278 ,n49);
    or g1669(n2139 ,n1454 ,n957);
    or g1670(n2001 ,n1363 ,n1701);
    dff g1671(.RN(n1), .SN(1'b1), .CK(n0), .D(n1836), .Q(n28[28]));
    not g1672(n518 ,n31[14]);
    not g1673(n606 ,n11[20]);
    nor g1674(n1384 ,n402 ,n46);
    not g1675(n151 ,n33[19]);
    dff g1676(.RN(n1), .SN(1'b1), .CK(n0), .D(n1909), .Q(n28[4]));
    or g1677(n2011 ,n1371 ,n945);
    not g1678(n554 ,n13[1]);
    or g1679(n2064 ,n1407 ,n832);
    nor g1680(n1202 ,n463 ,n65);
    xnor g1681(n809 ,n26[8] ,n33[4]);
    nor g1682(n938 ,n672 ,n56);
    dff g1683(.RN(n1), .SN(1'b1), .CK(n0), .D(n2005), .Q(n21[22]));
    not g1684(n607 ,n35[24]);
    or g1685(n2057 ,n1401 ,n830);
    nor g1686(n1467 ,n246 ,n44);
    not g1687(n149 ,n24[5]);
    not g1688(n486 ,n31[17]);
    not g1689(n263 ,n13[17]);
    nor g1690(n1157 ,n510 ,n61);
    nor g1691(n1163 ,n620 ,n44);
    dff g1692(.RN(n1), .SN(1'b1), .CK(n0), .D(n2193), .Q(n13[3]));
    nor g1693(n973 ,n638 ,n63);
    dff g1694(.RN(n1), .SN(1'b1), .CK(n0), .D(n2104), .Q(n24[20]));
    or g1695(n1788 ,n1169 ,n1547);
    dff g1696(.RN(n1), .SN(1'b1), .CK(n0), .D(n1913), .Q(n35[25]));
    not g1697(n229 ,n13[24]);
    xnor g1698(n707 ,n162 ,n406);
    nor g1699(n956 ,n629 ,n55);
    or g1700(n1804 ,n1188 ,n874);
    dff g1701(.RN(n1), .SN(1'b1), .CK(n0), .D(n1951), .Q(n35[1]));
    not g1702(n389 ,n30[5]);
    dff g1703(.RN(n1), .SN(1'b1), .CK(n0), .D(n1765), .Q(n11[24]));
    or g1704(n2132 ,n1451 ,n1651);
    nor g1705(n900 ,n755 ,n60);
    nor g1706(n1686 ,n414 ,n55);
    nor g1707(n1570 ,n575 ,n48);
    or g1708(n2070 ,n1504 ,n1512);
    dff g1709(.RN(n1), .SN(1'b1), .CK(n0), .D(n1980), .Q(n34[14]));
    dff g1710(.RN(n1), .SN(1'b1), .CK(n0), .D(n2065), .Q(n21[11]));
    not g1711(n390 ,n33[31]);
    dff g1712(.RN(n1), .SN(1'b1), .CK(n0), .D(n2034), .Q(n33[20]));
    nor g1713(n1179 ,n261 ,n43);
    nor g1714(n1327 ,n519 ,n68);
    xnor g1715(n748 ,n21[18] ,n24[18]);
    not g1716(n308 ,n4[19]);
    nor g1717(n1246 ,n164 ,n53);
    not g1718(n311 ,n4[2]);
    buf g1719(n14[29], n12[29]);
    dff g1720(.RN(n1), .SN(1'b1), .CK(n0), .D(n1894), .Q(n26[16]));
    xnor g1721(n671 ,n520 ,n518);
    nor g1722(n857 ,n815 ,n45);
    buf g1723(n14[11], n11[11]);
    or g1724(n1905 ,n1288 ,n995);
    not g1725(n528 ,n28[13]);
    not g1726(n521 ,n31[22]);
    nor g1727(n1366 ,n148 ,n61);
    nor g1728(n1224 ,n156 ,n57);
    or g1729(n1990 ,n1054 ,n1590);
    or g1730(n1754 ,n1133 ,n1526);
    nor g1731(n1079 ,n86 ,n61);
    nor g1732(n1350 ,n429 ,n61);
    nor g1733(n1511 ,n253 ,n43);
    not g1734(n543 ,n34[16]);
    or g1735(n2277 ,n2231 ,n21[16]);
    nor g1736(n1229 ,n538 ,n57);
    or g1737(n1998 ,n1254 ,n1698);
    not g1738(n404 ,n26[20]);
    or g1739(n2261 ,n20[1] ,n20[0]);
    buf g1740(n12[18], n11[18]);
    dff g1741(.RN(n1), .SN(1'b1), .CK(n0), .D(n1917), .Q(n35[22]));
    nor g1742(n1455 ,n600 ,n816);
    or g1743(n2126 ,n1445 ,n1647);
    not g1744(n470 ,n33[21]);
    nor g1745(n1660 ,n328 ,n49);
    nor g1746(n1595 ,n308 ,n49);
    not g1747(n475 ,n28[20]);
    xnor g1748(n775 ,n80 ,n421);
    nor g1749(n1701 ,n116 ,n55);
    nor g1750(n1117 ,n98 ,n66);
    nor g1751(n1702 ,n105 ,n63);
    nor g1752(n1169 ,n241 ,n46);
    xnor g1753(n20[1] ,n2224 ,n18[1]);
    xnor g1754(n718 ,n26[20] ,n33[16]);
    or g1755(n1765 ,n1145 ,n1530);
    nor g1756(n1722 ,n154 ,n66);
    or g1757(n1981 ,n1347 ,n1736);
    not g1758(n398 ,n30[8]);
    dff g1759(.RN(n1), .SN(1'b1), .CK(n0), .D(n2188), .Q(n15[8]));
    not g1760(n594 ,n11[27]);
    buf g1761(n14[23], n11[23]);
    nor g1762(n930 ,n703 ,n56);
    or g1763(n2073 ,n1076 ,n834);
    nor g1764(n1398 ,n608 ,n68);
    nor g1765(n1664 ,n415 ,n64);
    not g1766(n309 ,n5[11]);
    nor g1767(n841 ,n706 ,n47);
    nor g1768(n1693 ,n134 ,n55);
    dff g1769(.RN(n1), .SN(1'b1), .CK(n0), .D(n1755), .Q(n11[31]));
    or g1770(n2285 ,n2229 ,n2259);
    or g1771(n1923 ,n1437 ,n985);
    nor g1772(n878 ,n739 ,n63);
    xnor g1773(n636 ,n484 ,n420);
    or g1774(n2103 ,n1012 ,n1624);
    not g1775(n578 ,n25[30]);
    xnor g1776(n705 ,n204 ,n415);
    or g1777(n2287 ,n2249 ,n2257);
    not g1778(n514 ,n31[15]);
    nor g1779(n1542 ,n469 ,n45);
    or g1780(n1903 ,n1466 ,n930);
    or g1781(n1986 ,n1355 ,n1666);
    or g1782(n1810 ,n1193 ,n878);
    not g1783(n188 ,n31[1]);
    nor g1784(n1057 ,n97 ,n818);
    nor g1785(n1185 ,n163 ,n61);
    nor g1786(n1510 ,n122 ,n43);
    dff g1787(.RN(n1), .SN(1'b1), .CK(n0), .D(n1832), .Q(n28[31]));
    not g1788(n507 ,n29[13]);
    nor g1789(n1658 ,n290 ,n49);
    or g1790(n2181 ,n1502 ,n1117);
    nor g1791(n1244 ,n490 ,n53);
    nor g1792(n1125 ,n619 ,n65);
    nor g1793(n1328 ,n208 ,n54);
    nor g1794(n1589 ,n283 ,n817);
    or g1795(n2183 ,n1509 ,n968);
    dff g1796(.RN(n1), .SN(1'b1), .CK(n0), .D(n1985), .Q(n34[11]));
    nor g1797(n1086 ,n92 ,n47);
    nor g1798(n851 ,n719 ,n45);
    nor g1799(n846 ,n640 ,n45);
    nor g1800(n1441 ,n424 ,n51);
    not g1801(n167 ,n28[22]);
    nor g1802(n1732 ,n122 ,n66);
    not g1803(n210 ,n29[15]);
    dff g1804(.RN(n1), .SN(1'b1), .CK(n0), .D(n1743), .Q(n34[19]));
    or g1805(n1964 ,n1331 ,n1675);
    nor g1806(n1694 ,n396 ,n63);
    dff g1807(.RN(n1), .SN(1'b1), .CK(n0), .D(n2089), .Q(n21[6]));
    xnor g1808(n677 ,n175 ,n105);
    or g1809(n2303 ,n2276 ,n2274);
    xnor g1810(n790 ,n352 ,n377);
    not g1811(n150 ,n24[16]);
    dff g1812(.RN(n1), .SN(1'b1), .CK(n0), .D(n2040), .Q(n33[17]));
    nor g1813(n915 ,n643 ,n55);
    not g1814(n380 ,n21[24]);
    not g1815(n317 ,n5[1]);
    nor g1816(n1284 ,n514 ,n53);
    nor g1817(n933 ,n711 ,n55);
    not g1818(n576 ,n11[28]);
    dff g1819(.RN(n1), .SN(1'b1), .CK(n0), .D(n1891), .Q(n31[19]));
    buf g1820(n12[12], n11[12]);
    dff g1821(.RN(n1), .SN(1'b1), .CK(n0), .D(n1837), .Q(n32[10]));
    nor g1822(n1150 ,n227 ,n65);
    or g1823(n1745 ,n1124 ,n829);
    dff g1824(.RN(n1), .SN(1'b1), .CK(n0), .D(n2148), .Q(n13[29]));
    or g1825(n1926 ,n1430 ,n1002);
    nor g1826(n1025 ,n73 ,n818);
    not g1827(n377 ,n30[1]);
    dff g1828(.RN(n1), .SN(1'b1), .CK(n0), .D(n1850), .Q(n28[25]));
    nor g1829(n1108 ,n363 ,n60);
    or g1830(n2048 ,n1393 ,n971);
    dff g1831(.RN(n1), .SN(1'b1), .CK(n0), .D(n1768), .Q(n11[22]));
    nor g1832(n1341 ,n516 ,n53);
    nor g1833(n1411 ,n177 ,n54);
    nor g1834(n1298 ,n565 ,n68);
    nor g1835(n884 ,n772 ,n59);
    nor g1836(n1312 ,n611 ,n68);
    not g1837(n226 ,n26[3]);
    nor g1838(n1166 ,n221 ,n816);
    nor g1839(n1605 ,n268 ,n52);
    nor g1840(n1608 ,n342 ,n52);
    nor g1841(n1324 ,n499 ,n57);
    not g1842(n590 ,n11[0]);
    dff g1843(.RN(n1), .SN(1'b1), .CK(n0), .D(n2132), .Q(n24[2]));
    not g1844(n64 ,n62);
    not g1845(n353 ,n21[1]);
    xnor g1846(n799 ,n77 ,n80);
    nor g1847(n1122 ,n92 ,n69);
    nor g1848(n1654 ,n337 ,n52);
    nor g1849(n1612 ,n325 ,n49);
    not g1850(n138 ,n26[21]);
    nor g1851(n1712 ,n420 ,n64);
    or g1852(n2165 ,n1486 ,n963);
    or g1853(n1886 ,n1266 ,n1106);
    dff g1854(.RN(n1), .SN(1'b1), .CK(n0), .D(n1815), .Q(n29[3]));
    or g1855(n626 ,n346 ,n71);
    dff g1856(.RN(n1), .SN(1'b1), .CK(n0), .D(n1897), .Q(n26[14]));
    not g1857(n245 ,n25[29]);
    dff g1858(.RN(n1), .SN(1'b1), .CK(n0), .D(n1943), .Q(n35[6]));
    nor g1859(n1363 ,n506 ,n54);
    dff g1860(.RN(n1), .SN(1'b1), .CK(n0), .D(n2036), .Q(n33[19]));
    not g1861(n2242 ,n24[18]);
    or g1862(n1743 ,n1308 ,n1683);
    nor g1863(n825 ,n725 ,n47);
    or g1864(n2037 ,n1126 ,n1568);
    nor g1865(n1632 ,n331 ,n817);
    not g1866(n450 ,n30[6]);
    or g1867(n1907 ,n1507 ,n969);
    dff g1868(.RN(n1), .SN(1'b1), .CK(n0), .D(n2018), .Q(n33[29]));
    or g1869(n2031 ,n1382 ,n1564);
    nor g1870(n991 ,n657 ,n69);
    not g1871(n434 ,n24[8]);
    dff g1872(.RN(n1), .SN(1'b1), .CK(n0), .D(n1746), .Q(n29[15]));
    xnor g1873(n703 ,n198 ,n135);
    xnor g1874(n756 ,n21[9] ,n24[9]);
    not g1875(n562 ,n12[30]);
    not g1876(n381 ,n21[7]);
    nor g1877(n1192 ,n109 ,n58);
    or g1878(n1837 ,n1225 ,n900);
    dff g1879(.RN(n1), .SN(1'b1), .CK(n0), .D(n1777), .Q(n11[16]));
    dff g1880(.RN(n1), .SN(1'b1), .CK(n0), .D(n2094), .Q(n24[25]));
    dff g1881(.RN(n1), .SN(1'b1), .CK(n0), .D(n2019), .Q(n33[28]));
    not g1882(n84 ,n21[31]);
    nor g1883(n1182 ,n104 ,n44);
    nor g1884(n917 ,n646 ,n55);
    xor g1885(n19[4] ,n21[4] ,n22[4]);
    xnor g1886(n768 ,n21[12] ,n24[12]);
    or g1887(n1955 ,n1061 ,n1584);
    nor g1888(n995 ,n635 ,n69);
    nor g1889(n1323 ,n531 ,n53);
    not g1890(n438 ,n30[29]);
    nor g1891(n1604 ,n298 ,n49);
    not g1892(n277 ,n6[0]);
    nor g1893(n1236 ,n546 ,n58);
    not g1894(n178 ,n29[7]);
    or g1895(n42 ,n27[0] ,n27[1]);
    not g1896(n604 ,n35[17]);
    nor g1897(n1219 ,n123 ,n67);
    nor g1898(n1078 ,n381 ,n818);
    nor g1899(n1588 ,n307 ,n52);
    xnor g1900(n776 ,n353 ,n399);
    dff g1901(.RN(n1), .SN(1'b1), .CK(n0), .D(n1844), .Q(n32[7]));
    or g1902(n2269 ,n2239 ,n21[28]);
    nor g1903(n1141 ,n594 ,n43);
    dff g1904(.RN(n1), .SN(1'b1), .CK(n0), .D(n2124), .Q(n24[7]));
    or g1905(n1763 ,n1142 ,n1528);
    nor g1906(n1731 ,n407 ,n66);
    or g1907(n2312 ,n2302 ,n2294);
    nor g1908(n1725 ,n151 ,n66);
    not g1909(n295 ,n4[5]);
    not g1910(n583 ,n11[19]);
    or g1911(n2154 ,n1482 ,n1658);
    or g1912(n1832 ,n1217 ,n1087);
    not g1913(n57 ,n60);
    or g1914(n1802 ,n1185 ,n872);
    not g1915(n425 ,n33[6]);
    not g1916(n202 ,n28[11]);
    or g1917(n2062 ,n1405 ,n831);
    nor g1918(n1599 ,n336 ,n49);
    or g1919(n2153 ,n1469 ,n1004);
    nor g1920(n1226 ,n121 ,n58);
    xnor g1921(n698 ,n183 ,n490);
    nor g1922(n1655 ,n303 ,n52);
    xnor g1923(n770 ,n82 ,n443);
    nor g1924(n1106 ,n372 ,n59);
    nor g1925(n1292 ,n242 ,n68);
    or g1926(n2082 ,n1419 ,n1607);
    nor g1927(n1194 ,n436 ,n67);
    nor g1928(n1034 ,n76 ,n51);
    dff g1929(.RN(n1), .SN(1'b1), .CK(n0), .D(n1875), .Q(n31[27]));
    or g1930(n1766 ,n1147 ,n1531);
    nor g1931(n1020 ,n350 ,n66);
    nor g1932(n1420 ,n617 ,n819);
    dff g1933(.RN(n1), .SN(1'b1), .CK(n0), .D(n1910), .Q(n35[27]));
    dff g1934(.RN(n1), .SN(1'b1), .CK(n0), .D(n823), .Q(n17[0]));
    nor g1935(n1709 ,n444 ,n56);
    not g1936(n86 ,n30[0]);
    not g1937(n148 ,n30[18]);
    or g1938(n1883 ,n1263 ,n921);
    dff g1939(.RN(n1), .SN(1'b1), .CK(n0), .D(n1929), .Q(n35[16]));
    not g1940(n391 ,n24[21]);
    not g1941(n115 ,n24[27]);
    or g1942(n2072 ,n1073 ,n951);
    dff g1943(.RN(n1), .SN(1'b1), .CK(n0), .D(n1903), .Q(n31[14]));
    xnor g1944(n708 ,n26[28] ,n33[24]);
    nor g1945(n958 ,n665 ,n56);
    not g1946(n43 ,n45);
    or g1947(n1999 ,n1238 ,n1699);
    not g1948(n586 ,n11[12]);
    buf g1949(n17[3], 1'b0);
    or g1950(n1996 ,n1242 ,n1697);
    not g1951(n619 ,n15[4]);
    nor g1952(n950 ,n804 ,n64);
    nor g1953(n1615 ,n272 ,n52);
    or g1954(n2163 ,n1484 ,n847);
    dff g1955(.RN(n1), .SN(1'b1), .CK(n0), .D(n1759), .Q(n15[3]));
    or g1956(n1882 ,n1260 ,n1104);
    not g1957(n441 ,n30[19]);
    nor g1958(n831 ,n782 ,n45);
    not g1959(n143 ,n33[5]);
    or g1960(n1978 ,n1352 ,n1687);
    nor g1961(n867 ,n633 ,n63);
    or g1962(n2316 ,n2310 ,n2308);
    dff g1963(.RN(n1), .SN(1'b1), .CK(n0), .D(n2146), .Q(n25[30]));
    dff g1964(.RN(n1), .SN(1'b1), .CK(n0), .D(n2140), .Q(n14[2]));
    or g1965(n2184 ,n1462 ,n1652);
    nor g1966(n1493 ,n599 ,n67);
    nor g1967(n1395 ,n103 ,n816);
    nor g1968(n1040 ,n79 ,n50);
    not g1969(n55 ,n54);
    or g1970(n2145 ,n1463 ,n835);
    buf g1971(n12[11], n11[11]);
    nor g1972(n842 ,n645 ,n45);
    xnor g1973(n720 ,n26[18] ,n33[14]);
    nor g1974(n1172 ,n218 ,n44);
    buf g1975(n17[5], 1'b0);
    nor g1976(n892 ,n769 ,n59);
    dff g1977(.RN(n1), .SN(1'b1), .CK(n0), .D(n2160), .Q(n13[22]));
    nor g1978(n46 ,n40 ,n37);
    nor g1979(n944 ,n790 ,n55);
    or g1980(n2157 ,n1477 ,n843);
    xnor g1981(n637 ,n475 ,n132);
    nor g1982(n850 ,n718 ,n48);
    dff g1983(.RN(n1), .SN(1'b1), .CK(n0), .D(n1994), .Q(n34[8]));
    nor g1984(n1460 ,n225 ,n43);
    not g1985(n287 ,n6[2]);
    nor g1986(n1164 ,n185 ,n61);
    or g1987(n1965 ,n1058 ,n1585);
    nor g1988(n909 ,n778 ,n60);
    or g1989(n1995 ,n1360 ,n1696);
    nor g1990(n1233 ,n550 ,n53);
    nor g1991(n1087 ,n84 ,n60);
    nor g1992(n989 ,n683 ,n69);
    dff g1993(.RN(n1), .SN(1'b1), .CK(n0), .D(n2176), .Q(n13[12]));
    not g1994(n504 ,n31[8]);
    nor g1995(n1307 ,n504 ,n53);
    not g1996(n386 ,n24[18]);
    xnor g1997(n664 ,n161 ,n522);
    or g1998(n2201 ,n1304 ,n1681);
    not g1999(n569 ,n13[0]);
    buf g2000(n14[7], n11[31]);
    nor g2001(n1297 ,n258 ,n819);
    nor g2002(n1696 ,n125 ,n64);
    nor g2003(n1400 ,n101 ,n44);
    or g2004(n2105 ,n1082 ,n1620);
    nor g2005(n845 ,n713 ,n48);
    nor g2006(n1262 ,n528 ,n57);
    buf g2007(n14[24], n11[24]);
    nor g2008(n1562 ,n565 ,n45);
    xnor g2009(n656 ,n192 ,n148);
    not g2010(n2256 ,n24[5]);
    nor g2011(n1437 ,n596 ,n819);
    not g2012(n320 ,n5[24]);
    xnor g2013(n675 ,n482 ,n497);
    not g2014(n162 ,n28[24]);
    not g2015(n222 ,n13[21]);
    not g2016(n337 ,n5[0]);
    dff g2017(.RN(n1), .SN(1'b1), .CK(n0), .D(n1771), .Q(n11[20]));
    nor g2018(n1634 ,n311 ,n49);
    not g2019(n2206 ,n2205);
    nor g2020(n1659 ,n306 ,n817);
    nor g2021(n1287 ,n444 ,n61);
    nor g2022(n1520 ,n551 ,n61);
    not g2023(n269 ,n5[19]);
    or g2024(n2069 ,n1409 ,n827);
    not g2025(n488 ,n35[1]);
    nor g2026(n1227 ,n193 ,n58);
    not g2027(n587 ,n11[30]);
    or g2028(n2009 ,n1213 ,n944);
    nor g2029(n1424 ,n426 ,n818);
    dff g2030(.RN(n1), .SN(1'b1), .CK(n0), .D(n1855), .Q(n28[23]));
    nor g2031(n1716 ,n104 ,n66);
    dff g2032(.RN(n1), .SN(1'b1), .CK(n0), .D(n2147), .Q(n13[30]));
    nor g2033(n1190 ,n114 ,n57);
    or g2034(n2113 ,n1035 ,n1627);
    buf g2035(n14[10], n11[10]);
    not g2036(n439 ,n32[12]);
    nor g2037(n1698 ,n450 ,n55);
    or g2038(n1958 ,n1059 ,n1583);
    nor g2039(n1069 ,n378 ,n818);
    or g2040(n1914 ,n1299 ,n933);
    dff g2041(.RN(n1), .SN(1'b1), .CK(n0), .D(n1965), .Q(n21[29]));
    nor g2042(n1573 ,n589 ,n48);
    nor g2043(n899 ,n754 ,n60);
    dff g2044(.RN(n1), .SN(1'b1), .CK(n0), .D(n1762), .Q(n15[2]));
    not g2045(n292 ,n5[26]);
    dff g2046(.RN(n1), .SN(1'b1), .CK(n0), .D(n1748), .Q(n13[0]));
    nor g2047(n905 ,n765 ,n59);
    nor g2048(n1512 ,n464 ,n66);
    or g2049(n2075 ,n1075 ,n1604);
    not g2050(n264 ,n4[29]);
    buf g2051(n16[7], n15[3]);
    not g2052(n400 ,n33[27]);
    dff g2053(.RN(n1), .SN(1'b1), .CK(n0), .D(n2008), .Q(n26[4]));
    not g2054(n468 ,n33[4]);
    or g2055(n2276 ,n2248 ,n2251);
    dff g2056(.RN(n1), .SN(1'b1), .CK(n0), .D(n2123), .Q(n24[8]));
    not g2057(n154 ,n33[22]);
    not g2058(n419 ,n24[29]);
    dff g2059(.RN(n1), .SN(1'b1), .CK(n0), .D(n1884), .Q(n28[13]));
    not g2060(n359 ,n21[13]);
    nor g2061(n1597 ,n310 ,n52);
    not g2062(n818 ,n49);
    or g2063(n2100 ,n1011 ,n1622);
    buf g2064(n12[15], n11[15]);
    nor g2065(n1650 ,n293 ,n52);
    nor g2066(n877 ,n738 ,n60);
    dff g2067(.RN(n1), .SN(1'b1), .CK(n0), .D(n1852), .Q(n28[24]));
    nor g2068(n1412 ,n602 ,n68);
    nor g2069(n871 ,n731 ,n64);
    dff g2070(.RN(n1), .SN(1'b1), .CK(n0), .D(n1883), .Q(n31[23]));
    nor g2071(n1509 ,n192 ,n61);
    dff g2072(.RN(n1), .SN(1'b1), .CK(n0), .D(n1915), .Q(n28[3]));
    not g2073(n90 ,n21[18]);
    dff g2074(.RN(n1), .SN(1'b1), .CK(n0), .D(n1992), .Q(n30[22]));
    not g2075(n541 ,n31[11]);
    nor g2076(n979 ,n801 ,n69);
    nor g2077(n1345 ,n403 ,n61);
    not g2078(n561 ,n35[18]);
    nor g2079(n1539 ,n435 ,n48);
    nor g2080(n2216 ,n2141 ,n2213);
    nor g2081(n978 ,n698 ,n69);
    dff g2082(.RN(n1), .SN(1'b1), .CK(n0), .D(n2201), .Q(n30[27]));
    or g2083(n2156 ,n1475 ,n842);
    not g2084(n216 ,n11[6]);
    or g2085(n2107 ,n1432 ,n1630);
    or g2086(n1962 ,n1338 ,n1674);
    or g2087(n1991 ,n1251 ,n1695);
    or g2088(n2318 ,n2314 ,n2309);
    not g2089(n303 ,n8[1]);
    not g2090(n130 ,n26[24]);
    or g2091(n1936 ,n1399 ,n990);
    not g2092(n65 ,n66);
    not g2093(n160 ,n28[19]);
    nor g2094(n1333 ,n505 ,n68);
    dff g2095(.RN(n1), .SN(1'b1), .CK(n0), .D(n2053), .Q(n33[9]));
    nor g2096(n1299 ,n541 ,n53);
    nor g2097(n1320 ,n257 ,n68);
    nor g2098(n874 ,n735 ,n59);
    or g2099(n1834 ,n1220 ,n1088);
    dff g2100(.RN(n1), .SN(1'b1), .CK(n0), .D(n2042), .Q(n30[8]));
    or g2101(n2223 ,n623 ,n2221);
    nor g2102(n1621 ,n280 ,n49);
    not g2103(n506 ,n34[4]);
    buf g2104(n12[13], n11[13]);
    dff g2105(.RN(n1), .SN(1'b1), .CK(n0), .D(n2214), .Q(n28[1]));
    not g2106(n367 ,n21[22]);
    nor g2107(n1513 ,n577 ,n816);
    nor g2108(n1726 ,n411 ,n66);
    dff g2109(.RN(n1), .SN(1'b1), .CK(n0), .D(n2137), .Q(n18[0]));
    dff g2110(.RN(n1), .SN(1'b1), .CK(n0), .D(n2200), .Q(n34[18]));
    not g2111(n445 ,n32[23]);
    not g2112(n183 ,n34[31]);
    buf g2113(n14[14], n11[14]);
    dff g2114(.RN(n1), .SN(1'b1), .CK(n0), .D(n1802), .Q(n29[6]));
    dff g2115(.RN(n1), .SN(1'b1), .CK(n0), .D(n2039), .Q(n21[16]));
    nor g2116(n1413 ,n570 ,n68);
    not g2117(n431 ,n30[7]);
    dff g2118(.RN(n1), .SN(1'b1), .CK(n0), .D(n1967), .Q(n34[24]));
    dff g2119(.RN(n1), .SN(1'b1), .CK(n0), .D(n1814), .Q(n32[23]));
    or g2120(n2140 ,n1456 ,n1016);
    nor g2121(n1378 ,n397 ,n816);
    nor g2122(n2141 ,n27[2] ,n1281);
    or g2123(n1898 ,n1050 ,n928);
    or g2124(n2304 ,n2282 ,n2281);
    nor g2125(n1648 ,n333 ,n49);
    or g2126(n2322 ,n2320 ,n2321);
    or g2127(n2279 ,n2250 ,n24[24]);
    not g2128(n104 ,n33[28]);
    not g2129(n218 ,n11[5]);
    nor g2130(n1422 ,n419 ,n51);
    not g2131(n107 ,n26[26]);
    nor g2132(n1488 ,n545 ,n58);
    not g2133(n49 ,n51);
    not g2134(n205 ,n34[25]);
    not g2135(n286 ,n6[3]);
    dff g2136(.RN(n1), .SN(1'b1), .CK(n0), .D(n2117), .Q(n29[31]));
    xnor g2137(n791 ,n77 ,n379);
    nor g2138(n1614 ,n316 ,n49);
    nor g2139(n1067 ,n359 ,n50);
    xnor g2140(n742 ,n21[23] ,n24[23]);
    or g2141(n2021 ,n1175 ,n1551);
    nor g2142(n1633 ,n335 ,n817);
    or g2143(n2007 ,n1366 ,n1702);
    nor g2144(n1736 ,n142 ,n66);
    nor g2145(n1430 ,n604 ,n819);
    nor g2146(n1487 ,n584 ,n44);
    nor g2147(n1381 ,n501 ,n68);
    not g2148(n366 ,n21[4]);
    nor g2149(n1012 ,n348 ,n50);
    nor g2150(n1083 ,n95 ,n48);
    nor g2151(n1151 ,n568 ,n44);
    or g2152(n2056 ,n1067 ,n1660);
    nor g2153(n1518 ,n616 ,n816);
    not g2154(n585 ,n26[0]);
    nor g2155(n1232 ,n204 ,n57);
    nor g2156(n1386 ,n151 ,n44);
    nor g2157(n1357 ,n186 ,n53);
    nor g2158(n1107 ,n378 ,n60);
    xnor g2159(n695 ,n26[15] ,n33[11]);
    xnor g2160(n659 ,n551 ,n414);
    nor g2161(n1704 ,n118 ,n64);
    or g2162(n1829 ,n1216 ,n895);
    or g2163(n2302 ,n2287 ,n2271);
    dff g2164(.RN(n1), .SN(1'b1), .CK(n0), .D(n1811), .Q(n32[25]));
    or g2165(n1900 ,n1284 ,n929);
    or g2166(n2010 ,n1369 ,n1703);
    buf g2167(n16[4], n15[0]);
    dff g2168(.RN(n1), .SN(1'b1), .CK(n0), .D(n2026), .Q(n21[18]));
    nor g2169(n860 ,n811 ,n47);
    not g2170(n430 ,n33[25]);
    nor g2171(n1142 ,n552 ,n46);
    nor g2172(n1139 ,n576 ,n43);
    or g2173(n2127 ,n1446 ,n1648);
    xnor g2174(n738 ,n21[27] ,n24[27]);
    nor g2175(n856 ,n679 ,n47);
    nor g2176(n1459 ,n563 ,n819);
    nor g2177(n1552 ,n427 ,n47);
    nor g2178(n1265 ,n521 ,n53);
    nor g2179(n1581 ,n282 ,n49);
    nor g2180(n1091 ,n87 ,n60);
    nor g2181(n1561 ,n258 ,n48);
    nor g2182(n1567 ,n596 ,n48);
    not g2183(n462 ,n26[15]);
    nor g2184(n1547 ,n111 ,n45);
    dff g2185(.RN(n1), .SN(1'b1), .CK(n0), .D(n1979), .Q(n30[25]));
    not g2186(n355 ,n21[0]);
    buf g2187(n14[13], n11[13]);
    nor g2188(n1550 ,n99 ,n45);
    nor g2189(n1213 ,n476 ,n53);
    or g2190(n2314 ,n2305 ,n2301);
    nor g2191(n1342 ,n438 ,n61);
    dff g2192(.RN(n1), .SN(1'b1), .CK(n0), .D(n1941), .Q(n31[4]));
    nor g2193(n1683 ,n441 ,n55);
    dff g2194(.RN(n1), .SN(1'b1), .CK(n0), .D(n1758), .Q(n29[13]));
    not g2195(n523 ,n31[28]);
    or g2196(n2013 ,n1370 ,n1704);
    or g2197(n1985 ,n1356 ,n1692);
    xnor g2198(n692 ,n529 ,n514);
    dff g2199(.RN(n1), .SN(1'b1), .CK(n0), .D(n1879), .Q(n28[15]));
    nor g2200(n1583 ,n322 ,n52);
    xnor g2201(n733 ,n21[31] ,n24[31]);
    dff g2202(.RN(n1), .SN(1'b1), .CK(n0), .D(n2161), .Q(n13[21]));
    not g2203(n251 ,n11[14]);
    buf g2204(n12[20], n11[20]);
    nor g2205(n855 ,n695 ,n45);
    or g2206(n2085 ,n1422 ,n1611);
    dff g2207(.RN(n1), .SN(1'b1), .CK(n0), .D(n1970), .Q(n21[28]));
    nor g2208(n1196 ,n390 ,n43);
    nor g2209(n1490 ,n417 ,n44);
    or g2210(n1875 ,n1273 ,n917);
    dff g2211(.RN(n1), .SN(1'b1), .CK(n0), .D(n1009), .Q(n17[2]));
    nor g2212(n997 ,n681 ,n69);
    nor g2213(n1295 ,n187 ,n53);
    not g2214(n306 ,n4[12]);
    dff g2215(.RN(n1), .SN(1'b1), .CK(n0), .D(n1756), .Q(n11[30]));
    not g2216(n408 ,n32[30]);
    dff g2217(.RN(n1), .SN(1'b1), .CK(n0), .D(n2195), .Q(n13[2]));
    or g2218(n2295 ,n2272 ,n2270);
    or g2219(n39 ,n346 ,n27[0]);
    nor g2220(n1527 ,n436 ,n47);
    nor g2221(n1742 ,n593 ,n65);
    nor g2222(n1239 ,n530 ,n58);
    dff g2223(.RN(n1), .SN(1'b1), .CK(n0), .D(n1745), .Q(n13[1]));
    not g2224(n591 ,n11[1]);
    nor g2225(n1464 ,n247 ,n44);
    nor g2226(n1296 ,n536 ,n53);
    nor g2227(n1611 ,n304 ,n817);
    not g2228(n254 ,n13[11]);
    nor g2229(n1526 ,n128 ,n47);
    not g2230(n457 ,n30[21]);
    nor g2231(n1286 ,n117 ,n61);
    not g2232(n123 ,n26[23]);
    or g2233(n2213 ,n70 ,n2199);
    not g2234(n351 ,n22[5]);
    not g2235(n186 ,n34[10]);
    nor g2236(n1336 ,n395 ,n61);
    not g2237(n176 ,n29[28]);
    nor g2238(n881 ,n773 ,n60);
    xnor g2239(n773 ,n21[24] ,n24[24]);
    nor g2240(n1314 ,n248 ,n68);
    or g2241(n1945 ,n1326 ,n994);
    not g2242(n101 ,n33[8]);
    or g2243(n2025 ,n1160 ,n1562);
    or g2244(n1807 ,n1186 ,n1716);
    dff g2245(.RN(n1), .SN(1'b1), .CK(n0), .D(n1931), .Q(n31[7]));
    dff g2246(.RN(n1), .SN(1'b1), .CK(n0), .D(n2119), .Q(n21[2]));
    not g2247(n817 ,n818);
    or g2248(n2093 ,n1022 ,n1615);
    nor g2249(n1249 ,n527 ,n57);
    xnor g2250(n810 ,n507 ,n152);
    not g2251(n505 ,n35[0]);
    not g2252(n473 ,n29[17]);
    or g2253(n1753 ,n1125 ,n1026);
    or g2254(n1846 ,n1046 ,n905);
    nor g2255(n1266 ,n474 ,n57);
    or g2256(n1746 ,n1123 ,n973);
    nor g2257(n1586 ,n301 ,n49);
    or g2258(n2197 ,n1350 ,n1667);
    nor g2259(n1367 ,n99 ,n67);
    not g2260(n79 ,n18[0]);
    or g2261(n1828 ,n1215 ,n893);
    xnor g2262(n794 ,n78 ,n373);
    not g2263(n248 ,n35[13]);
    nor g2264(n1044 ,n85 ,n51);
    xnor g2265(n696 ,n542 ,n121);
    not g2266(n532 ,n29[29]);
    dff g2267(.RN(n1), .SN(1'b1), .CK(n0), .D(n2170), .Q(n13[15]));
    or g2268(n2308 ,n2296 ,n2292);
    or g2269(n2080 ,n1410 ,n1122);
    not g2270(n82 ,n36[2]);
    or g2271(n1839 ,n1219 ,n1721);
    dff g2272(.RN(n1), .SN(1'b1), .CK(n0), .D(n1753), .Q(n15[4]));
    nor g2273(n1556 ,n585 ,n48);
    dff g2274(.RN(n1), .SN(1'b1), .CK(n0), .D(n2215), .Q(n28[0]));
    or g2275(n2005 ,n1062 ,n1592);
    not g2276(n410 ,n26[30]);
    nor g2277(n824 ,n729 ,n45);
    nor g2278(n1421 ,n155 ,n51);
    nor g2279(n894 ,n751 ,n59);
    or g2280(n2150 ,n1468 ,n839);
    not g2281(n589 ,n35[11]);
    dff g2282(.RN(n1), .SN(1'b1), .CK(n0), .D(n2041), .Q(n33[16]));
    or g2283(n41 ,n70 ,n27[2]);
    or g2284(n1940 ,n1321 ,n1005);
    dff g2285(.RN(n1), .SN(1'b1), .CK(n0), .D(n2074), .Q(n21[9]));
    dff g2286(.RN(n1), .SN(1'b1), .CK(n0), .D(n1969), .Q(n34[23]));
    not g2287(n157 ,n29[12]);
    or g2288(n1858 ,n1052 ,n911);
    nor g2289(n1174 ,n615 ,n44);
    nor g2290(n1092 ,n371 ,n59);
    nor g2291(n1001 ,n673 ,n69);
    not g2292(n545 ,n28[4]);
    not g2293(n376 ,n32[4]);
    dff g2294(.RN(n1), .SN(1'b1), .CK(n0), .D(n1960), .Q(n34[27]));
    nor g2295(n1310 ,n477 ,n54);
    xnor g2296(n766 ,n26[5] ,n33[1]);
    not g2297(n300 ,n5[12]);
    or g2298(n1819 ,n1204 ,n885);
    xnor g2299(n651 ,n539 ,n461);
    dff g2300(.RN(n1), .SN(1'b1), .CK(n0), .D(n1838), .Q(n28[29]));
    nor g2301(n1137 ,n581 ,n43);
    xnor g2302(n706 ,n26[30] ,n33[26]);
    not g2303(n156 ,n28[29]);
    dff g2304(.RN(n1), .SN(1'b1), .CK(n0), .D(n1854), .Q(n32[2]));
    not g2305(n256 ,n12[31]);
    or g2306(n2191 ,n1518 ,n860);
    not g2307(n189 ,n31[25]);
    or g2308(n1931 ,n1418 ,n937);
    nor g2309(n928 ,n659 ,n56);
    or g2310(n2217 ,n70 ,n2212);
    dff g2311(.RN(n1), .SN(1'b1), .CK(n0), .D(n1781), .Q(n11[14]));
    or g2312(n625 ,n182 ,n7[3]);
    not g2313(n333 ,n5[5]);
    nor g2314(n1167 ,n214 ,n46);
    not g2315(n396 ,n32[22]);
    not g2316(n271 ,n4[11]);
    or g2317(n1988 ,n1343 ,n1668);
    nor g2318(n1075 ,n369 ,n51);
    xnor g2319(n644 ,n176 ,n403);
    or g2320(n2131 ,n1339 ,n941);
    nor g2321(n1148 ,n388 ,n61);
    not g2322(n565 ,n35[25]);
    dff g2323(.RN(n1), .SN(1'b1), .CK(n0), .D(n1937), .Q(n31[5]));
    dff g2324(.RN(n1), .SN(1'b1), .CK(n0), .D(n1973), .Q(n30[28]));
    or g2325(n1992 ,n1252 ,n1694);
    nor g2326(n879 ,n774 ,n59);
    buf g2327(n12[0], n11[28]);
    nor g2328(n864 ,n628 ,n63);
    xnor g2329(n741 ,n172 ,n357);
    nor g2330(n1109 ,n360 ,n60);
    dff g2331(.RN(n1), .SN(1'b1), .CK(n0), .D(n2047), .Q(n33[13]));
    or g2332(n1816 ,n1202 ,n1719);
    dff g2333(.RN(n1), .SN(1'b1), .CK(n0), .D(n1749), .Q(n12[31]));
    or g2334(n1952 ,n1330 ,n913);
    or g2335(n2124 ,n1444 ,n1644);
    or g2336(n2074 ,n1074 ,n1603);
    xnor g2337(n727 ,n352 ,n353);
    nor g2338(n866 ,n699 ,n64);
    nor g2339(n1429 ,n391 ,n50);
    nor g2340(n1643 ,n266 ,n52);
    or g2341(n2283 ,n2247 ,n24[21]);
    xnor g2342(n750 ,n499 ,n83);
    nor g2343(n1104 ,n361 ,n60);
    dff g2344(.RN(n1), .SN(1'b1), .CK(n0), .D(n2152), .Q(n29[25]));
    not g2345(n236 ,n11[16]);
    or g2346(n1933 ,n1314 ,n989);
    dff g2347(.RN(n1), .SN(1'b1), .CK(n0), .D(n2011), .Q(n34[0]));
    nor g2348(n1073 ,n373 ,n61);
    nor g2349(n873 ,n734 ,n59);
    buf g2350(n12[16], n11[16]);
    or g2351(n1969 ,n1322 ,n1678);
    nor g2352(n921 ,n650 ,n55);
    not g2353(n466 ,n33[16]);
    or g2354(n1971 ,n1323 ,n1679);
    nor g2355(n1203 ,n125 ,n58);
    xnor g2356(n654 ,n548 ,n147);
    not g2357(n547 ,n28[2]);
    nor g2358(n1479 ,n252 ,n816);
    nor g2359(n1260 ,n191 ,n57);
    nor g2360(n1283 ,n469 ,n67);
    dff g2361(.RN(n1), .SN(1'b1), .CK(n0), .D(n2129), .Q(n21[0]));
    or g2362(n1761 ,n1141 ,n1527);
    nor g2363(n906 ,n758 ,n60);
    or g2364(n37 ,n347 ,n27[1]);
    or g2365(n1821 ,n1205 ,n887);
    or g2366(n1966 ,n1332 ,n1735);
    dff g2367(.RN(n1), .SN(1'b1), .CK(n0), .D(n1856), .Q(n32[1]));
    not g2368(n128 ,n26[28]);
    or g2369(n2046 ,n1391 ,n1571);
    nor g2370(n1369 ,n416 ,n61);
    nor g2371(n2211 ,n182 ,n2206);
    not g2372(n526 ,n29[11]);
    nor g2373(n1560 ,n242 ,n48);
    not g2374(n522 ,n31[23]);
    nor g2375(n67 ,n40 ,n39);
    nor g2376(n1463 ,n228 ,n43);
    not g2377(n237 ,n11[13]);
    not g2378(n478 ,n29[1]);
    dff g2379(.RN(n1), .SN(1'b1), .CK(n0), .D(n1964), .Q(n30[30]));
    not g2380(n339 ,n9[2]);
    dff g2381(.RN(n1), .SN(1'b1), .CK(n0), .D(n2097), .Q(n22[4]));
    nor g2382(n1680 ,n457 ,n55);
    nor g2383(n1212 ,n118 ,n57);
    nor g2384(n1494 ,n574 ,n44);
    xnor g2385(n730 ,n169 ,n379);
    not g2386(n225 ,n14[0]);
    not g2387(n262 ,n13[23]);
    not g2388(n460 ,n24[19]);
    nor g2389(n1018 ,n72 ,n66);
    not g2390(n89 ,n33[0]);
    nor g2391(n1155 ,n610 ,n46);
    nor g2392(n51 ,n41 ,n42);
    or g2393(n2038 ,n1148 ,n1711);
    dff g2394(.RN(n1), .SN(1'b1), .CK(n0), .D(n1763), .Q(n11[26]));
    nor g2395(n1657 ,n302 ,n52);
    or g2396(n2146 ,n1458 ,n1657);
    or g2397(n2267 ,n2252 ,n24[13]);
    buf g2398(n17[7], 1'b0);
    dff g2399(.RN(n1), .SN(1'b1), .CK(n0), .D(n1866), .Q(n31[31]));
    not g2400(n87 ,n21[27]);
    or g2401(n1860 ,n1032 ,n1580);
    nor g2402(n1388 ,n226 ,n65);
    nor g2403(n1666 ,n445 ,n63);
    nor g2404(n1211 ,n124 ,n57);
    or g2405(n1919 ,n1472 ,n984);
    not g2406(n219 ,n13[4]);
    or g2407(n2012 ,n1063 ,n1593);
    dff g2408(.RN(n1), .SN(1'b1), .CK(n0), .D(n2092), .Q(n24[26]));
    not g2409(n595 ,n35[31]);
    not g2410(n243 ,n15[6]);
    dff g2411(.RN(n1), .SN(1'b1), .CK(n0), .D(n1808), .Q(n32[27]));
    or g2412(n2263 ,n21[9] ,n21[8]);
    or g2413(n1783 ,n1162 ,n1543);
    xnor g2414(n635 ,n496 ,n164);
    or g2415(n2278 ,n2232 ,n21[18]);
    or g2416(n1932 ,n1312 ,n988);
    nor g2417(n1178 ,n178 ,n61);
    or g2418(n2178 ,n1503 ,n855);
    nor g2419(n1606 ,n305 ,n49);
    dff g2420(.RN(n1), .SN(1'b1), .CK(n0), .D(n1766), .Q(n11[23]));
    nor g2421(n1127 ,n569 ,n44);
    dff g2422(.RN(n1), .SN(1'b1), .CK(n0), .D(n2099), .Q(n24[22]));
    dff g2423(.RN(n1), .SN(1'b1), .CK(n0), .D(n1993), .Q(n26[6]));
    dff g2424(.RN(n1), .SN(1'b1), .CK(n0), .D(n1901), .Q(n28[6]));
    xnor g2425(n792 ,n79 ,n89);
    nor g2426(n1101 ,n94 ,n59);
    xnor g2427(n712 ,n546 ,n445);
    not g2428(n71 ,n27[2]);
    nor g2429(n1446 ,n149 ,n50);
    dff g2430(.RN(n1), .SN(1'b1), .CK(n0), .D(n1889), .Q(n28[11]));
    or g2431(n2286 ,n2245 ,n2238);
    buf g2432(n12[3], n11[31]);
    xnor g2433(n711 ,n526 ,n392);
    nor g2434(n1285 ,n492 ,n57);
    nor g2435(n1645 ,n299 ,n52);
    nor g2436(n1456 ,n582 ,n43);
    xnor g2437(n717 ,n530 ,n125);
    nor g2438(n1703 ,n124 ,n63);
    dff g2439(.RN(n1), .SN(1'b1), .CK(n0), .D(n2098), .Q(n24[23]));
    nor g2440(n1032 ,n78 ,n818);
    or g2441(n2317 ,n2311 ,n2312);
    xnor g2442(n758 ,n21[5] ,n24[5]);
    nor g2443(n932 ,n764 ,n55);
    dff g2444(.RN(n1), .SN(1'b1), .CK(n0), .D(n1817), .Q(n32[22]));
    not g2445(n557 ,n13[25]);
    nor g2446(n1516 ,n556 ,n65);
    nor g2447(n1695 ,n388 ,n56);
    or g2448(n2014 ,n1196 ,n1557);
    dff g2449(.RN(n1), .SN(1'b1), .CK(n0), .D(n1750), .Q(n12[30]));
    or g2450(n1920 ,n1291 ,n1732);
    xor g2451(n19[2] ,n21[2] ,n22[2]);
    or g2452(n2102 ,n1081 ,n1613);
    dff g2453(.RN(n1), .SN(1'b1), .CK(n0), .D(n1868), .Q(n28[19]));
    nor g2454(n945 ,n789 ,n56);
    not g2455(n194 ,n29[30]);
    nor g2456(n826 ,n710 ,n47);
    nor g2457(n1396 ,n409 ,n44);
    not g2458(n383 ,n21[21]);
    or g2459(n38 ,n347 ,n346);
    not g2460(n307 ,n4[26]);
    not g2461(n2240 ,n24[26]);
    xnor g2462(n643 ,n532 ,n438);
    nor g2463(n965 ,n637 ,n63);
    nor g2464(n2203 ,n625 ,n1030);
    nor g2465(n904 ,n757 ,n59);
    not g2466(n612 ,n35[8]);
    nor g2467(n1123 ,n210 ,n62);
    not g2468(n492 ,n28[6]);
    dff g2469(.RN(n1), .SN(1'b1), .CK(n0), .D(n1860), .Q(n23[2]));
    nor g2470(n1729 ,n454 ,n66);
    or g2471(n1880 ,n1259 ,n919);
    nor g2472(n1385 ,n134 ,n62);
    nor g2473(n1544 ,n412 ,n45);
    dff g2474(.RN(n1), .SN(1'b1), .CK(n0), .D(n2093), .Q(n22[5]));
    or g2475(n1977 ,n1055 ,n1588);
    or g2476(n1890 ,n1270 ,n1108);
    or g2477(n2090 ,n1077 ,n952);
    or g2478(n2095 ,n1349 ,n974);
    or g2479(n1944 ,n1376 ,n946);
    xnor g2480(n778 ,n356 ,n139);
    buf g2481(n14[26], n11[26]);
    not g2482(n136 ,n32[19]);
    or g2483(n1857 ,n1237 ,n1096);
    xnor g2484(n704 ,n538 ,n422);
    xnor g2485(n813 ,n527 ,n124);
    or g2486(n1974 ,n1346 ,n1682);
    or g2487(n2173 ,n1498 ,n965);
    nor g2488(n1538 ,n405 ,n45);
    xnor g2489(n661 ,n515 ,n118);
    or g2490(n2106 ,n1431 ,n1628);
    dff g2491(.RN(n1), .SN(1'b1), .CK(n0), .D(n1950), .Q(n35[2]));
    nor g2492(n1081 ,n91 ,n818);
    not g2493(n315 ,n9[6]);
    nor g2494(n1662 ,n132 ,n64);
    or g2495(n1867 ,n1246 ,n914);
    nor g2496(n830 ,n780 ,n45);
    not g2497(n278 ,n9[1]);
    dff g2498(.RN(n1), .SN(1'b1), .CK(n0), .D(n2068), .Q(n21[10]));
    nor g2499(n980 ,n721 ,n69);
    or g2500(n2290 ,n2234 ,n2228);
    nor g2501(n1630 ,n319 ,n49);
    dff g2502(.RN(n1), .SN(1'b1), .CK(n0), .D(n2183), .Q(n29[18]));
    or g2503(n1752 ,n1130 ,n864);
    not g2504(n78 ,n23[2]);
    not g2505(n2258 ,n24[28]);
    nor g2506(n2207 ,n27[1] ,n2203);
    dff g2507(.RN(n1), .SN(1'b1), .CK(n0), .D(n2159), .Q(n13[23]));
    nor g2508(n875 ,n736 ,n63);
    or g2509(n2260 ,n2242 ,n24[19]);
    not g2510(n484 ,n28[8]);
    nor g2511(n1711 ,n121 ,n63);
    or g2512(n2299 ,n2284 ,n2283);
    nor g2513(n1601 ,n271 ,n49);
    not g2514(n192 ,n29[18]);
    nor g2515(n1481 ,n222 ,n43);
    nor g2516(n1555 ,n573 ,n45);
    nor g2517(n1590 ,n330 ,n49);
    dff g2518(.RN(n1), .SN(1'b1), .CK(n0), .D(n1949), .Q(n26[9]));
    dff g2519(.RN(n1), .SN(1'b1), .CK(n0), .D(n1851), .Q(n32[4]));
    not g2520(n533 ,n31[10]);
    dff g2521(.RN(n1), .SN(1'b1), .CK(n0), .D(n2102), .Q(n21[5]));
    not g2522(n319 ,n5[18]);
    nor g2523(n1535 ,n458 ,n48);
    dff g2524(.RN(n1), .SN(1'b1), .CK(n0), .D(n1881), .Q(n31[24]));
    xnor g2525(n753 ,n21[13] ,n24[13]);
    nor g2526(n1274 ,n481 ,n53);
    not g2527(n252 ,n13[22]);
    or g2528(n2164 ,n1487 ,n848);
    not g2529(n588 ,n10[0]);
    dff g2530(.RN(n1), .SN(1'b1), .CK(n0), .D(n1963), .Q(n34[29]));
    nor g2531(n1105 ,n359 ,n59);
    or g2532(n1838 ,n1224 ,n1089);
    or g2533(n1870 ,n1248 ,n915);
    nor g2534(n983 ,n666 ,n69);
    nor g2535(n1027 ,n75 ,n66);
    nor g2536(n1186 ,n128 ,n67);
    xnor g2537(n648 ,n184 ,n117);
    nor g2538(n888 ,n746 ,n60);
    xnor g2539(n798 ,n73 ,n376);
    or g2540(n2166 ,n1489 ,n849);
    or g2541(n1825 ,n1211 ,n891);
    buf g2542(n12[1], n11[29]);
    xnor g2543(n722 ,n26[17] ,n33[13]);
    not g2544(n187 ,n34[17]);
    dff g2545(.RN(n1), .SN(1'b1), .CK(n0), .D(n2067), .Q(n30[3]));
    xnor g2546(n754 ,n21[11] ,n24[11]);
    or g2547(n1881 ,n1261 ,n920);
    nor g2548(n1598 ,n289 ,n52);
    or g2549(n2142 ,n1457 ,n1014);
    not g2550(n172 ,n28[3]);
    nor g2551(n949 ,n798 ,n64);
    nor g2552(n1159 ,n251 ,n43);
    xor g2553(n20[3] ,n23[3] ,n24[3]);
    nor g2554(n1214 ,n145 ,n57);
    not g2555(n196 ,n34[8]);
    or g2556(n2043 ,n1483 ,n1578);
    dff g2557(.RN(n1), .SN(1'b1), .CK(n0), .D(n1942), .Q(n35[7]));
    dff g2558(.RN(n1), .SN(1'b1), .CK(n0), .D(n1898), .Q(n31[16]));
    or g2559(n1877 ,n1256 ,n918);
    dff g2560(.RN(n1), .SN(1'b1), .CK(n0), .D(n1798), .Q(n11[1]));
    or g2561(n2222 ,n622 ,n2220);
    dff g2562(.RN(n1), .SN(1'b1), .CK(n0), .D(n2186), .Q(n13[7]));
    nor g2563(n893 ,n750 ,n64);
    nor g2564(n1515 ,n473 ,n61);
    not g2565(n242 ,n35[28]);
    not g2566(n327 ,n5[4]);
    or g2567(n2138 ,n1455 ,n1015);
    nor g2568(n1715 ,n100 ,n66);
    or g2569(n2065 ,n1069 ,n1601);
    or g2570(n2092 ,n1424 ,n1616);
    nor g2571(n990 ,n691 ,n69);
    not g2572(n80 ,n21[3]);
    not g2573(n66 ,n67);
    nor g2574(n1368 ,n126 ,n51);
    dff g2575(.RN(n1), .SN(1'b1), .CK(n0), .D(n1886), .Q(n28[12]));
    dff g2576(.RN(n1), .SN(1'b1), .CK(n0), .D(n2010), .Q(n30[17]));
    not g2577(n340 ,n5[15]);
    dff g2578(.RN(n1), .SN(1'b1), .CK(n0), .D(n1902), .Q(n35[31]));
    dff g2579(.RN(n1), .SN(1'b1), .CK(n0), .D(n1805), .Q(n29[5]));
    buf g2580(n14[21], n11[21]);
    not g2581(n2232 ,n21[19]);
    dff g2582(.RN(n1), .SN(1'b1), .CK(n0), .D(n1778), .Q(n11[15]));
    not g2583(n349 ,n22[0]);
    nor g2584(n1248 ,n199 ,n53);
    or g2585(n1861 ,n1239 ,n1097);
    xnor g2586(n781 ,n73 ,n519);
    buf g2587(n12[17], n11[17]);
    nor g2588(n985 ,n701 ,n69);
    not g2589(n2247 ,n24[20]);
    not g2590(n223 ,n35[20]);
    nor g2591(n1566 ,n223 ,n48);
    nor g2592(n1474 ,n488 ,n68);
    nor g2593(n1036 ,n356 ,n818);
    xnor g2594(n762 ,n95 ,n390);
    nor g2595(n1543 ,n401 ,n45);
    dff g2596(.RN(n1), .SN(1'b1), .CK(n0), .D(n2082), .Q(n24[31]));
    not g2597(n139 ,n24[2]);
    nor g2598(n1180 ,n591 ,n44);
    not g2599(n515 ,n28[16]);
    nor g2600(n1577 ,n572 ,n45);
    or g2601(n2188 ,n1506 ,n1118);
    nor g2602(n1033 ,n352 ,n818);
    or g2603(n1913 ,n1298 ,n981);
    or g2604(n2162 ,n1480 ,n962);
    nor g2605(n1613 ,n295 ,n49);
    dff g2606(.RN(n1), .SN(1'b1), .CK(n0), .D(n2138), .Q(n14[3]));
    xnor g2607(n800 ,n78 ,n356);
    not g2608(n96 ,n33[1]);
    not g2609(n233 ,n11[7]);
    nor g2610(n1145 ,n564 ,n44);
    nor g2611(n925 ,n655 ,n55);
    nor g2612(n1303 ,n412 ,n65);
    dff g2613(.RN(n1), .SN(1'b1), .CK(n0), .D(n1984), .Q(n34[12]));
    xnor g2614(n690 ,n167 ,n396);
    buf g2615(n15[12], 1'b0);
    nor g2616(n882 ,n741 ,n64);
    nor g2617(n1063 ,n383 ,n51);
    dff g2618(.RN(n1), .SN(1'b1), .CK(n0), .D(n1761), .Q(n11[27]));
    xnor g2619(n734 ,n21[30] ,n24[30]);
    nor g2620(n1373 ,n100 ,n816);
    nor g2621(n929 ,n660 ,n56);
    nor g2622(n1243 ,n160 ,n57);
    not g2623(n324 ,n3[31]);
    dff g2624(.RN(n1), .SN(1'b1), .CK(n0), .D(n2122), .Q(n24[9]));
    or g2625(n2104 ,n1374 ,n1626);
    not g2626(n184 ,n29[25]);
    xnor g2627(n725 ,n26[14] ,n33[10]);
    or g2628(n1798 ,n1180 ,n1555);
    nor g2629(n1628 ,n269 ,n49);
    or g2630(n40 ,n71 ,n70);
    or g2631(n1749 ,n1128 ,n1523);
    nor g2632(n1156 ,n236 ,n43);
    or g2633(n1972 ,n1310 ,n1680);
    nor g2634(n998 ,n678 ,n69);
    nor g2635(n1644 ,n312 ,n49);
    or g2636(n1808 ,n1191 ,n877);
    dff g2637(.RN(n1), .SN(1'b1), .CK(n0), .D(n2081), .Q(n21[7]));
    not g2638(n608 ,n35[10]);
    or g2639(n2079 ,n1079 ,n953);
    nor g2640(n1331 ,n432 ,n61);
    or g2641(n1809 ,n1192 ,n879);
    not g2642(n209 ,n28[31]);
    not g2643(n362 ,n32[6]);
    dff g2644(.RN(n1), .SN(1'b1), .CK(n0), .D(n2127), .Q(n24[5]));
    or g2645(n2044 ,n1065 ,n1599);
    dff g2646(.RN(n1), .SN(1'b1), .CK(n0), .D(n1924), .Q(n26[11]));
    or g2647(n1983 ,n1287 ,n1689);
    nor g2648(n1046 ,n362 ,n57);
    buf g2649(n16[8], n15[4]);
    xnor g2650(n678 ,n506 ,n177);
    nor g2651(n1557 ,n595 ,n48);
    xnor g2652(n686 ,n476 ,n188);
    xnor g2653(n760 ,n478 ,n377);
    nor g2654(n1574 ,n608 ,n47);
    not g2655(n70 ,n2);
    nor g2656(n1727 ,n447 ,n66);
    nor g2657(n1699 ,n389 ,n56);
    nor g2658(n1278 ,n484 ,n57);
    nor g2659(n1210 ,n130 ,n67);
    dff g2660(.RN(n1), .SN(1'b1), .CK(n0), .D(n1888), .Q(n31[20]));
    or g2661(n1831 ,n1218 ,n896);
    not g2662(n476 ,n34[1]);
    nor g2663(n1128 ,n256 ,n43);
    dff g2664(.RN(n1), .SN(1'b1), .CK(n0), .D(n2027), .Q(n33[24]));
    xnor g2665(n687 ,n26[11] ,n33[7]);
    not g2666(n368 ,n32[2]);
    or g2667(n1897 ,n1264 ,n1729);
    or g2668(n1934 ,n1316 ,n1001);
    xnor g2669(n653 ,n26[31] ,n33[27]);
    or g2670(n1790 ,n1168 ,n870);
    nor g2671(n1723 ,n470 ,n66);
    not g2672(n230 ,n12[28]);
    or g2673(n2119 ,n1036 ,n1634);
    not g2674(n370 ,n32[1]);
    nor g2675(n1718 ,n451 ,n66);
    not g2676(n45 ,n46);
    nor g2677(n1465 ,n495 ,n61);
    nor g2678(n898 ,n768 ,n59);
    xnor g2679(n688 ,n472 ,n398);
    nor g2680(n1428 ,n418 ,n818);
    nor g2681(n1134 ,n255 ,n816);
    or g2682(n1957 ,n1344 ,n932);
    not g2683(n119 ,n24[23]);
    or g2684(n1960 ,n1337 ,n1673);
    nor g2685(n865 ,n632 ,n63);
    nor g2686(n1669 ,n395 ,n56);
    or g2687(n2058 ,n1398 ,n1000);
    or g2688(n1814 ,n1199 ,n883);
    dff g2689(.RN(n1), .SN(1'b1), .CK(n0), .D(n1829), .Q(n32[14]));
    or g2690(n2195 ,n1522 ,n863);
    not g2691(n599 ,n15[11]);
    dff g2692(.RN(n1), .SN(1'b1), .CK(n0), .D(n1835), .Q(n32[11]));
    nor g2693(n918 ,n647 ,n55);
    dff g2694(.RN(n1), .SN(1'b1), .CK(n0), .D(n2075), .Q(n21[8]));
    not g2695(n208 ,n31[2]);
    dff g2696(.RN(n1), .SN(1'b1), .CK(n0), .D(n1978), .Q(n34[15]));
    not g2697(n2236 ,n21[20]);
    not g2698(n401 ,n26[12]);
    or g2699(n1863 ,n1033 ,n1581);
    xor g2700(n20[2] ,n23[2] ,n24[2]);
    not g2701(n549 ,n28[10]);
    nor g2702(n1261 ,n489 ,n53);
    nor g2703(n937 ,n694 ,n55);
    dff g2704(.RN(n1), .SN(1'b1), .CK(n0), .D(n1801), .Q(n32[31]));
    or g2705(n1989 ,n1357 ,n1693);
    nor g2706(n896 ,n753 ,n59);
    nor g2707(n1133 ,n230 ,n816);
    nor g2708(n1022 ,n351 ,n818);
    xnor g2709(n805 ,n348 ,n368);
    nor g2710(n1714 ,n443 ,n66);
    or g2711(n1799 ,n1181 ,n1715);
    nor g2712(n1478 ,n262 ,n816);
    dff g2713(.RN(n1), .SN(1'b1), .CK(n0), .D(n2058), .Q(n35[10]));
    not g2714(n203 ,n34[12]);
    or g2715(n1758 ,n1138 ,n942);
    dff g2716(.RN(n1), .SN(1'b1), .CK(n0), .D(n1839), .Q(n26[23]));
    nor g2717(n1273 ,n517 ,n53);
    not g2718(n417 ,n33[9]);
    not g2719(n323 ,n5[31]);
    nor g2720(n1682 ,n147 ,n55);
    not g2721(n137 ,n26[18]);
    or g2722(n1774 ,n1161 ,n1713);
    nor g2723(n1129 ,n562 ,n43);
    not g2724(n142 ,n33[7]);
    nor g2725(n834 ,n786 ,n48);
    nor g2726(n1165 ,n410 ,n67);
    not g2727(n373 ,n30[2]);
    nor g2728(n1183 ,n590 ,n43);
    not g2729(n452 ,n30[27]);
    not g2730(n235 ,n13[18]);
    xnor g2731(n737 ,n21[28] ,n24[28]);
    not g2732(n126 ,n24[12]);
    nor g2733(n1426 ,n119 ,n818);
    dff g2734(.RN(n1), .SN(1'b1), .CK(n0), .D(n1795), .Q(n11[3]));
    nor g2735(n1375 ,n451 ,n816);
    or g2736(n1777 ,n1156 ,n1539);
    nor g2737(n1024 ,n74 ,n51);
    dff g2738(.RN(n1), .SN(1'b1), .CK(n0), .D(n1916), .Q(n35[23]));
    nor g2739(n1587 ,n265 ,n52);
    buf g2740(n14[22], n11[22]);
    not g2741(n91 ,n21[5]);
    nor g2742(n1402 ,n389 ,n61);
    not g2743(n59 ,n58);
    xnor g2744(n689 ,n480 ,n166);
    or g2745(n1866 ,n1244 ,n912);
    nor g2746(n1689 ,n406 ,n64);
    nor g2747(n1152 ,n606 ,n44);
    nor g2748(n1049 ,n357 ,n58);
    not g2749(n442 ,n26[14]);
    nor g2750(n982 ,n664 ,n69);
    dff g2751(.RN(n1), .SN(1'b1), .CK(n0), .D(n1952), .Q(n31[1]));
    nor g2752(n987 ,n692 ,n69);
    nor g2753(n1427 ,n547 ,n57);
    not g2754(n190 ,n34[19]);
    nor g2755(n1088 ,n364 ,n60);
    dff g2756(.RN(n1), .SN(1'b1), .CK(n0), .D(n2177), .Q(n35[28]));
    not g2757(n302 ,n3[30]);
    nor g2758(n1223 ,n108 ,n67);
    xnor g2759(n697 ,n209 ,n127);
    xnor g2760(n655 ,n525 ,n441);
    dff g2761(.RN(n1), .SN(1'b1), .CK(n0), .D(n1864), .Q(n23[0]));
    nor g2762(n1371 ,n483 ,n54);
    or g2763(n2189 ,n1514 ,n859);
    nor g2764(n1154 ,n601 ,n43);
    dff g2765(.RN(n1), .SN(1'b1), .CK(n0), .D(n1806), .Q(n32[28]));
    not g2766(n347 ,n27[0]);
    nor g2767(n1713 ,n390 ,n66);
    not g2768(n609 ,n13[13]);
    or g2769(n1796 ,n1179 ,n1554);
    not g2770(n399 ,n24[1]);
    nor g2771(n901 ,n756 ,n60);
    nor g2772(n1525 ,n455 ,n47);
    or g2773(n1888 ,n1269 ,n924);
    or g2774(n1755 ,n1134 ,n1083);
    nor g2775(n971 ,n795 ,n64);
    or g2776(n1764 ,n1143 ,n1529);
    or g2777(n2017 ,n1372 ,n1705);
    nor g2778(n1062 ,n367 ,n51);
    or g2779(n2076 ,n1417 ,n1119);
    nor g2780(n1679 ,n461 ,n56);
    dff g2781(.RN(n1), .SN(1'b1), .CK(n0), .D(n1859), .Q(n23[3]));
    nor g2782(n62 ,n39 ,n41);
    dff g2783(.RN(n1), .SN(1'b1), .CK(n0), .D(n2103), .Q(n22[2]));
    not g2784(n240 ,n15[8]);
    nor g2785(n1050 ,n500 ,n53);
    nor g2786(n1440 ,n394 ,n818);
    nor g2787(n839 ,n771 ,n47);
    nor g2788(n1231 ,n138 ,n67);
    or g2789(n2310 ,n2295 ,n2297);
    dff g2790(.RN(n1), .SN(1'b1), .CK(n0), .D(n1793), .Q(n11[5]));
    nor g2791(n1308 ,n190 ,n53);
    buf g2792(n15[13], 1'b0);
    nor g2793(n1206 ,n136 ,n57);
    or g2794(n1959 ,n1335 ,n1677);
    or g2795(n1891 ,n1271 ,n925);
    nor g2796(n1476 ,n180 ,n62);
    nor g2797(n1177 ,n427 ,n67);
    or g2798(n2059 ,n1402 ,n948);
    dff g2799(.RN(n1), .SN(1'b1), .CK(n0), .D(n1948), .Q(n31[2]));
    not g2800(n413 ,n32[10]);
    dff g2801(.RN(n1), .SN(1'b1), .CK(n0), .D(n2106), .Q(n24[19]));
    not g2802(n177 ,n31[4]);
    not g2803(n592 ,n11[3]);
    or g2804(n2042 ,n1390 ,n1712);
    nor g2805(n1668 ,n117 ,n56);
    or g2806(n2054 ,n1397 ,n966);
    not g2807(n318 ,n3[28]);
    nor g2808(n970 ,n813 ,n64);
    nor g2809(n1491 ,n263 ,n44);
    dff g2810(.RN(n1), .SN(1'b1), .CK(n0), .D(n2120), .Q(n21[1]));
    not g2811(n409 ,n33[10]);
    xnor g2812(n793 ,n354 ,n96);
    dff g2813(.RN(n1), .SN(1'b1), .CK(n0), .D(n1986), .Q(n30[23]));
    nor g2814(n1635 ,n340 ,n52);
    nor g2815(n1380 ,n102 ,n816);
    not g2816(n2237 ,n24[9]);
    dff g2817(.RN(n1), .SN(1'b1), .CK(n0), .D(n1922), .Q(n31[9]));
    nor g2818(n1497 ,n259 ,n44);
    xnor g2819(n691 ,n201 ,n541);
    dff g2820(.RN(n1), .SN(1'b1), .CK(n0), .D(n2197), .Q(n30[26]));
    not g2821(n259 ,n13[14]);
    dff g2822(.RN(n1), .SN(1'b1), .CK(n0), .D(n2052), .Q(n33[10]));
    buf g2823(n14[28], n12[28]);
    not g2824(n485 ,n34[28]);
    or g2825(n1792 ,n1165 ,n1714);
    nor g2826(n1294 ,n603 ,n819);
    nor g2827(n1640 ,n309 ,n49);
    or g2828(n1767 ,n1144 ,n865);
    nor g2829(n1504 ,n238 ,n65);
    not g2830(n483 ,n34[0]);
    nor g2831(n1344 ,n170 ,n53);
    nor g2832(n1015 ,n72 ,n45);
    nor g2833(n1452 ,n399 ,n818);
    nor g2834(n1306 ,n561 ,n819);
    xnor g2835(n631 ,n471 ,n489);
    or g2836(n1929 ,n1309 ,n999);
    not g2837(n500 ,n31[16]);
    not g2838(n2253 ,n24[14]);
    or g2839(n1772 ,n1438 ,n866);
    not g2840(n536 ,n31[12]);
    not g2841(n551 ,n29[16]);
    not g2842(n113 ,n24[25]);
    not g2843(n479 ,n31[21]);
    not g2844(n284 ,n8[0]);
    not g2845(n73 ,n22[4]);
    dff g2846(.RN(n1), .SN(1'b1), .CK(n0), .D(n2038), .Q(n30[9]));
endmodule
